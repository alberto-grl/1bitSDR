// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.11.2.446
// Netlist written on Mon Apr 06 13:41:19 2020
//
// Verilog Description of module top
//

module top (i_Rx_Serial, o_Tx_Serial, MYLED, XOut, RFIn, DiffOut, 
            PWMOut, PWMOutP1, PWMOutP2, PWMOutP3, PWMOutP4, PWMOutN1, 
            PWMOutN2, PWMOutN3, PWMOutN4, sinGen, sin_out, CIC_out_clkSin) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(45[8:11])
    input i_Rx_Serial;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(47[13:24])
    output o_Tx_Serial;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(48[11:22])
    output [7:0]MYLED;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(49[18:23])
    output XOut;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(53[9:13])
    input RFIn;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(54[9:13])
    output DiffOut;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(55[9:16])
    output PWMOut;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(56[9:15])
    output PWMOutP1;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(57[9:17])
    output PWMOutP2;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(58[9:17])
    output PWMOutP3;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(59[9:17])
    output PWMOutP4;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(60[9:17])
    output PWMOutN1;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(61[9:17])
    output PWMOutN2;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(62[9:17])
    output PWMOutN3;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(63[9:17])
    output PWMOutN4;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(64[9:17])
    output sinGen;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(65[9:15])
    output sin_out;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(66[9:16])
    output CIC_out_clkSin;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(67[9:23])
    
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(69[8:15])
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(85[6:21])
    
    wire GND_net, VCC_net, i_Rx_Serial_c, MYLED_c_6, MYLED_c_5, MYLED_c_4, 
        MYLED_c_3, MYLED_c_2, MYLED_c_1, MYLED_c_0, RFIn_c, DiffOut_c, 
        PWMOutP4_c, PWMOutN4_c, sinGen_c, n2323, o_Rx_DV;
    wire [7:0]o_Rx_Byte;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(73[10:19])
    
    wire o_Rx_DV1;
    wire [7:0]o_Rx_Byte1;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(76[11:21])
    wire [11:0]MixerOutSin;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(81[20:31])
    wire [11:0]MixerOutCos;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(82[20:31])
    wire [11:0]CIC1_outSin;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(84[20:31])
    wire [11:0]CIC1_outCos;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(87[20:31])
    wire [63:0]phase_accum;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(89[13:24])
    wire [12:0]LOSine;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(90[20:26])
    wire [12:0]LOCosine;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(91[20:28])
    wire [63:0]phase_inc_carrGen;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(93[19:36])
    wire [63:0]phase_inc_carrGen1;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(94[19:37])
    wire [11:0]DemodOut;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(97[20:28])
    wire [7:0]CICGain;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(99[11:18])
    
    wire n1154, n1153, n1152, n1151, n1150, n1149, n1148, n1147, 
        n1146, n1145, n1144, n1143, n1142, n1141, n1140, n1139, 
        n1138, n1137, n1136, n1135, n1134, n1133, n1132, n1131, 
        n1130, n1129, n1128, n1127, n1126, n1125, n1124, n1123, 
        n1122, n1121, n1120, n1119, n1118, n1117, n1116, n1115, 
        n1114, n1113, n1112, n1111, n1110, n1109, n1108, n1107, 
        n1106, n1105, n1104, n1103, n1102, n1101, n1100, n1099, 
        n1098, n1097, n1096, n1092, n1093, n1094, n1095, n12533, 
        n7760, n7762, n2384, n2379, n2373, n1032, n1031, n1033, 
        n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, 
        n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, 
        n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, 
        n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, 
        n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, 
        n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, 
        n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, 
        n1090, n11047, n11046, n11045, n11044, n11043, n11042, 
        n11041, n11040, n11039, n11038, n11037, n11036, n11035, 
        n11034, n11033, n11032, n11031, n11030, n11029, n11028, 
        n11027, n11026, n11025, n11024, n11023, n11022, n11021, 
        n11020, n11019, n11018, n11017, n11009, n11008, n11007, 
        n11006, n11005, n11004, n11003, n11002, n11001, n11000, 
        n10999, n10998, n10997, n10996, n10995, n10994, n10993, 
        n10992, n10991, n10990, n10989, n10988, n10987, n10986, 
        n10985, n10984, n10983, n10982, n10981, n10980, n10979, 
        n10978, n10836, n10835, n10834, n10833, n10832, n10831, 
        n10830, n10829, n10828, n10827, n10826, n10825, n10824, 
        n10823, n10822, n10821, n10820, n10819, n10818, n10817, 
        n10816, n10815, n10814, n10813, n10812, n10811, n10810, 
        n10809, n10808, n10807;
    wire [71:0]d10_adj_2554;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(47[26:29])
    wire [71:0]d_out_11__N_1819_adj_2579;
    wire [11:0]DataInReg_11__N_1856;
    
    wire n2325, n2322, n2320, n2319, n2318, n2317, n2316, n2315, 
        n2314, n2313, n2312, n2311, n2309, n2308, n2307, n2306, 
        n2305, n2304, n2303, n2302, n3686, n3682, n3678, n3653, 
        n7603, n3634, n2326, n2327, n8257, n41, n13063, n2328, 
        n2324, n13061, n13060, n13056, n2361, n2360, n2359, n2358, 
        n2357, n2355, n2354, n2353, n2352, n2351, n2350, n2348, 
        n2347, n2346, n2344, n2555, n2551, n2550, n2547, n2541, 
        n2540, n2533, n8391, n2522, n8043, n2512, n13094, n2506, 
        n2505, osc_clk_enable_1411, n13093, n13092, n2628, n2880, 
        n2879, n2878, n2877, n2876, n2875, n2874, n2873, n2872, 
        n2871, n2870, n2869, n2868, n2867, n2866, n2865, n2864, 
        n2863, n2862, n2861, n2860, n2859, n2858, n2857, n2856, 
        n2855, n2854, n2853, n2852, n2851, n2850, n2849, n2848, 
        n2847, n2846, n2845, n2844, n2843, n2842, n61, n62, 
        n63, n64, n65, n66, n67, n68, n70, n2342, n2341, n2340, 
        n2339, n2338, n2337, n2336, n2335, n2334, n2333, n2332, 
        n2331, n2330, n2329, n12947, n2563, n2841, n2840, n2839, 
        n2838, n2837, n2836, n2835, n2834, n2833, n2832, n2831, 
        n2830, n2829, n2828, n2827, n2826, n2825, n2824, n2823, 
        n2822, n2821, n2820, n2819, n2818, n2817, n2815, osc_clk_enable_1471, 
        n12954, n12953, osc_clk_enable_1461, n13212, n13179, n6, 
        n13054, n8252, n7766, n7768, n7770, n7776, n7778, n7782, 
        n7786, n7790, n7792, n7794, n7796, n7798, n7800, n7804, 
        n7806, n7808, n7810, n7812, n7814, n7816, n7818, n7820, 
        n7822, n7826, n7828, n7830, n7832, n7834, n7836, n7840, 
        n7844, n7846, n7852, n7854, n7856, n13068, n13067, n12946, 
        osc_clk_enable_1407, osc_clk_enable_1408, n8041, n8039, n8037, 
        n8035, n8033, n7997, n8031, n8029, n8027;
    
    VHI i2 (.Z(VCC_net));
    PUR PUR_INST (.PUR(VCC_net)) /* synthesis syn_instantiated=1 */ ;
    defparam PUR_INST.RST_PULSE = 1;
    FD1S3AX o_Rx_DV_40 (.D(o_Rx_DV1), .CK(osc_clk), .Q(o_Rx_DV));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam o_Rx_DV_40.GSR = "ENABLED";
    OSCH OSCH_inst (.STDBY(GND_net), .OSC(osc_clk)) /* synthesis syn_instantiated=1 */ ;
    defparam OSCH_inst.NOM_FREQ = "88.67";
    LUT4 mux_322_i15_4_lut (.A(n7776), .B(n1141), .C(n13056), .D(n2563), 
         .Z(n2348)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i15_4_lut.init = 16'hcfca;
    FD1S3AX phase_inc_carrGen1_i0 (.D(phase_inc_carrGen[0]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[0]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i0.GSR = "ENABLED";
    LUT4 n12947_bdd_4_lut (.A(n12947), .B(n12946), .C(MYLED_c_6), .D(o_Rx_Byte[6]), 
         .Z(n13054)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n12947_bdd_4_lut.init = 16'hca00;
    LUT4 mux_322_i43_4_lut (.A(n7826), .B(n1113), .C(n13056), .D(n2563), 
         .Z(n2320)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i43_4_lut.init = 16'hc0ca;
    PWM PWM1 (.osc_clk(osc_clk), .\DataInReg_11__N_1856[0] (DataInReg_11__N_1856[0]), 
        .PWMOutP4_c(PWMOutP4_c), .GND_net(GND_net), .\DemodOut[9] (DemodOut[9]), 
        .\DataInReg_11__N_1856[1] (DataInReg_11__N_1856[1]), .\DataInReg_11__N_1856[2] (DataInReg_11__N_1856[2]), 
        .\DataInReg_11__N_1856[3] (DataInReg_11__N_1856[3]), .\DataInReg_11__N_1856[4] (DataInReg_11__N_1856[4]), 
        .\DataInReg_11__N_1856[5] (DataInReg_11__N_1856[5]), .\DataInReg_11__N_1856[6] (DataInReg_11__N_1856[6]), 
        .\DataInReg_11__N_1856[7] (DataInReg_11__N_1856[7]), .\DataInReg_11__N_1856[8] (DataInReg_11__N_1856[8])) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(189[5] 195[2])
    FD1S3AX phase_inc_carrGen1_i41 (.D(phase_inc_carrGen[41]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[41]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i41.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i40 (.D(phase_inc_carrGen[40]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[40]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i40.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i39 (.D(phase_inc_carrGen[39]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[39]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i39.GSR = "ENABLED";
    LUT4 i1765_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(n13179), 
         .D(n1063), .Z(n7806)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1765_3_lut_4_lut.init = 16'hf404;
    FD1P3AX CICGain__i1 (.D(o_Rx_Byte[0]), .SP(osc_clk_enable_1407), .CK(osc_clk), 
            .Q(CICGain[0]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam CICGain__i1.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i7 (.D(o_Rx_Byte1[7]), .CK(osc_clk), .Q(o_Rx_Byte[7]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam o_Rx_Byte_i7.GSR = "ENABLED";
    LUT4 i1759_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(o_Rx_Byte[3]), 
         .D(n1066), .Z(n7800)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1759_3_lut_4_lut.init = 16'hf404;
    FD1S3AX phase_inc_carrGen1_i38 (.D(phase_inc_carrGen[38]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[38]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i38.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i6 (.D(o_Rx_Byte1[6]), .CK(osc_clk), .Q(o_Rx_Byte[6]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam o_Rx_Byte_i6.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i37 (.D(phase_inc_carrGen[37]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[37]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i37.GSR = "ENABLED";
    LUT4 o_Rx_Byte_4__bdd_3_lut_5467 (.A(o_Rx_Byte[2]), .B(n13179), .C(o_Rx_Byte[0]), 
         .Z(n12947)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam o_Rx_Byte_4__bdd_3_lut_5467.init = 16'h1010;
    FD1S3AX o_Rx_Byte_i5 (.D(o_Rx_Byte1[5]), .CK(osc_clk), .Q(o_Rx_Byte[5]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam o_Rx_Byte_i5.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i36 (.D(phase_inc_carrGen[36]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[36]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i36.GSR = "ENABLED";
    LUT4 mux_322_i44_4_lut (.A(n7828), .B(n1112), .C(n13056), .D(n2563), 
         .Z(n2319)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i44_4_lut.init = 16'hc0ca;
    FD1S3AX o_Rx_Byte_i4 (.D(o_Rx_Byte1[4]), .CK(osc_clk), .Q(o_Rx_Byte[4]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam o_Rx_Byte_i4.GSR = "ENABLED";
    LUT4 mux_322_i41_4_lut (.A(n2522), .B(n1115), .C(n13056), .D(n2563), 
         .Z(n2322)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i41_4_lut.init = 16'hcfca;
    OB MYLED_pad_6 (.I(MYLED_c_6), .O(MYLED[6]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(49[18:23])
    FD1S3AX o_Rx_Byte_i3 (.D(o_Rx_Byte1[3]), .CK(osc_clk), .Q(o_Rx_Byte[3]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam o_Rx_Byte_i3.GSR = "ENABLED";
    LUT4 mux_322_i16_4_lut (.A(n2547), .B(n1140), .C(n13056), .D(n2563), 
         .Z(n2347)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i16_4_lut.init = 16'hcfca;
    LUT4 i1982_4_lut (.A(n1114), .B(n1053), .C(o_Rx_Byte[3]), .D(n13060), 
         .Z(n8035)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1982_4_lut.init = 16'hcac0;
    FD1S3AX phase_inc_carrGen1_i35 (.D(phase_inc_carrGen[35]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[35]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i35.GSR = "ENABLED";
    LUT4 i1787_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(n13179), 
         .D(n1051), .Z(n7828)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1787_3_lut_4_lut.init = 16'hfb0b;
    FD1S3AX phase_inc_carrGen1_i34 (.D(phase_inc_carrGen[34]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[34]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i34.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i33 (.D(phase_inc_carrGen[33]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[33]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i33.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i32 (.D(phase_inc_carrGen[32]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[32]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i32.GSR = "ENABLED";
    LUT4 mux_322_i39_4_lut (.A(n7820), .B(n1117), .C(n13056), .D(n2563), 
         .Z(n2324)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i39_4_lut.init = 16'hc0ca;
    FD1S3AX phase_inc_carrGen1_i31 (.D(phase_inc_carrGen[31]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[31]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i31.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i30 (.D(phase_inc_carrGen[30]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[30]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i30.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i2 (.D(o_Rx_Byte1[2]), .CK(osc_clk), .Q(o_Rx_Byte[2]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam o_Rx_Byte_i2.GSR = "ENABLED";
    LUT4 mux_322_i40_4_lut (.A(n7822), .B(n1116), .C(n13056), .D(n2563), 
         .Z(n2323)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i40_4_lut.init = 16'hcfca;
    FD1S3AX phase_inc_carrGen1_i29 (.D(phase_inc_carrGen[29]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[29]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i29.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i28 (.D(phase_inc_carrGen[28]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[28]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i28.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i27 (.D(phase_inc_carrGen[27]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[27]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i27.GSR = "ENABLED";
    LUT4 mux_322_i37_4_lut (.A(n7816), .B(n1119), .C(n13056), .D(n2563), 
         .Z(n2326)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i37_4_lut.init = 16'hcfca;
    LUT4 i1767_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(o_Rx_Byte[3]), 
         .D(n1062), .Z(n7808)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1767_3_lut_4_lut.init = 16'hfb0b;
    LUT4 n2644_bdd_4_lut_5398 (.A(o_Rx_Byte[0]), .B(o_Rx_Byte[4]), .C(MYLED_c_6), 
         .D(o_Rx_Byte[3]), .Z(n12954)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam n2644_bdd_4_lut_5398.init = 16'h0004;
    LUT4 i1749_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(n13179), 
         .D(n1071), .Z(n7790)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1749_3_lut_4_lut.init = 16'hf404;
    LUT4 mux_322_i13_4_lut (.A(n2550), .B(n1143), .C(n13056), .D(n2563), 
         .Z(n2350)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i13_4_lut.init = 16'hc0ca;
    LUT4 i1976_4_lut (.A(n1142), .B(n1081), .C(o_Rx_Byte[3]), .D(n13060), 
         .Z(n8029)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1976_4_lut.init = 16'hcac0;
    LUT4 mux_322_i11_4_lut (.A(n7770), .B(n1145), .C(n13056), .D(n2563), 
         .Z(n2352)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i11_4_lut.init = 16'hcfca;
    FD1S3AX phase_inc_carrGen1_i26 (.D(phase_inc_carrGen[26]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[26]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i26.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i25 (.D(phase_inc_carrGen[25]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[25]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i25.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i24 (.D(phase_inc_carrGen[24]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[24]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i24.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i1 (.D(o_Rx_Byte1[1]), .CK(osc_clk), .Q(MYLED_c_6));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam o_Rx_Byte_i1.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i23 (.D(phase_inc_carrGen[23]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[23]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i23.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i22 (.D(phase_inc_carrGen[22]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[22]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i22.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i21 (.D(phase_inc_carrGen[21]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[21]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i21.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i20 (.D(phase_inc_carrGen[20]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[20]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i20.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i19 (.D(phase_inc_carrGen[19]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[19]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i19.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i18 (.D(phase_inc_carrGen[18]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[18]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i18.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i17 (.D(phase_inc_carrGen[17]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[17]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i17.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i16 (.D(phase_inc_carrGen[16]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[16]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i16.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i15 (.D(phase_inc_carrGen[15]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[15]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i15.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i14 (.D(phase_inc_carrGen[14]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[14]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i14.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i13 (.D(phase_inc_carrGen[13]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[13]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i13.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i12 (.D(phase_inc_carrGen[12]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[12]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i12.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i11 (.D(phase_inc_carrGen[11]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[11]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i11.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i10 (.D(phase_inc_carrGen[10]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[10]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i10.GSR = "ENABLED";
    LUT4 i2579_2_lut (.A(o_Rx_Byte[4]), .B(n2815), .Z(n3682)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i2579_2_lut.init = 16'hbbbb;
    LUT4 mux_322_i12_4_lut (.A(n2551), .B(n1144), .C(n13056), .D(n2563), 
         .Z(n2351)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i12_4_lut.init = 16'hcfca;
    LUT4 i2720_2_lut (.A(n1083), .B(o_Rx_Byte[3]), .Z(n2551)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i2720_2_lut.init = 16'h8888;
    LUT4 mux_322_i38_4_lut (.A(n7818), .B(n1118), .C(n13056), .D(n2563), 
         .Z(n2325)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i38_4_lut.init = 16'hc0ca;
    LUT4 mux_322_i9_4_lut (.A(n7766), .B(n1147), .C(n13056), .D(n2563), 
         .Z(n2354)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i9_4_lut.init = 16'hcfca;
    LUT4 mux_322_i10_4_lut (.A(n7768), .B(n1146), .C(n13056), .D(n2563), 
         .Z(n2353)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i10_4_lut.init = 16'hcfca;
    FD1S3AX phase_inc_carrGen1_i9 (.D(phase_inc_carrGen[9]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[9]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i9.GSR = "ENABLED";
    LUT4 i1974_4_lut (.A(n1149), .B(n1088), .C(o_Rx_Byte[3]), .D(n13060), 
         .Z(n8027)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1974_4_lut.init = 16'hcacf;
    LUT4 i1737_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(o_Rx_Byte[3]), 
         .D(n1078), .Z(n7778)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1737_3_lut_4_lut.init = 16'hf404;
    LUT4 mux_322_i8_4_lut (.A(n2555), .B(n1148), .C(n13056), .D(n2563), 
         .Z(n2355)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i8_4_lut.init = 16'hcfca;
    LUT4 mux_322_i35_4_lut (.A(n7812), .B(n1121), .C(n13056), .D(n2563), 
         .Z(n2328)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i35_4_lut.init = 16'hcfca;
    LUT4 mux_322_i5_4_lut (.A(n7760), .B(n1151), .C(n13056), .D(n2563), 
         .Z(n2358)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i5_4_lut.init = 16'hc0ca;
    LUT4 mux_322_i6_4_lut (.A(n7762), .B(n1150), .C(n13056), .D(n2563), 
         .Z(n2357)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i6_4_lut.init = 16'hcfca;
    FD1S3AX phase_inc_carrGen1_i8 (.D(phase_inc_carrGen[8]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[8]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i8.GSR = "ENABLED";
    LUT4 mux_322_i36_4_lut (.A(n7814), .B(n1120), .C(n13056), .D(n2563), 
         .Z(n2327)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i36_4_lut.init = 16'hcfca;
    FD1S3AX phase_inc_carrGen1_i7 (.D(phase_inc_carrGen[7]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[7]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i7.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i6 (.D(phase_inc_carrGen[6]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[6]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i6.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i5 (.D(phase_inc_carrGen[5]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[5]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i5.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i4 (.D(phase_inc_carrGen[4]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[4]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i4.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i3 (.D(phase_inc_carrGen[3]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[3]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i3.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i2 (.D(phase_inc_carrGen[2]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[2]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i2.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i1 (.D(phase_inc_carrGen[1]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[1]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i1.GSR = "ENABLED";
    OB MYLED_pad_5 (.I(MYLED_c_5), .O(MYLED[5]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(49[18:23])
    LUT4 mux_322_i33_4_lut (.A(n7808), .B(n1123), .C(n13056), .D(n2563), 
         .Z(n2330)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i33_4_lut.init = 16'hc0ca;
    LUT4 i1_3_lut (.A(o_Rx_Byte[3]), .B(n13063), .C(o_Rx_Byte[2]), .Z(n2628)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_3_lut.init = 16'h4040;
    LUT4 mux_322_i2_4_lut (.A(n8391), .B(n1154), .C(n13056), .D(n2563), 
         .Z(n2361)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i2_4_lut.init = 16'hcfc5;
    LUT4 mux_322_i34_4_lut (.A(n7810), .B(n1122), .C(n13056), .D(n2563), 
         .Z(n2329)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i34_4_lut.init = 16'hcfca;
    LUT4 i1729_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(n13179), 
         .D(n1084), .Z(n7770)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1729_3_lut_4_lut.init = 16'hf404;
    LUT4 i1769_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(n13179), 
         .D(n1061), .Z(n7810)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1769_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i1751_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(o_Rx_Byte[3]), 
         .D(n1070), .Z(n7792)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1751_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i1719_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(n13179), 
         .D(n1090), .Z(n7760)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1719_3_lut_4_lut.init = 16'hf404;
    LUT4 mux_322_i31_4_lut (.A(n7804), .B(n1125), .C(n13056), .D(n2563), 
         .Z(n2332)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i31_4_lut.init = 16'hc0ca;
    LUT4 mux_747_i2_3_lut (.A(o_Rx_Byte[2]), .B(o_Rx_Byte[4]), .C(n2815), 
         .Z(n3686)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_747_i2_3_lut.init = 16'hc5c5;
    LUT4 i1803_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(o_Rx_Byte[3]), 
         .D(n1041), .Z(n7844)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1803_3_lut_4_lut.init = 16'hf707;
    LUT4 mux_322_i32_4_lut (.A(n7806), .B(n1124), .C(n13056), .D(n2563), 
         .Z(n2331)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i32_4_lut.init = 16'hcfca;
    LUT4 mux_322_i29_4_lut (.A(n7800), .B(n1127), .C(n13056), .D(n2563), 
         .Z(n2334)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i29_4_lut.init = 16'hc0ca;
    LUT4 mux_322_i30_4_lut (.A(n2533), .B(n1126), .C(n13056), .D(n2563), 
         .Z(n2333)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i30_4_lut.init = 16'hc0ca;
    OB MYLED_pad_7 (.I(GND_net), .O(MYLED[7]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(49[18:23])
    OB o_Tx_Serial_pad (.I(GND_net), .O(o_Tx_Serial));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(48[11:22])
    \uart_rx(CLKS_PER_BIT=87)  uart_rx1 (.osc_clk(osc_clk), .i_Rx_Serial_c(i_Rx_Serial_c), 
            .o_Rx_Byte1({o_Rx_Byte1}), .GND_net(GND_net), .o_Rx_DV1(o_Rx_DV1)) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(220[32] 225[2])
    LUT4 i5373_4_lut_rep_131 (.A(n13067), .B(n8252), .C(o_Rx_Byte[6]), 
         .D(n13094), .Z(n13212)) /* synthesis lut_function=(!(A+!(B (C)+!B (C (D))))) */ ;
    defparam i5373_4_lut_rep_131.init = 16'h5040;
    OB MYLED_pad_4 (.I(MYLED_c_4), .O(MYLED[4]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(49[18:23])
    OB MYLED_pad_3 (.I(MYLED_c_3), .O(MYLED[3]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(49[18:23])
    OB MYLED_pad_2 (.I(MYLED_c_2), .O(MYLED[2]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(49[18:23])
    OB MYLED_pad_1 (.I(MYLED_c_1), .O(MYLED[1]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(49[18:23])
    OB MYLED_pad_0 (.I(MYLED_c_0), .O(MYLED[0]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(49[18:23])
    OB XOut_pad (.I(GND_net), .O(XOut));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(53[9:13])
    OB DiffOut_pad (.I(DiffOut_c), .O(DiffOut));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(55[9:16])
    OB PWMOut_pad (.I(PWMOutP4_c), .O(PWMOut));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(56[9:15])
    OB PWMOutP1_pad (.I(PWMOutP4_c), .O(PWMOutP1));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(57[9:17])
    OB PWMOutP2_pad (.I(PWMOutP4_c), .O(PWMOutP2));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(58[9:17])
    OB PWMOutP3_pad (.I(PWMOutP4_c), .O(PWMOutP3));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(59[9:17])
    OB PWMOutP4_pad (.I(PWMOutP4_c), .O(PWMOutP4));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(60[9:17])
    OB PWMOutN1_pad (.I(PWMOutN4_c), .O(PWMOutN1));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(61[9:17])
    OB PWMOutN2_pad (.I(PWMOutN4_c), .O(PWMOutN2));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(62[9:17])
    OB PWMOutN3_pad (.I(PWMOutN4_c), .O(PWMOutN3));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(63[9:17])
    OB PWMOutN4_pad (.I(PWMOutN4_c), .O(PWMOutN4));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(64[9:17])
    OB sinGen_pad (.I(sinGen_c), .O(sinGen));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(65[9:15])
    OB sin_out_pad (.I(GND_net), .O(sin_out));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(66[9:16])
    OB CIC_out_clkSin_pad (.I(GND_net), .O(CIC_out_clkSin));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(67[9:23])
    IB i_Rx_Serial_pad (.I(i_Rx_Serial), .O(i_Rx_Serial_c));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(47[13:24])
    IB RFIn_pad (.I(RFIn), .O(RFIn_c));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(54[9:13])
    LUT4 i1_3_lut_rep_93 (.A(o_Rx_DV), .B(o_Rx_Byte[5]), .C(o_Rx_Byte[7]), 
         .Z(n13067)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_3_lut_rep_93.init = 16'hf7f7;
    LUT4 i1_2_lut_rep_87_4_lut (.A(o_Rx_DV), .B(o_Rx_Byte[5]), .C(o_Rx_Byte[7]), 
         .D(n13054), .Z(n13061)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_87_4_lut.init = 16'h0800;
    LUT4 i1_2_lut_4_lut (.A(o_Rx_DV), .B(o_Rx_Byte[5]), .C(o_Rx_Byte[7]), 
         .D(o_Rx_Byte[4]), .Z(n6)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam i1_2_lut_4_lut.init = 16'hf7ff;
    LUT4 i1741_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(o_Rx_Byte[3]), 
         .D(n1076), .Z(n7782)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1741_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i1_2_lut_rep_94 (.A(MYLED_c_6), .B(o_Rx_Byte[0]), .Z(n13068)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam i1_2_lut_rep_94.init = 16'h2222;
    LUT4 i1_3_lut_rep_89_3_lut_4_lut (.A(MYLED_c_6), .B(o_Rx_Byte[0]), .C(n8257), 
         .D(o_Rx_Byte[4]), .Z(n13063)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam i1_3_lut_rep_89_3_lut_4_lut.init = 16'h0020;
    LUT4 i2727_2_lut (.A(n1065), .B(n13179), .Z(n2533)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i2727_2_lut.init = 16'hbbbb;
    LUT4 i1815_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(n13179), 
         .D(n1034), .Z(n7856)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1815_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i1811_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(o_Rx_Byte[3]), 
         .D(n1036), .Z(n7852)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1811_3_lut_4_lut.init = 16'hfb0b;
    FD1S3AX phase_inc_carrGen1_i42 (.D(phase_inc_carrGen[42]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[42]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i42.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i43 (.D(phase_inc_carrGen[43]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[43]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i43.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i44 (.D(phase_inc_carrGen[44]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[44]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i44.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i45 (.D(phase_inc_carrGen[45]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[45]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i45.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i46 (.D(phase_inc_carrGen[46]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[46]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i46.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i47 (.D(phase_inc_carrGen[47]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[47]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i47.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i48 (.D(phase_inc_carrGen[48]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[48]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i48.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i49 (.D(phase_inc_carrGen[49]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[49]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i49.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i50 (.D(phase_inc_carrGen[50]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[50]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i50.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i51 (.D(phase_inc_carrGen[51]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[51]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i51.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i52 (.D(phase_inc_carrGen[52]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[52]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i52.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i53 (.D(phase_inc_carrGen[53]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[53]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i53.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i54 (.D(phase_inc_carrGen[54]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[54]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i54.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i55 (.D(phase_inc_carrGen[55]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[55]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i55.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i56 (.D(phase_inc_carrGen[56]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[56]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i56.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i57 (.D(phase_inc_carrGen[57]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[57]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i57.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i58 (.D(phase_inc_carrGen[58]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[58]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i58.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i59 (.D(phase_inc_carrGen[59]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[59]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i59.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i60 (.D(phase_inc_carrGen[60]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[60]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i60.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i61 (.D(phase_inc_carrGen[61]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[61]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i61.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i62 (.D(phase_inc_carrGen[62]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[62]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i62.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i63 (.D(phase_inc_carrGen[63]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[63]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen1_i63.GSR = "ENABLED";
    FD1P3AX CICGain__i2 (.D(MYLED_c_6), .SP(osc_clk_enable_1407), .CK(osc_clk), 
            .Q(CICGain[1]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam CICGain__i2.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i0 (.D(n2880), .SP(osc_clk_enable_1408), 
            .CK(osc_clk), .Q(phase_inc_carrGen[0]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i0.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i1 (.D(n2879), .SP(osc_clk_enable_1411), 
            .CK(osc_clk), .Q(phase_inc_carrGen[1]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i1.GSR = "ENABLED";
    LUT4 i5373_4_lut_rep_132 (.A(n13067), .B(n8252), .C(o_Rx_Byte[6]), 
         .D(n13094), .Z(osc_clk_enable_1461)) /* synthesis lut_function=(!(A+!(B (C)+!B (C (D))))) */ ;
    defparam i5373_4_lut_rep_132.init = 16'h5040;
    LUT4 i5364_4_lut (.A(n13212), .B(o_Rx_Byte[3]), .C(n13061), .D(n13060), 
         .Z(osc_clk_enable_1408)) /* synthesis lut_function=(!((B (C)+!B (C (D)))+!A)) */ ;
    defparam i5364_4_lut.init = 16'h0a2a;
    LUT4 i1795_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(o_Rx_Byte[3]), 
         .D(n1046), .Z(n7836)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1795_3_lut_4_lut.init = 16'hf808;
    LUT4 i5373_4_lut (.A(n13067), .B(n8252), .C(o_Rx_Byte[6]), .D(n13094), 
         .Z(osc_clk_enable_1471)) /* synthesis lut_function=(!(A+!(B (C)+!B (C (D))))) */ ;
    defparam i5373_4_lut.init = 16'h5040;
    LUT4 i1_4_lut (.A(n41), .B(o_Rx_Byte[2]), .C(o_Rx_Byte[3]), .D(MYLED_c_6), 
         .Z(n8252)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (B+((D)+!C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(271[4] 285[10])
    defparam i1_4_lut.init = 16'h0012;
    CCU2D sub_46_add_2_63 (.A0(phase_inc_carrGen[62]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[63]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11047), .S0(n1093), .S1(n1092));
    defparam sub_46_add_2_63.INIT0 = 16'h5555;
    defparam sub_46_add_2_63.INIT1 = 16'h5555;
    defparam sub_46_add_2_63.INJECT1_0 = "NO";
    defparam sub_46_add_2_63.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_61 (.A0(phase_inc_carrGen[60]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[61]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11046), .COUT(n11047), .S0(n1095), .S1(n1094));
    defparam sub_46_add_2_61.INIT0 = 16'h5555;
    defparam sub_46_add_2_61.INIT1 = 16'h5555;
    defparam sub_46_add_2_61.INJECT1_0 = "NO";
    defparam sub_46_add_2_61.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_59 (.A0(phase_inc_carrGen[58]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[59]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11045), .COUT(n11046), .S0(n1097), .S1(n1096));
    defparam sub_46_add_2_59.INIT0 = 16'h5555;
    defparam sub_46_add_2_59.INIT1 = 16'h5555;
    defparam sub_46_add_2_59.INJECT1_0 = "NO";
    defparam sub_46_add_2_59.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_57 (.A0(phase_inc_carrGen[56]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[57]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11044), .COUT(n11045), .S0(n1099), .S1(n1098));
    defparam sub_46_add_2_57.INIT0 = 16'h5555;
    defparam sub_46_add_2_57.INIT1 = 16'h5555;
    defparam sub_46_add_2_57.INJECT1_0 = "NO";
    defparam sub_46_add_2_57.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_55 (.A0(phase_inc_carrGen[54]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[55]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11043), .COUT(n11044), .S0(n1101), .S1(n1100));
    defparam sub_46_add_2_55.INIT0 = 16'h5555;
    defparam sub_46_add_2_55.INIT1 = 16'h5555;
    defparam sub_46_add_2_55.INJECT1_0 = "NO";
    defparam sub_46_add_2_55.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_53 (.A0(phase_inc_carrGen[52]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[53]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11042), .COUT(n11043), .S0(n1103), .S1(n1102));
    defparam sub_46_add_2_53.INIT0 = 16'h5555;
    defparam sub_46_add_2_53.INIT1 = 16'h5555;
    defparam sub_46_add_2_53.INJECT1_0 = "NO";
    defparam sub_46_add_2_53.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_51 (.A0(phase_inc_carrGen[50]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[51]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11041), .COUT(n11042), .S0(n1105), .S1(n1104));
    defparam sub_46_add_2_51.INIT0 = 16'h5aaa;
    defparam sub_46_add_2_51.INIT1 = 16'h5aaa;
    defparam sub_46_add_2_51.INJECT1_0 = "NO";
    defparam sub_46_add_2_51.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_49 (.A0(phase_inc_carrGen[48]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[49]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11040), .COUT(n11041), .S0(n1107), .S1(n1106));
    defparam sub_46_add_2_49.INIT0 = 16'h5555;
    defparam sub_46_add_2_49.INIT1 = 16'h5555;
    defparam sub_46_add_2_49.INJECT1_0 = "NO";
    defparam sub_46_add_2_49.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_47 (.A0(phase_inc_carrGen[46]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[47]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11039), .COUT(n11040), .S0(n1109), .S1(n1108));
    defparam sub_46_add_2_47.INIT0 = 16'h5555;
    defparam sub_46_add_2_47.INIT1 = 16'h5aaa;
    defparam sub_46_add_2_47.INJECT1_0 = "NO";
    defparam sub_46_add_2_47.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_45 (.A0(phase_inc_carrGen[44]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[45]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11038), .COUT(n11039), .S0(n1111), .S1(n1110));
    defparam sub_46_add_2_45.INIT0 = 16'h5555;
    defparam sub_46_add_2_45.INIT1 = 16'h5aaa;
    defparam sub_46_add_2_45.INJECT1_0 = "NO";
    defparam sub_46_add_2_45.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_43 (.A0(phase_inc_carrGen[42]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[43]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11037), .COUT(n11038), .S0(n1113), .S1(n1112));
    defparam sub_46_add_2_43.INIT0 = 16'h5555;
    defparam sub_46_add_2_43.INIT1 = 16'h5555;
    defparam sub_46_add_2_43.INJECT1_0 = "NO";
    defparam sub_46_add_2_43.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_41 (.A0(phase_inc_carrGen[40]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[41]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11036), .COUT(n11037), .S0(n1115), .S1(n1114));
    defparam sub_46_add_2_41.INIT0 = 16'h5555;
    defparam sub_46_add_2_41.INIT1 = 16'h5aaa;
    defparam sub_46_add_2_41.INJECT1_0 = "NO";
    defparam sub_46_add_2_41.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_39 (.A0(phase_inc_carrGen[38]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[39]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11035), .COUT(n11036), .S0(n1117), .S1(n1116));
    defparam sub_46_add_2_39.INIT0 = 16'h5555;
    defparam sub_46_add_2_39.INIT1 = 16'h5555;
    defparam sub_46_add_2_39.INJECT1_0 = "NO";
    defparam sub_46_add_2_39.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_37 (.A0(phase_inc_carrGen[36]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[37]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11034), .COUT(n11035), .S0(n1119), .S1(n1118));
    defparam sub_46_add_2_37.INIT0 = 16'h5555;
    defparam sub_46_add_2_37.INIT1 = 16'h5aaa;
    defparam sub_46_add_2_37.INJECT1_0 = "NO";
    defparam sub_46_add_2_37.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_35 (.A0(phase_inc_carrGen[34]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[35]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11033), .COUT(n11034), .S0(n1121), .S1(n1120));
    defparam sub_46_add_2_35.INIT0 = 16'h5555;
    defparam sub_46_add_2_35.INIT1 = 16'h5aaa;
    defparam sub_46_add_2_35.INJECT1_0 = "NO";
    defparam sub_46_add_2_35.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_33 (.A0(phase_inc_carrGen[32]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[33]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11032), .COUT(n11033), .S0(n1123), .S1(n1122));
    defparam sub_46_add_2_33.INIT0 = 16'h5aaa;
    defparam sub_46_add_2_33.INIT1 = 16'h5555;
    defparam sub_46_add_2_33.INJECT1_0 = "NO";
    defparam sub_46_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_31 (.A0(phase_inc_carrGen[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11031), .COUT(n11032), .S0(n1125), .S1(n1124));
    defparam sub_46_add_2_31.INIT0 = 16'h5555;
    defparam sub_46_add_2_31.INIT1 = 16'h5aaa;
    defparam sub_46_add_2_31.INJECT1_0 = "NO";
    defparam sub_46_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_29 (.A0(phase_inc_carrGen[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11030), .COUT(n11031), .S0(n1127), .S1(n1126));
    defparam sub_46_add_2_29.INIT0 = 16'h5555;
    defparam sub_46_add_2_29.INIT1 = 16'h5555;
    defparam sub_46_add_2_29.INJECT1_0 = "NO";
    defparam sub_46_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_27 (.A0(phase_inc_carrGen[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11029), .COUT(n11030), .S0(n1129), .S1(n1128));
    defparam sub_46_add_2_27.INIT0 = 16'h5555;
    defparam sub_46_add_2_27.INIT1 = 16'h5555;
    defparam sub_46_add_2_27.INJECT1_0 = "NO";
    defparam sub_46_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_25 (.A0(phase_inc_carrGen[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11028), .COUT(n11029), .S0(n1131), .S1(n1130));
    defparam sub_46_add_2_25.INIT0 = 16'h5555;
    defparam sub_46_add_2_25.INIT1 = 16'h5555;
    defparam sub_46_add_2_25.INJECT1_0 = "NO";
    defparam sub_46_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_23 (.A0(phase_inc_carrGen[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11027), .COUT(n11028), .S0(n1133), .S1(n1132));
    defparam sub_46_add_2_23.INIT0 = 16'h5555;
    defparam sub_46_add_2_23.INIT1 = 16'h5aaa;
    defparam sub_46_add_2_23.INJECT1_0 = "NO";
    defparam sub_46_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_21 (.A0(phase_inc_carrGen[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11026), .COUT(n11027), .S0(n1135), .S1(n1134));
    defparam sub_46_add_2_21.INIT0 = 16'h5aaa;
    defparam sub_46_add_2_21.INIT1 = 16'h5aaa;
    defparam sub_46_add_2_21.INJECT1_0 = "NO";
    defparam sub_46_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_19 (.A0(phase_inc_carrGen[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11025), .COUT(n11026), .S0(n1137), .S1(n1136));
    defparam sub_46_add_2_19.INIT0 = 16'h5555;
    defparam sub_46_add_2_19.INIT1 = 16'h5aaa;
    defparam sub_46_add_2_19.INJECT1_0 = "NO";
    defparam sub_46_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_17 (.A0(phase_inc_carrGen[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11024), .COUT(n11025), .S0(n1139), .S1(n1138));
    defparam sub_46_add_2_17.INIT0 = 16'h5555;
    defparam sub_46_add_2_17.INIT1 = 16'h5aaa;
    defparam sub_46_add_2_17.INJECT1_0 = "NO";
    defparam sub_46_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_15 (.A0(phase_inc_carrGen[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11023), .COUT(n11024), .S0(n1141), .S1(n1140));
    defparam sub_46_add_2_15.INIT0 = 16'h5aaa;
    defparam sub_46_add_2_15.INIT1 = 16'h5555;
    defparam sub_46_add_2_15.INJECT1_0 = "NO";
    defparam sub_46_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_13 (.A0(phase_inc_carrGen[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11022), .COUT(n11023), .S0(n1143), .S1(n1142));
    defparam sub_46_add_2_13.INIT0 = 16'h5aaa;
    defparam sub_46_add_2_13.INIT1 = 16'h5555;
    defparam sub_46_add_2_13.INJECT1_0 = "NO";
    defparam sub_46_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_11 (.A0(phase_inc_carrGen[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11021), .COUT(n11022), .S0(n1145), .S1(n1144));
    defparam sub_46_add_2_11.INIT0 = 16'h5aaa;
    defparam sub_46_add_2_11.INIT1 = 16'h5555;
    defparam sub_46_add_2_11.INJECT1_0 = "NO";
    defparam sub_46_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_9 (.A0(phase_inc_carrGen[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11020), .COUT(n11021), .S0(n1147), .S1(n1146));
    defparam sub_46_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_46_add_2_9.INIT1 = 16'h5aaa;
    defparam sub_46_add_2_9.INJECT1_0 = "NO";
    defparam sub_46_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_7 (.A0(phase_inc_carrGen[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11019), .COUT(n11020), .S0(n1149), .S1(n1148));
    defparam sub_46_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_46_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_46_add_2_7.INJECT1_0 = "NO";
    defparam sub_46_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_5 (.A0(phase_inc_carrGen[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11018), .COUT(n11019), .S0(n1151), .S1(n1150));
    defparam sub_46_add_2_5.INIT0 = 16'h5555;
    defparam sub_46_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_46_add_2_5.INJECT1_0 = "NO";
    defparam sub_46_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_3 (.A0(phase_inc_carrGen[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11017), .COUT(n11018), .S0(n1153), .S1(n1152));
    defparam sub_46_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_46_add_2_3.INIT1 = 16'h5555;
    defparam sub_46_add_2_3.INJECT1_0 = "NO";
    defparam sub_46_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(phase_inc_carrGen[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n11017), .S1(n1154));
    defparam sub_46_add_2_1.INIT0 = 16'hF000;
    defparam sub_46_add_2_1.INIT1 = 16'h5555;
    defparam sub_46_add_2_1.INJECT1_0 = "NO";
    defparam sub_46_add_2_1.INJECT1_1 = "NO";
    CCU2D add_749_65 (.A0(n3634), .B0(n13061), .C0(n8041), .D0(phase_inc_carrGen[62]), 
          .A1(n3634), .B1(n13061), .C1(n8043), .D1(phase_inc_carrGen[63]), 
          .CIN(n11009), .S0(n2818), .S1(n2817));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_65.INIT0 = 16'hd1e2;
    defparam add_749_65.INIT1 = 16'hd1e2;
    defparam add_749_65.INJECT1_0 = "NO";
    defparam add_749_65.INJECT1_1 = "NO";
    CCU2D add_749_63 (.A0(n3634), .B0(n13061), .C0(n2302), .D0(phase_inc_carrGen[60]), 
          .A1(n3634), .B1(n13061), .C1(n8039), .D1(phase_inc_carrGen[61]), 
          .CIN(n11008), .COUT(n11009), .S0(n2820), .S1(n2819));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_63.INIT0 = 16'hd1e2;
    defparam add_749_63.INIT1 = 16'hd1e2;
    defparam add_749_63.INJECT1_0 = "NO";
    defparam add_749_63.INJECT1_1 = "NO";
    CCU2D add_749_61 (.A0(n3634), .B0(n13061), .C0(n2304), .D0(phase_inc_carrGen[58]), 
          .A1(n3634), .B1(n13061), .C1(n2303), .D1(phase_inc_carrGen[59]), 
          .CIN(n11007), .COUT(n11008), .S0(n2822), .S1(n2821));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_61.INIT0 = 16'hd1e2;
    defparam add_749_61.INIT1 = 16'hd1e2;
    defparam add_749_61.INJECT1_0 = "NO";
    defparam add_749_61.INJECT1_1 = "NO";
    CCU2D add_749_59 (.A0(n3634), .B0(n13061), .C0(n2306), .D0(phase_inc_carrGen[56]), 
          .A1(n3634), .B1(n13061), .C1(n2305), .D1(phase_inc_carrGen[57]), 
          .CIN(n11006), .COUT(n11007), .S0(n2824), .S1(n2823));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_59.INIT0 = 16'hd1e2;
    defparam add_749_59.INIT1 = 16'hd1e2;
    defparam add_749_59.INJECT1_0 = "NO";
    defparam add_749_59.INJECT1_1 = "NO";
    CCU2D add_749_57 (.A0(n3634), .B0(n13061), .C0(n2308), .D0(phase_inc_carrGen[54]), 
          .A1(n3634), .B1(n13061), .C1(n2307), .D1(phase_inc_carrGen[55]), 
          .CIN(n11005), .COUT(n11006), .S0(n2826), .S1(n2825));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_57.INIT0 = 16'hd1e2;
    defparam add_749_57.INIT1 = 16'hd1e2;
    defparam add_749_57.INJECT1_0 = "NO";
    defparam add_749_57.INJECT1_1 = "NO";
    CCU2D add_749_55 (.A0(n3634), .B0(n13061), .C0(n8037), .D0(phase_inc_carrGen[52]), 
          .A1(n3634), .B1(n13061), .C1(n2309), .D1(phase_inc_carrGen[53]), 
          .CIN(n11004), .COUT(n11005), .S0(n2828), .S1(n2827));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_55.INIT0 = 16'hd1e2;
    defparam add_749_55.INIT1 = 16'hd1e2;
    defparam add_749_55.INJECT1_0 = "NO";
    defparam add_749_55.INJECT1_1 = "NO";
    CCU2D add_749_53 (.A0(n13061), .B0(n3678), .C0(n2312), .D0(phase_inc_carrGen[50]), 
          .A1(n13061), .B1(n7603), .C1(n2311), .D1(phase_inc_carrGen[51]), 
          .CIN(n11003), .COUT(n11004), .S0(n2830), .S1(n2829));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_53.INIT0 = 16'he4b1;
    defparam add_749_53.INIT1 = 16'he4b1;
    defparam add_749_53.INJECT1_0 = "NO";
    defparam add_749_53.INJECT1_1 = "NO";
    CCU2D add_749_51 (.A0(n3653), .B0(n13061), .C0(n2314), .D0(phase_inc_carrGen[48]), 
          .A1(n3653), .B1(n13061), .C1(n2313), .D1(phase_inc_carrGen[49]), 
          .CIN(n11002), .COUT(n11003), .S0(n2832), .S1(n2831));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_51.INIT0 = 16'hd1e2;
    defparam add_749_51.INIT1 = 16'hd1e2;
    defparam add_749_51.INJECT1_0 = "NO";
    defparam add_749_51.INJECT1_1 = "NO";
    CCU2D add_749_49 (.A0(n3634), .B0(n13061), .C0(n2316), .D0(phase_inc_carrGen[46]), 
          .A1(n13061), .B1(n7603), .C1(n2315), .D1(phase_inc_carrGen[47]), 
          .CIN(n11001), .COUT(n11002), .S0(n2834), .S1(n2833));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_49.INIT0 = 16'hd1e2;
    defparam add_749_49.INIT1 = 16'he4b1;
    defparam add_749_49.INJECT1_0 = "NO";
    defparam add_749_49.INJECT1_1 = "NO";
    CCU2D add_749_47 (.A0(n7603), .B0(n13061), .C0(n2318), .D0(phase_inc_carrGen[44]), 
          .A1(n13061), .B1(n7603), .C1(n2317), .D1(phase_inc_carrGen[45]), 
          .CIN(n11000), .COUT(n11001), .S0(n2836), .S1(n2835));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_47.INIT0 = 16'hd1e2;
    defparam add_749_47.INIT1 = 16'he4b1;
    defparam add_749_47.INJECT1_0 = "NO";
    defparam add_749_47.INJECT1_1 = "NO";
    CCU2D add_749_45 (.A0(n3678), .B0(n13061), .C0(n2320), .D0(phase_inc_carrGen[42]), 
          .A1(n3653), .B1(n13061), .C1(n2319), .D1(phase_inc_carrGen[43]), 
          .CIN(n10999), .COUT(n11000), .S0(n2838), .S1(n2837));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_45.INIT0 = 16'hd1e2;
    defparam add_749_45.INIT1 = 16'hd1e2;
    defparam add_749_45.INJECT1_0 = "NO";
    defparam add_749_45.INJECT1_1 = "NO";
    CCU2D add_749_43 (.A0(n3653), .B0(n13061), .C0(n2322), .D0(phase_inc_carrGen[40]), 
          .A1(n13061), .B1(n3678), .C1(n8035), .D1(phase_inc_carrGen[41]), 
          .CIN(n10998), .COUT(n10999), .S0(n2840), .S1(n2839));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_43.INIT0 = 16'hd1e2;
    defparam add_749_43.INIT1 = 16'he4b1;
    defparam add_749_43.INJECT1_0 = "NO";
    defparam add_749_43.INJECT1_1 = "NO";
    CCU2D add_749_41 (.A0(n3634), .B0(n13061), .C0(n2324), .D0(phase_inc_carrGen[38]), 
          .A1(n3634), .B1(n13061), .C1(n2323), .D1(phase_inc_carrGen[39]), 
          .CIN(n10997), .COUT(n10998), .S0(n2842), .S1(n2841));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_41.INIT0 = 16'hd1e2;
    defparam add_749_41.INIT1 = 16'hd1e2;
    defparam add_749_41.INJECT1_0 = "NO";
    defparam add_749_41.INJECT1_1 = "NO";
    CCU2D add_749_39 (.A0(n7603), .B0(n13061), .C0(n2326), .D0(phase_inc_carrGen[36]), 
          .A1(n3682), .B1(n13061), .C1(n2325), .D1(phase_inc_carrGen[37]), 
          .CIN(n10996), .COUT(n10997), .S0(n2844), .S1(n2843));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_39.INIT0 = 16'hd1e2;
    defparam add_749_39.INIT1 = 16'hd1e2;
    defparam add_749_39.INJECT1_0 = "NO";
    defparam add_749_39.INJECT1_1 = "NO";
    CCU2D add_749_37 (.A0(n7603), .B0(n13061), .C0(n2328), .D0(phase_inc_carrGen[34]), 
          .A1(n13061), .B1(n7603), .C1(n2327), .D1(phase_inc_carrGen[35]), 
          .CIN(n10995), .COUT(n10996), .S0(n2846), .S1(n2845));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_37.INIT0 = 16'hd1e2;
    defparam add_749_37.INIT1 = 16'he4b1;
    defparam add_749_37.INJECT1_0 = "NO";
    defparam add_749_37.INJECT1_1 = "NO";
    CCU2D add_749_35 (.A0(n13061), .B0(n3678), .C0(n2330), .D0(phase_inc_carrGen[32]), 
          .A1(n7603), .B1(n13061), .C1(n2329), .D1(phase_inc_carrGen[33]), 
          .CIN(n10994), .COUT(n10995), .S0(n2848), .S1(n2847));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_35.INIT0 = 16'he4b1;
    defparam add_749_35.INIT1 = 16'hd1e2;
    defparam add_749_35.INJECT1_0 = "NO";
    defparam add_749_35.INJECT1_1 = "NO";
    CCU2D add_749_33 (.A0(n3653), .B0(n13061), .C0(n2332), .D0(phase_inc_carrGen[30]), 
          .A1(n3686), .B1(n13061), .C1(n2331), .D1(phase_inc_carrGen[31]), 
          .CIN(n10993), .COUT(n10994), .S0(n2850), .S1(n2849));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_33.INIT0 = 16'hd1e2;
    defparam add_749_33.INIT1 = 16'hd1e2;
    defparam add_749_33.INJECT1_0 = "NO";
    defparam add_749_33.INJECT1_1 = "NO";
    CCU2D add_749_31 (.A0(n3653), .B0(n13061), .C0(n2334), .D0(phase_inc_carrGen[28]), 
          .A1(n3678), .B1(n13061), .C1(n2333), .D1(phase_inc_carrGen[29]), 
          .CIN(n10992), .COUT(n10993), .S0(n2852), .S1(n2851));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_31.INIT0 = 16'hd1e2;
    defparam add_749_31.INIT1 = 16'hd1e2;
    defparam add_749_31.INJECT1_0 = "NO";
    defparam add_749_31.INJECT1_1 = "NO";
    CCU2D add_749_29 (.A0(n3634), .B0(n13061), .C0(n2336), .D0(phase_inc_carrGen[26]), 
          .A1(n7603), .B1(n13061), .C1(n2335), .D1(phase_inc_carrGen[27]), 
          .CIN(n10991), .COUT(n10992), .S0(n2854), .S1(n2853));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_29.INIT0 = 16'hd1e2;
    defparam add_749_29.INIT1 = 16'hd1e2;
    defparam add_749_29.INJECT1_0 = "NO";
    defparam add_749_29.INJECT1_1 = "NO";
    CCU2D add_749_27 (.A0(n3634), .B0(n13061), .C0(n2338), .D0(phase_inc_carrGen[24]), 
          .A1(n3634), .B1(n13061), .C1(n2337), .D1(phase_inc_carrGen[25]), 
          .CIN(n10990), .COUT(n10991), .S0(n2856), .S1(n2855));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_27.INIT0 = 16'hd1e2;
    defparam add_749_27.INIT1 = 16'hd1e2;
    defparam add_749_27.INJECT1_0 = "NO";
    defparam add_749_27.INJECT1_1 = "NO";
    CCU2D add_749_25 (.A0(n7603), .B0(n13061), .C0(n2340), .D0(phase_inc_carrGen[22]), 
          .A1(n3686), .B1(n13061), .C1(n2339), .D1(phase_inc_carrGen[23]), 
          .CIN(n10989), .COUT(n10990), .S0(n2858), .S1(n2857));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_25.INIT0 = 16'hd1e2;
    defparam add_749_25.INIT1 = 16'hd1e2;
    defparam add_749_25.INJECT1_0 = "NO";
    defparam add_749_25.INJECT1_1 = "NO";
    CCU2D add_749_23 (.A0(n13061), .B0(n7603), .C0(n2342), .D0(phase_inc_carrGen[20]), 
          .A1(n13061), .B1(n3678), .C1(n2341), .D1(phase_inc_carrGen[21]), 
          .CIN(n10988), .COUT(n10989), .S0(n2860), .S1(n2859));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_23.INIT0 = 16'he4b1;
    defparam add_749_23.INIT1 = 16'he4b1;
    defparam add_749_23.INJECT1_0 = "NO";
    defparam add_749_23.INJECT1_1 = "NO";
    CCU2D add_749_21 (.A0(n3678), .B0(n13061), .C0(n2344), .D0(phase_inc_carrGen[18]), 
          .A1(n3682), .B1(n13061), .C1(n8033), .D1(phase_inc_carrGen[19]), 
          .CIN(n10987), .COUT(n10988), .S0(n2862), .S1(n2861));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_21.INIT0 = 16'hd1e2;
    defparam add_749_21.INIT1 = 16'hd1e2;
    defparam add_749_21.INJECT1_0 = "NO";
    defparam add_749_21.INJECT1_1 = "NO";
    CCU2D add_749_19 (.A0(n3678), .B0(n13061), .C0(n2346), .D0(phase_inc_carrGen[16]), 
          .A1(n13061), .B1(n7603), .C1(n8031), .D1(phase_inc_carrGen[17]), 
          .CIN(n10986), .COUT(n10987), .S0(n2864), .S1(n2863));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_19.INIT0 = 16'hd1e2;
    defparam add_749_19.INIT1 = 16'he4b1;
    defparam add_749_19.INJECT1_0 = "NO";
    defparam add_749_19.INJECT1_1 = "NO";
    CCU2D add_749_17 (.A0(n3682), .B0(n13061), .C0(n2348), .D0(phase_inc_carrGen[14]), 
          .A1(n7603), .B1(n13061), .C1(n2347), .D1(phase_inc_carrGen[15]), 
          .CIN(n10985), .COUT(n10986), .S0(n2866), .S1(n2865));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_17.INIT0 = 16'hd1e2;
    defparam add_749_17.INIT1 = 16'hd1e2;
    defparam add_749_17.INJECT1_0 = "NO";
    defparam add_749_17.INJECT1_1 = "NO";
    CCU2D add_749_15 (.A0(n3682), .B0(n13061), .C0(n2350), .D0(phase_inc_carrGen[12]), 
          .A1(n3678), .B1(n13061), .C1(n8029), .D1(phase_inc_carrGen[13]), 
          .CIN(n10984), .COUT(n10985), .S0(n2868), .S1(n2867));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_15.INIT0 = 16'hd1e2;
    defparam add_749_15.INIT1 = 16'hd1e2;
    defparam add_749_15.INJECT1_0 = "NO";
    defparam add_749_15.INJECT1_1 = "NO";
    CCU2D add_749_13 (.A0(n3686), .B0(n13061), .C0(n2352), .D0(phase_inc_carrGen[10]), 
          .A1(n3634), .B1(n13061), .C1(n2351), .D1(phase_inc_carrGen[11]), 
          .CIN(n10983), .COUT(n10984), .S0(n2870), .S1(n2869));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_13.INIT0 = 16'hd1e2;
    defparam add_749_13.INIT1 = 16'hd1e2;
    defparam add_749_13.INJECT1_0 = "NO";
    defparam add_749_13.INJECT1_1 = "NO";
    CCU2D add_749_11 (.A0(n13061), .B0(n3678), .C0(n2354), .D0(phase_inc_carrGen[8]), 
          .A1(n3686), .B1(n13061), .C1(n2353), .D1(phase_inc_carrGen[9]), 
          .CIN(n10982), .COUT(n10983), .S0(n2872), .S1(n2871));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_11.INIT0 = 16'he4b1;
    defparam add_749_11.INIT1 = 16'hd1e2;
    defparam add_749_11.INJECT1_0 = "NO";
    defparam add_749_11.INJECT1_1 = "NO";
    CCU2D add_749_9 (.A0(n3682), .B0(n13061), .C0(n8027), .D0(phase_inc_carrGen[6]), 
          .A1(n3686), .B1(n13061), .C1(n2355), .D1(phase_inc_carrGen[7]), 
          .CIN(n10981), .COUT(n10982), .S0(n2874), .S1(n2873));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_9.INIT0 = 16'hd1e2;
    defparam add_749_9.INIT1 = 16'hd1e2;
    defparam add_749_9.INJECT1_0 = "NO";
    defparam add_749_9.INJECT1_1 = "NO";
    CCU2D add_749_7 (.A0(n7603), .B0(n13061), .C0(n2358), .D0(phase_inc_carrGen[4]), 
          .A1(n3682), .B1(n13061), .C1(n2357), .D1(phase_inc_carrGen[5]), 
          .CIN(n10980), .COUT(n10981), .S0(n2876), .S1(n2875));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_7.INIT0 = 16'hd1e2;
    defparam add_749_7.INIT1 = 16'hd1e2;
    defparam add_749_7.INJECT1_0 = "NO";
    defparam add_749_7.INJECT1_1 = "NO";
    CCU2D add_749_5 (.A0(n13061), .B0(n7603), .C0(n2360), .D0(phase_inc_carrGen[2]), 
          .A1(n3634), .B1(n13061), .C1(n2359), .D1(phase_inc_carrGen[3]), 
          .CIN(n10979), .COUT(n10980), .S0(n2878), .S1(n2877));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_5.INIT0 = 16'he4b1;
    defparam add_749_5.INIT1 = 16'hd1e2;
    defparam add_749_5.INJECT1_0 = "NO";
    defparam add_749_5.INJECT1_1 = "NO";
    CCU2D add_749_3 (.A0(n3678), .B0(n13061), .C0(n2628), .D0(phase_inc_carrGen[0]), 
          .A1(n3686), .B1(n13061), .C1(n2361), .D1(phase_inc_carrGen[1]), 
          .CIN(n10978), .COUT(n10979), .S0(n2880), .S1(n2879));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_3.INIT0 = 16'hd1e2;
    defparam add_749_3.INIT1 = 16'hd1e2;
    defparam add_749_3.INJECT1_0 = "NO";
    defparam add_749_3.INJECT1_1 = "NO";
    CCU2D add_749_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n3634), .B1(n13061), .C1(GND_net), .D1(GND_net), .COUT(n10978));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam add_749_1.INIT0 = 16'hF000;
    defparam add_749_1.INIT1 = 16'hdddd;
    defparam add_749_1.INJECT1_0 = "NO";
    defparam add_749_1.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_61 (.A0(phase_inc_carrGen[63]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n10836), .S0(n1031));
    defparam sub_45_add_2_61.INIT0 = 16'h5555;
    defparam sub_45_add_2_61.INIT1 = 16'h0000;
    defparam sub_45_add_2_61.INJECT1_0 = "NO";
    defparam sub_45_add_2_61.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_59 (.A0(phase_inc_carrGen[61]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[62]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10835), .COUT(n10836), .S0(n1033), .S1(n1032));
    defparam sub_45_add_2_59.INIT0 = 16'h5555;
    defparam sub_45_add_2_59.INIT1 = 16'h5555;
    defparam sub_45_add_2_59.INJECT1_0 = "NO";
    defparam sub_45_add_2_59.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_57 (.A0(phase_inc_carrGen[59]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[60]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10834), .COUT(n10835), .S0(n1035), .S1(n1034));
    defparam sub_45_add_2_57.INIT0 = 16'h5555;
    defparam sub_45_add_2_57.INIT1 = 16'h5555;
    defparam sub_45_add_2_57.INJECT1_0 = "NO";
    defparam sub_45_add_2_57.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_55 (.A0(phase_inc_carrGen[57]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[58]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10833), .COUT(n10834), .S0(n1037), .S1(n1036));
    defparam sub_45_add_2_55.INIT0 = 16'h5555;
    defparam sub_45_add_2_55.INIT1 = 16'h5555;
    defparam sub_45_add_2_55.INJECT1_0 = "NO";
    defparam sub_45_add_2_55.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_53 (.A0(phase_inc_carrGen[55]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[56]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10832), .COUT(n10833), .S0(n1039), .S1(n1038));
    defparam sub_45_add_2_53.INIT0 = 16'h5555;
    defparam sub_45_add_2_53.INIT1 = 16'h5555;
    defparam sub_45_add_2_53.INJECT1_0 = "NO";
    defparam sub_45_add_2_53.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_51 (.A0(phase_inc_carrGen[53]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[54]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10831), .COUT(n10832), .S0(n1041), .S1(n1040));
    defparam sub_45_add_2_51.INIT0 = 16'h5555;
    defparam sub_45_add_2_51.INIT1 = 16'h5555;
    defparam sub_45_add_2_51.INJECT1_0 = "NO";
    defparam sub_45_add_2_51.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_49 (.A0(phase_inc_carrGen[51]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[52]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10830), .COUT(n10831), .S0(n1043), .S1(n1042));
    defparam sub_45_add_2_49.INIT0 = 16'h5555;
    defparam sub_45_add_2_49.INIT1 = 16'h5555;
    defparam sub_45_add_2_49.INJECT1_0 = "NO";
    defparam sub_45_add_2_49.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_47 (.A0(phase_inc_carrGen[49]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[50]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10829), .COUT(n10830), .S0(n1045), .S1(n1044));
    defparam sub_45_add_2_47.INIT0 = 16'h5aaa;
    defparam sub_45_add_2_47.INIT1 = 16'h5aaa;
    defparam sub_45_add_2_47.INJECT1_0 = "NO";
    defparam sub_45_add_2_47.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_45 (.A0(phase_inc_carrGen[47]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[48]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10828), .COUT(n10829), .S0(n1047), .S1(n1046));
    defparam sub_45_add_2_45.INIT0 = 16'h5555;
    defparam sub_45_add_2_45.INIT1 = 16'h5aaa;
    defparam sub_45_add_2_45.INJECT1_0 = "NO";
    defparam sub_45_add_2_45.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_43 (.A0(phase_inc_carrGen[45]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[46]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10827), .COUT(n10828), .S0(n1049), .S1(n1048));
    defparam sub_45_add_2_43.INIT0 = 16'h5555;
    defparam sub_45_add_2_43.INIT1 = 16'h5555;
    defparam sub_45_add_2_43.INJECT1_0 = "NO";
    defparam sub_45_add_2_43.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_41 (.A0(phase_inc_carrGen[43]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[44]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10826), .COUT(n10827), .S0(n1051), .S1(n1050));
    defparam sub_45_add_2_41.INIT0 = 16'h5aaa;
    defparam sub_45_add_2_41.INIT1 = 16'h5aaa;
    defparam sub_45_add_2_41.INJECT1_0 = "NO";
    defparam sub_45_add_2_41.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_39 (.A0(phase_inc_carrGen[41]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[42]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10825), .COUT(n10826), .S0(n1053), .S1(n1052));
    defparam sub_45_add_2_39.INIT0 = 16'h5aaa;
    defparam sub_45_add_2_39.INIT1 = 16'h5555;
    defparam sub_45_add_2_39.INJECT1_0 = "NO";
    defparam sub_45_add_2_39.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_37 (.A0(phase_inc_carrGen[39]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[40]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10824), .COUT(n10825), .S0(n1055), .S1(n1054));
    defparam sub_45_add_2_37.INIT0 = 16'h5555;
    defparam sub_45_add_2_37.INIT1 = 16'h5aaa;
    defparam sub_45_add_2_37.INJECT1_0 = "NO";
    defparam sub_45_add_2_37.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_35 (.A0(phase_inc_carrGen[37]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[38]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10823), .COUT(n10824), .S0(n1057), .S1(n1056));
    defparam sub_45_add_2_35.INIT0 = 16'h5aaa;
    defparam sub_45_add_2_35.INIT1 = 16'h5555;
    defparam sub_45_add_2_35.INJECT1_0 = "NO";
    defparam sub_45_add_2_35.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_33 (.A0(phase_inc_carrGen[35]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[36]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10822), .COUT(n10823), .S0(n1059), .S1(n1058));
    defparam sub_45_add_2_33.INIT0 = 16'h5555;
    defparam sub_45_add_2_33.INIT1 = 16'h5aaa;
    defparam sub_45_add_2_33.INJECT1_0 = "NO";
    defparam sub_45_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_31 (.A0(phase_inc_carrGen[33]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[34]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10821), .COUT(n10822), .S0(n1061), .S1(n1060));
    defparam sub_45_add_2_31.INIT0 = 16'h5aaa;
    defparam sub_45_add_2_31.INIT1 = 16'h5aaa;
    defparam sub_45_add_2_31.INJECT1_0 = "NO";
    defparam sub_45_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_29 (.A0(phase_inc_carrGen[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[32]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10820), .COUT(n10821), .S0(n1063), .S1(n1062));
    defparam sub_45_add_2_29.INIT0 = 16'h5555;
    defparam sub_45_add_2_29.INIT1 = 16'h5aaa;
    defparam sub_45_add_2_29.INJECT1_0 = "NO";
    defparam sub_45_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_27 (.A0(phase_inc_carrGen[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10819), .COUT(n10820), .S0(n1065), .S1(n1064));
    defparam sub_45_add_2_27.INIT0 = 16'h5555;
    defparam sub_45_add_2_27.INIT1 = 16'h5aaa;
    defparam sub_45_add_2_27.INJECT1_0 = "NO";
    defparam sub_45_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_25 (.A0(phase_inc_carrGen[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10818), .COUT(n10819), .S0(n1067), .S1(n1066));
    defparam sub_45_add_2_25.INIT0 = 16'h5aaa;
    defparam sub_45_add_2_25.INIT1 = 16'h5aaa;
    defparam sub_45_add_2_25.INJECT1_0 = "NO";
    defparam sub_45_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_23 (.A0(phase_inc_carrGen[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10817), .COUT(n10818), .S0(n1069), .S1(n1068));
    defparam sub_45_add_2_23.INIT0 = 16'h5555;
    defparam sub_45_add_2_23.INIT1 = 16'h5555;
    defparam sub_45_add_2_23.INJECT1_0 = "NO";
    defparam sub_45_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_21 (.A0(phase_inc_carrGen[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10816), .COUT(n10817), .S0(n1071), .S1(n1070));
    defparam sub_45_add_2_21.INIT0 = 16'h5555;
    defparam sub_45_add_2_21.INIT1 = 16'h5555;
    defparam sub_45_add_2_21.INJECT1_0 = "NO";
    defparam sub_45_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_19 (.A0(phase_inc_carrGen[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10815), .COUT(n10816), .S0(n1073), .S1(n1072));
    defparam sub_45_add_2_19.INIT0 = 16'h5aaa;
    defparam sub_45_add_2_19.INIT1 = 16'h5aaa;
    defparam sub_45_add_2_19.INJECT1_0 = "NO";
    defparam sub_45_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_17 (.A0(phase_inc_carrGen[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10814), .COUT(n10815), .S0(n1075), .S1(n1074));
    defparam sub_45_add_2_17.INIT0 = 16'h5aaa;
    defparam sub_45_add_2_17.INIT1 = 16'h5555;
    defparam sub_45_add_2_17.INJECT1_0 = "NO";
    defparam sub_45_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_15 (.A0(phase_inc_carrGen[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10813), .COUT(n10814), .S0(n1077), .S1(n1076));
    defparam sub_45_add_2_15.INIT0 = 16'h5555;
    defparam sub_45_add_2_15.INIT1 = 16'h5555;
    defparam sub_45_add_2_15.INJECT1_0 = "NO";
    defparam sub_45_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_13 (.A0(phase_inc_carrGen[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10812), .COUT(n10813), .S0(n1079), .S1(n1078));
    defparam sub_45_add_2_13.INIT0 = 16'h5aaa;
    defparam sub_45_add_2_13.INIT1 = 16'h5555;
    defparam sub_45_add_2_13.INJECT1_0 = "NO";
    defparam sub_45_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_11 (.A0(phase_inc_carrGen[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10811), .COUT(n10812), .S0(n1081), .S1(n1080));
    defparam sub_45_add_2_11.INIT0 = 16'h5555;
    defparam sub_45_add_2_11.INIT1 = 16'h5aaa;
    defparam sub_45_add_2_11.INJECT1_0 = "NO";
    defparam sub_45_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_9 (.A0(phase_inc_carrGen[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10810), .COUT(n10811), .S0(n1083), .S1(n1082));
    defparam sub_45_add_2_9.INIT0 = 16'h5555;
    defparam sub_45_add_2_9.INIT1 = 16'h5aaa;
    defparam sub_45_add_2_9.INJECT1_0 = "NO";
    defparam sub_45_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_7 (.A0(phase_inc_carrGen[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10809), .COUT(n10810), .S0(n1085), .S1(n1084));
    defparam sub_45_add_2_7.INIT0 = 16'h5555;
    defparam sub_45_add_2_7.INIT1 = 16'h5555;
    defparam sub_45_add_2_7.INJECT1_0 = "NO";
    defparam sub_45_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_5 (.A0(phase_inc_carrGen[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10808), .COUT(n10809), .S0(n1087), .S1(n1086));
    defparam sub_45_add_2_5.INIT0 = 16'h5555;
    defparam sub_45_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_45_add_2_5.INJECT1_0 = "NO";
    defparam sub_45_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_3 (.A0(phase_inc_carrGen[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10807), .COUT(n10808), .S0(n1089), .S1(n1088));
    defparam sub_45_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_45_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_45_add_2_3.INJECT1_0 = "NO";
    defparam sub_45_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_45_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(phase_inc_carrGen[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n10807), .S1(n1090));
    defparam sub_45_add_2_1.INIT0 = 16'hF000;
    defparam sub_45_add_2_1.INIT1 = 16'h5555;
    defparam sub_45_add_2_1.INJECT1_0 = "NO";
    defparam sub_45_add_2_1.INJECT1_1 = "NO";
    LUT4 mux_322_i27_4_lut (.A(n7796), .B(n1129), .C(n13056), .D(n2563), 
         .Z(n2336)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i27_4_lut.init = 16'hc0ca;
    LUT4 i1_2_lut (.A(o_Rx_Byte[4]), .B(o_Rx_Byte[0]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(271[4] 285[10])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 mux_322_i28_4_lut (.A(n7798), .B(n1128), .C(n13056), .D(n2563), 
         .Z(n2335)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i28_4_lut.init = 16'hcfca;
    LUT4 i5367_3_lut_4_lut (.A(n13067), .B(n13054), .C(n13212), .D(o_Rx_Byte[3]), 
         .Z(osc_clk_enable_1411)) /* synthesis lut_function=(A (C)+!A !(B ((D)+!C)+!B !(C))) */ ;
    defparam i5367_3_lut_4_lut.init = 16'hb0f0;
    LUT4 i1813_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(n13179), 
         .D(n1035), .Z(n7854)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1813_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_322_i25_4_lut (.A(n7792), .B(n1131), .C(n13056), .D(n2563), 
         .Z(n2338)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i25_4_lut.init = 16'hc0ca;
    LUT4 i1805_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(n13179), 
         .D(n1040), .Z(n7846)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1805_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_322_i26_4_lut (.A(n7794), .B(n1130), .C(n13056), .D(n2563), 
         .Z(n2337)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i26_4_lut.init = 16'hc0ca;
    LUT4 i2665_3_lut_3_lut (.A(o_Rx_Byte[3]), .B(n13063), .C(n1072), .Z(n2540)) /* synthesis lut_function=(A (C)+!A !(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam i2665_3_lut_3_lut.init = 16'hb1b1;
    LUT4 mux_322_i23_4_lut (.A(n2540), .B(n1133), .C(n13056), .D(n2563), 
         .Z(n2340)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i23_4_lut.init = 16'hcfca;
    LUT4 i1793_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(n13179), 
         .D(n1047), .Z(n7834)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1793_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i2666_3_lut_3_lut (.A(n13179), .B(n13063), .C(n1054), .Z(n2522)) /* synthesis lut_function=(A (C)+!A !(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam i2666_3_lut_3_lut.init = 16'hb1b1;
    LUT4 mux_322_i24_4_lut (.A(n7790), .B(n1132), .C(n13056), .D(n2563), 
         .Z(n2339)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i24_4_lut.init = 16'hcfca;
    LUT4 i2663_3_lut_3_lut (.A(o_Rx_Byte[3]), .B(n13063), .C(n1082), .Z(n2550)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam i2663_3_lut_3_lut.init = 16'he4e4;
    LUT4 i2664_3_lut_3_lut (.A(o_Rx_Byte[3]), .B(n13063), .C(n1079), .Z(n2547)) /* synthesis lut_function=(A (C)+!A !(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam i2664_3_lut_3_lut.init = 16'hb1b1;
    LUT4 mux_322_i21_4_lut (.A(n7786), .B(n1135), .C(n13056), .D(n2563), 
         .Z(n2342)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i21_4_lut.init = 16'hcfca;
    LUT4 i2662_3_lut_3_lut (.A(o_Rx_Byte[3]), .B(n13063), .C(n1087), .Z(n2555)) /* synthesis lut_function=(A (C)+!A !(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam i2662_3_lut_3_lut.init = 16'hb1b1;
    LUT4 mux_322_i22_4_lut (.A(n2541), .B(n1134), .C(n13056), .D(n2563), 
         .Z(n2341)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i22_4_lut.init = 16'hcfca;
    LUT4 i1799_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(o_Rx_Byte[3]), 
         .D(n1043), .Z(n7840)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1799_3_lut_4_lut.init = 16'hf404;
    LUT4 i1789_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(n13179), 
         .D(n1049), .Z(n7830)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1789_3_lut_4_lut.init = 16'hf404;
    LUT4 i2726_2_lut (.A(n1073), .B(n13179), .Z(n2541)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i2726_2_lut.init = 16'h8888;
    LUT4 i1779_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(o_Rx_Byte[3]), 
         .D(n1056), .Z(n7820)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1779_3_lut_4_lut.init = 16'hf404;
    LUT4 mux_322_i19_4_lut (.A(n7782), .B(n1137), .C(n13056), .D(n2563), 
         .Z(n2344)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i19_4_lut.init = 16'hc0ca;
    LUT4 i1980_4_lut (.A(n1136), .B(n1075), .C(o_Rx_Byte[3]), .D(n13060), 
         .Z(n8033)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1980_4_lut.init = 16'hcac0;
    LUT4 mux_322_i17_4_lut (.A(n7778), .B(n1139), .C(n13056), .D(n2563), 
         .Z(n2346)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i17_4_lut.init = 16'hcfca;
    LUT4 i1781_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(n13179), 
         .D(n1055), .Z(n7822)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1781_3_lut_4_lut.init = 16'hf404;
    LUT4 i1775_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(n13179), 
         .D(n1058), .Z(n7816)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1775_3_lut_4_lut.init = 16'hf404;
    LUT4 i1773_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(o_Rx_Byte[3]), 
         .D(n1059), .Z(n7814)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1773_3_lut_4_lut.init = 16'hf404;
    LUT4 o_Rx_Byte_4__bdd_4_lut_5399 (.A(o_Rx_Byte[4]), .B(o_Rx_Byte[2]), 
         .C(o_Rx_Byte[3]), .D(o_Rx_Byte[0]), .Z(n12946)) /* synthesis lut_function=(!(A+(B (C (D))+!B (C+(D))))) */ ;
    defparam o_Rx_Byte_4__bdd_4_lut_5399.init = 16'h0445;
    LUT4 i1_2_lut_rep_86 (.A(o_Rx_Byte[4]), .B(n12533), .Z(n13060)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(271[4] 285[10])
    defparam i1_2_lut_rep_86.init = 16'h8888;
    LUT4 i1978_4_lut (.A(n1138), .B(n1077), .C(o_Rx_Byte[3]), .D(n13060), 
         .Z(n8031)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1978_4_lut.init = 16'hcac0;
    LUT4 i1791_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(o_Rx_Byte[3]), 
         .D(n1048), .Z(n7832)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1791_3_lut_4_lut.init = 16'hf707;
    LUT4 i1_4_lut_adj_60 (.A(n8257), .B(o_Rx_Byte[2]), .C(o_Rx_Byte[0]), 
         .D(MYLED_c_6), .Z(n12533)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(271[4] 285[10])
    defparam i1_4_lut_adj_60.init = 16'h0020;
    LUT4 i1_4_lut_adj_61 (.A(o_Rx_Byte[5]), .B(o_Rx_Byte[7]), .C(o_Rx_Byte[6]), 
         .D(o_Rx_DV), .Z(n8257)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam i1_4_lut_adj_61.init = 16'h2000;
    LUT4 i1785_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(o_Rx_Byte[3]), 
         .D(n1052), .Z(n7826)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1785_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_322_i56_4_lut (.A(n2373), .B(n1100), .C(n13056), .D(n7997), 
         .Z(n2307)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i56_4_lut.init = 16'hcfca;
    LUT4 mux_322_i3_4_lut_4_lut_4_lut (.A(o_Rx_Byte[3]), .B(o_Rx_Byte[4]), 
         .C(n12533), .D(n1153), .Z(n2360)) /* synthesis lut_function=(!(A+!(B ((D)+!C)+!B !(C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam mux_322_i3_4_lut_4_lut_4_lut.init = 16'h4505;
    LUT4 i1745_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(o_Rx_Byte[3]), 
         .D(n1074), .Z(n7786)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1745_3_lut_4_lut.init = 16'hf707;
    LUT4 i1735_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(n13179), 
         .D(n1080), .Z(n7776)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1735_3_lut_4_lut.init = 16'hf808;
    LUT4 i1725_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(n13179), 
         .D(n1086), .Z(n7766)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1725_3_lut_4_lut.init = 16'hf808;
    LUT4 i2674_2_lut (.A(n1039), .B(o_Rx_Byte[3]), .Z(n2373)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i2674_2_lut.init = 16'h8888;
    LUT4 i1727_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(o_Rx_Byte[3]), 
         .D(n1085), .Z(n7768)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1727_3_lut_4_lut.init = 16'hf707;
    LUT4 i1984_4_lut (.A(n1103), .B(n1042), .C(o_Rx_Byte[3]), .D(n13060), 
         .Z(n8037)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1984_4_lut.init = 16'hcac0;
    LUT4 i1721_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(o_Rx_Byte[3]), 
         .D(n1089), .Z(n7762)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1721_3_lut_4_lut.init = 16'hf808;
    LUT4 n12954_bdd_4_lut (.A(n12954), .B(n12953), .C(o_Rx_Byte[2]), .D(n8257), 
         .Z(n2815)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n12954_bdd_4_lut.init = 16'hca00;
    LUT4 PWMOut_I_0_1_lut (.A(PWMOutP4_c), .Z(PWMOutN4_c)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(135[19:26])
    defparam PWMOut_I_0_1_lut.init = 16'h5555;
    LUT4 mux_322_i4_3_lut_4_lut (.A(o_Rx_Byte[3]), .B(n13060), .C(n1152), 
         .D(n2628), .Z(n2359)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam mux_322_i4_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1988_4_lut (.A(n1093), .B(n1032), .C(o_Rx_Byte[3]), .D(n13060), 
         .Z(n8041)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1988_4_lut.init = 16'hcac0;
    LUT4 mux_322_i54_4_lut (.A(n7844), .B(n1102), .C(n13056), .D(n2563), 
         .Z(n2309)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i54_4_lut.init = 16'hc0ca;
    LUT4 i345_2_lut_rep_82_3_lut (.A(o_Rx_Byte[4]), .B(n12533), .C(n13179), 
         .Z(n13056)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(271[4] 285[10])
    defparam i345_2_lut_rep_82_3_lut.init = 16'h0808;
    LUT4 i1990_4_lut (.A(n1092), .B(n1031), .C(o_Rx_Byte[3]), .D(n13060), 
         .Z(n8043)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1990_4_lut.init = 16'hcac0;
    LUT4 i1777_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(o_Rx_Byte[3]), 
         .D(n1057), .Z(n7818)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1777_3_lut_4_lut.init = 16'hf707;
    LUT4 mux_322_i61_4_lut (.A(n7856), .B(n1095), .C(n13056), .D(n2563), 
         .Z(n2302)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i61_4_lut.init = 16'hc0ca;
    Mixer Mixer1 (.MixerOutSin({MixerOutSin}), .osc_clk(osc_clk), .DiffOut_c(DiffOut_c), 
          .MixerOutCos({MixerOutCos}), .RFIn_c(RFIn_c), .\LOCosine[12] (LOCosine[12]), 
          .GND_net(GND_net), .\LOCosine[10] (LOCosine[10]), .\LOCosine[11] (LOCosine[11]), 
          .\LOCosine[8] (LOCosine[8]), .\LOCosine[9] (LOCosine[9]), .\LOCosine[6] (LOCosine[6]), 
          .\LOCosine[7] (LOCosine[7]), .\LOCosine[4] (LOCosine[4]), .\LOCosine[5] (LOCosine[5]), 
          .\LOCosine[2] (LOCosine[2]), .\LOCosine[3] (LOCosine[3]), .\LOCosine[1] (LOCosine[1]), 
          .\LOSine[12] (LOSine[12]), .\LOSine[10] (LOSine[10]), .\LOSine[11] (LOSine[11]), 
          .\LOSine[8] (LOSine[8]), .\LOSine[9] (LOSine[9]), .\LOSine[6] (LOSine[6]), 
          .\LOSine[7] (LOSine[7]), .\LOSine[4] (LOSine[4]), .\LOSine[5] (LOSine[5]), 
          .\LOSine[2] (LOSine[2]), .\LOSine[3] (LOSine[3]), .\LOSine[1] (LOSine[1])) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(160[7] 168[2])
    LUT4 i1986_4_lut (.A(n1094), .B(n1033), .C(o_Rx_Byte[3]), .D(n13060), 
         .Z(n8039)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1986_4_lut.init = 16'hcac0;
    FD1S3AX o_Rx_Byte_i3_rep_98 (.D(o_Rx_Byte1[3]), .CK(osc_clk), .Q(n13179));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam o_Rx_Byte_i3_rep_98.GSR = "ENABLED";
    LUT4 i1771_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(n13179), 
         .D(n1060), .Z(n7812)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1771_3_lut_4_lut.init = 16'hf808;
    LUT4 i1763_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(o_Rx_Byte[3]), 
         .D(n1064), .Z(n7804)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1763_3_lut_4_lut.init = 16'hf808;
    LUT4 i1755_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(o_Rx_Byte[3]), 
         .D(n1068), .Z(n7796)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1755_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_322_i59_4_lut (.A(n7852), .B(n1097), .C(n13056), .D(n2563), 
         .Z(n2304)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i59_4_lut.init = 16'hc0ca;
    LUT4 i1757_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(n13179), 
         .D(n1067), .Z(n7798)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1757_3_lut_4_lut.init = 16'hf707;
    LUT4 mux_322_i60_4_lut (.A(n7854), .B(n1096), .C(n13056), .D(n2563), 
         .Z(n2303)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i60_4_lut.init = 16'hc0ca;
    LUT4 i1753_3_lut_4_lut (.A(o_Rx_Byte[2]), .B(n13063), .C(n13179), 
         .D(n1069), .Z(n7794)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i1753_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_322_i57_4_lut (.A(n2506), .B(n1099), .C(n13056), .D(n2563), 
         .Z(n2306)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i57_4_lut.init = 16'hc0ca;
    LUT4 i2734_2_lut (.A(n1038), .B(o_Rx_Byte[3]), .Z(n2506)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i2734_2_lut.init = 16'hbbbb;
    LUT4 mux_322_i58_4_lut (.A(n2505), .B(n1098), .C(n13056), .D(n2563), 
         .Z(n2305)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i58_4_lut.init = 16'hcfca;
    LUT4 i2735_2_lut (.A(n1037), .B(o_Rx_Byte[3]), .Z(n2505)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i2735_2_lut.init = 16'h8888;
    FD1S3AX o_Rx_Byte_i0 (.D(o_Rx_Byte1[0]), .CK(osc_clk), .Q(o_Rx_Byte[0]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam o_Rx_Byte_i0.GSR = "ENABLED";
    LUT4 mux_322_i55_4_lut (.A(n7846), .B(n1101), .C(n13056), .D(n2563), 
         .Z(n2308)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i55_4_lut.init = 16'hcfca;
    LUT4 i5381_4_lut (.A(o_Rx_Byte[3]), .B(o_Rx_Byte[2]), .C(o_Rx_Byte[6]), 
         .D(n6), .Z(osc_clk_enable_1407)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i5381_4_lut.init = 16'h0001;
    LUT4 i2589_2_lut (.A(o_Rx_Byte[4]), .B(n2815), .Z(n3678)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i2589_2_lut.init = 16'h8888;
    FD1P3AX phase_inc_carrGen_i0_i2 (.D(n2878), .SP(osc_clk_enable_1411), 
            .CK(osc_clk), .Q(phase_inc_carrGen[2]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i2.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i3 (.D(n2877), .SP(osc_clk_enable_1411), 
            .CK(osc_clk), .Q(phase_inc_carrGen[3]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i3.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i4 (.D(n2876), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[4]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i4.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i5 (.D(n2875), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[5]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i5.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i6 (.D(n2874), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[6]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i6.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i7 (.D(n2873), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[7]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i7.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i8 (.D(n2872), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[8]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i8.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i9 (.D(n2871), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[9]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i9.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i10 (.D(n2870), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[10]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i10.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i11 (.D(n2869), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[11]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i11.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i12 (.D(n2868), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[12]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i12.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i13 (.D(n2867), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[13]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i13.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i14 (.D(n2866), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[14]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i14.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i15 (.D(n2865), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[15]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i15.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i16 (.D(n2864), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[16]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i16.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i17 (.D(n2863), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[17]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i17.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i18 (.D(n2862), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[18]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i18.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i19 (.D(n2861), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[19]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i19.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i20 (.D(n2860), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[20]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i20.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i21 (.D(n2859), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[21]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i21.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i22 (.D(n2858), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[22]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i22.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i23 (.D(n2857), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[23]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i23.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i24 (.D(n2856), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[24]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i24.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i25 (.D(n2855), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[25]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i25.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i26 (.D(n2854), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[26]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i26.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i27 (.D(n2853), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[27]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i27.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i28 (.D(n2852), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[28]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i28.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i29 (.D(n2851), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[29]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i29.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i30 (.D(n2850), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[30]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i30.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i31 (.D(n2849), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[31]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i31.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i32 (.D(n2848), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[32]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i32.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i33 (.D(n2847), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[33]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i33.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i34 (.D(n2846), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[34]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i34.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i35 (.D(n2845), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[35]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i35.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i36 (.D(n2844), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[36]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i36.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i37 (.D(n2843), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[37]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i37.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i38 (.D(n2842), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[38]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i38.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i39 (.D(n2841), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[39]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i39.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i40 (.D(n2840), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[40]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i40.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i41 (.D(n2839), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[41]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i41.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i42 (.D(n2838), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[42]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i42.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i43 (.D(n2837), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[43]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i43.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i44 (.D(n2836), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[44]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i44.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i45 (.D(n2835), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[45]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i45.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i46 (.D(n2834), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[46]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i46.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i47 (.D(n2833), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[47]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i47.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i48 (.D(n2832), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[48]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i48.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i49 (.D(n2831), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[49]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i49.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i50 (.D(n2830), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[50]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i50.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i51 (.D(n2829), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[51]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i51.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i52 (.D(n2828), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[52]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i52.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i53 (.D(n2827), .SP(osc_clk_enable_1461), 
            .CK(osc_clk), .Q(phase_inc_carrGen[53]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i53.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i54 (.D(n2826), .SP(osc_clk_enable_1471), 
            .CK(osc_clk), .Q(phase_inc_carrGen[54]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i54.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i55 (.D(n2825), .SP(osc_clk_enable_1471), 
            .CK(osc_clk), .Q(phase_inc_carrGen[55]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i55.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i56 (.D(n2824), .SP(osc_clk_enable_1471), 
            .CK(osc_clk), .Q(phase_inc_carrGen[56]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i56.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i57 (.D(n2823), .SP(osc_clk_enable_1471), 
            .CK(osc_clk), .Q(phase_inc_carrGen[57]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i57.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i58 (.D(n2822), .SP(osc_clk_enable_1471), 
            .CK(osc_clk), .Q(phase_inc_carrGen[58]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i58.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i59 (.D(n2821), .SP(osc_clk_enable_1471), 
            .CK(osc_clk), .Q(phase_inc_carrGen[59]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i59.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i60 (.D(n2820), .SP(osc_clk_enable_1471), 
            .CK(osc_clk), .Q(phase_inc_carrGen[60]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i60.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i61 (.D(n2819), .SP(osc_clk_enable_1471), 
            .CK(osc_clk), .Q(phase_inc_carrGen[61]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i61.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i62 (.D(n2818), .SP(osc_clk_enable_1471), 
            .CK(osc_clk), .Q(phase_inc_carrGen[62]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i62.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i63 (.D(n2817), .SP(osc_clk_enable_1471), 
            .CK(osc_clk), .Q(phase_inc_carrGen[63]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam phase_inc_carrGen_i0_i63.GSR = "ENABLED";
    VLO i1 (.Z(GND_net));
    TSALL TSALL_INST (.TSALL(GND_net));
    LUT4 mux_322_i51_4_lut (.A(n2512), .B(n1105), .C(n13056), .D(n2563), 
         .Z(n2312)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i51_4_lut.init = 16'hcfca;
    PFUMX i5446 (.BLUT(n13092), .ALUT(n13093), .C0(o_Rx_Byte[0]), .Z(n13094));
    LUT4 i2729_2_lut (.A(n1044), .B(n13179), .Z(n2512)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i2729_2_lut.init = 16'h8888;
    LUT4 mux_747_i3_3_lut (.A(o_Rx_Byte[2]), .B(o_Rx_Byte[4]), .C(n2815), 
         .Z(n7603)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_747_i3_3_lut.init = 16'hcaca;
    LUT4 mux_322_i52_4_lut (.A(n7840), .B(n1104), .C(n13056), .D(n2563), 
         .Z(n2311)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i52_4_lut.init = 16'hc0ca;
    LUT4 i2338_2_lut_4_lut_4_lut (.A(o_Rx_Byte[4]), .B(n13179), .C(n13068), 
         .D(n8257), .Z(n8391)) /* synthesis lut_function=(A (B)+!A (B+(C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam i2338_2_lut_4_lut_4_lut.init = 16'hdccc;
    LUT4 i356_2_lut_3_lut_3_lut (.A(o_Rx_Byte[4]), .B(o_Rx_Byte[3]), .C(n12533), 
         .Z(n2563)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam i356_2_lut_3_lut_3_lut.init = 16'h1010;
    SinCos SinCos1 (.osc_clk(osc_clk), .VCC_net(VCC_net), .GND_net(GND_net), 
           .\phase_accum[57] (phase_accum[57]), .\phase_accum[58] (phase_accum[58]), 
           .\phase_accum[59] (phase_accum[59]), .\phase_accum[60] (phase_accum[60]), 
           .\phase_accum[61] (phase_accum[61]), .\phase_accum[62] (phase_accum[62]), 
           .\phase_accum[63] (phase_accum[63]), .\LOSine[1] (LOSine[1]), 
           .\LOSine[2] (LOSine[2]), .\LOSine[3] (LOSine[3]), .\LOSine[4] (LOSine[4]), 
           .\LOSine[5] (LOSine[5]), .\LOSine[6] (LOSine[6]), .\LOSine[7] (LOSine[7]), 
           .\LOSine[8] (LOSine[8]), .\LOSine[9] (LOSine[9]), .\LOSine[10] (LOSine[10]), 
           .\LOSine[11] (LOSine[11]), .\LOSine[12] (LOSine[12]), .\LOCosine[1] (LOCosine[1]), 
           .\LOCosine[2] (LOCosine[2]), .\LOCosine[3] (LOCosine[3]), .\LOCosine[4] (LOCosine[4]), 
           .\LOCosine[5] (LOCosine[5]), .\LOCosine[6] (LOCosine[6]), .\LOCosine[7] (LOCosine[7]), 
           .\LOCosine[8] (LOCosine[8]), .\LOCosine[9] (LOCosine[9]), .\LOCosine[10] (LOCosine[10]), 
           .\LOCosine[11] (LOCosine[11]), .\LOCosine[12] (LOCosine[12]), 
           .\phase_accum[56] (phase_accum[56])) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    \CIC(width=72,decimation_ratio=4096)  CIC1Sin (.MixerOutSin({MixerOutSin}), 
            .osc_clk(osc_clk), .GND_net(GND_net), .CIC1_out_clkSin(CIC1_out_clkSin), 
            .\CIC1_outSin[0] (CIC1_outSin[0]), .\CICGain[0] (CICGain[0]), 
            .\CICGain[1] (CICGain[1]), .n62(n62), .\d10[60] (d10_adj_2554[60]), 
            .n63(n63), .\d_out_11__N_1819[2] (d_out_11__N_1819_adj_2579[2]), 
            .n64(n64), .\d_out_11__N_1819[3] (d_out_11__N_1819_adj_2579[3]), 
            .n65(n65), .\d_out_11__N_1819[4] (d_out_11__N_1819_adj_2579[4]), 
            .n66(n66), .\d_out_11__N_1819[5] (d_out_11__N_1819_adj_2579[5]), 
            .n67(n67), .\d_out_11__N_1819[6] (d_out_11__N_1819_adj_2579[6]), 
            .n68(n68), .\d_out_11__N_1819[7] (d_out_11__N_1819_adj_2579[7]), 
            .\d10[68] (d10_adj_2554[68]), .\d_out_11__N_1819[8] (d_out_11__N_1819_adj_2579[8]), 
            .n70(n70), .\d_out_11__N_1819[9] (d_out_11__N_1819_adj_2579[9]), 
            .\d10[71] (d10_adj_2554[71]), .\d_out_11__N_1819[11] (d_out_11__N_1819_adj_2579[11]), 
            .\CIC1_outSin[1] (CIC1_outSin[1]), .\CIC1_outSin[2] (CIC1_outSin[2]), 
            .\CIC1_outSin[3] (CIC1_outSin[3]), .\CIC1_outSin[4] (CIC1_outSin[4]), 
            .\CIC1_outSin[5] (CIC1_outSin[5]), .MYLED_c_0(MYLED_c_0), .MYLED_c_1(MYLED_c_1), 
            .MYLED_c_2(MYLED_c_2), .MYLED_c_3(MYLED_c_3), .MYLED_c_4(MYLED_c_4), 
            .MYLED_c_5(MYLED_c_5), .\d10[67] (d10_adj_2554[67]), .\d10[69] (d10_adj_2554[69]), 
            .\d10[70] (d10_adj_2554[70]), .\d10[65] (d10_adj_2554[65]), 
            .\d10[66] (d10_adj_2554[66]), .\d10[63] (d10_adj_2554[63]), 
            .\d_out_11__N_1819[10] (d_out_11__N_1819_adj_2579[10]), .\d10[64] (d10_adj_2554[64]), 
            .\d10[61] (d10_adj_2554[61]), .\d10[62] (d10_adj_2554[62]), 
            .n61(n61), .\d10[59] (d10_adj_2554[59])) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(171[45] 177[2])
    LUT4 i2580_2_lut_2_lut (.A(o_Rx_Byte[4]), .B(n2815), .Z(n3634)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam i2580_2_lut_2_lut.init = 16'h4444;
    LUT4 n2644_bdd_4_lut_5390_4_lut (.A(o_Rx_Byte[4]), .B(o_Rx_Byte[3]), 
         .C(MYLED_c_6), .D(o_Rx_Byte[0]), .Z(n12953)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam n2644_bdd_4_lut_5390_4_lut.init = 16'h4000;
    LUT4 i1949_3_lut_4_lut_4_lut (.A(o_Rx_Byte[4]), .B(o_Rx_Byte[3]), .C(n13063), 
         .D(n12533), .Z(n7997)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+(D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam i1949_3_lut_4_lut_4_lut.init = 16'h3130;
    LUT4 i1_4_lut_4_lut_then_4_lut (.A(o_Rx_Byte[4]), .B(o_Rx_Byte[3]), 
         .C(MYLED_c_6), .D(o_Rx_Byte[2]), .Z(n13093)) /* synthesis lut_function=(!(A+!(B (D)+!B (C (D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam i1_4_lut_4_lut_then_4_lut.init = 16'h5400;
    LUT4 mux_322_i49_4_lut (.A(n7836), .B(n1107), .C(n13056), .D(n2563), 
         .Z(n2314)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i49_4_lut.init = 16'hc0ca;
    LUT4 mux_747_i29_3_lut_3_lut (.A(o_Rx_Byte[4]), .B(n2815), .C(o_Rx_Byte[2]), 
         .Z(n3653)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam mux_747_i29_3_lut_3_lut.init = 16'h7474;
    LUT4 i1_4_lut_4_lut_else_4_lut (.A(o_Rx_Byte[4]), .B(o_Rx_Byte[3]), 
         .C(MYLED_c_6), .D(o_Rx_Byte[2]), .Z(n13092)) /* synthesis lut_function=(!(A+!(B (C (D))+!B (C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(238[8] 288[4])
    defparam i1_4_lut_4_lut_else_4_lut.init = 16'h5010;
    LUT4 mux_322_i50_4_lut (.A(n2379), .B(n1106), .C(n13056), .D(n7997), 
         .Z(n2313)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i50_4_lut.init = 16'hcfca;
    LUT4 i2673_2_lut (.A(n1045), .B(n13179), .Z(n2379)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i2673_2_lut.init = 16'h8888;
    GSR GSR_INST (.GSR(VCC_net));
    LUT4 mux_322_i47_4_lut (.A(n7832), .B(n1109), .C(n13056), .D(n2563), 
         .Z(n2316)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i47_4_lut.init = 16'hc0ca;
    LUT4 mux_322_i48_4_lut (.A(n7834), .B(n1108), .C(n13056), .D(n2563), 
         .Z(n2315)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i48_4_lut.init = 16'hcfca;
    LUT4 mux_322_i45_4_lut (.A(n2384), .B(n1111), .C(n13056), .D(n7997), 
         .Z(n2318)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i45_4_lut.init = 16'hc0ca;
    LUT4 i2672_2_lut (.A(n1050), .B(o_Rx_Byte[3]), .Z(n2384)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam i2672_2_lut.init = 16'hbbbb;
    LUT4 mux_322_i46_4_lut (.A(n7830), .B(n1110), .C(n13056), .D(n2563), 
         .Z(n2317)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(245[2] 287[6])
    defparam mux_322_i46_4_lut.init = 16'hcfca;
    nco_sig ncoGen (.osc_clk(osc_clk), .\phase_accum[56] (phase_accum[56]), 
            .\phase_accum[57] (phase_accum[57]), .\phase_accum[58] (phase_accum[58]), 
            .\phase_accum[59] (phase_accum[59]), .\phase_accum[60] (phase_accum[60]), 
            .\phase_accum[61] (phase_accum[61]), .\phase_accum[62] (phase_accum[62]), 
            .\phase_accum[63] (phase_accum[63]), .phase_inc_carrGen1({phase_inc_carrGen1}), 
            .GND_net(GND_net), .sinGen_c(sinGen_c)) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(151[10] 157[2])
    \CIC(width=72,decimation_ratio=4096)_U1  CIC1Cos (.GND_net(GND_net), .MixerOutCos({MixerOutCos}), 
            .osc_clk(osc_clk), .CIC1_outCos({CIC1_outCos}), .\d10[61] (d10_adj_2554[61]), 
            .\d10[62] (d10_adj_2554[62]), .\CICGain[0] (CICGain[0]), .n62(n62), 
            .\d10[63] (d10_adj_2554[63]), .n63(n63), .\d10[64] (d10_adj_2554[64]), 
            .n64(n64), .\d10[65] (d10_adj_2554[65]), .n65(n65), .\d10[66] (d10_adj_2554[66]), 
            .n66(n66), .\d10[60] (d10_adj_2554[60]), .n61(n61), .\d10[67] (d10_adj_2554[67]), 
            .n67(n67), .\d10[68] (d10_adj_2554[68]), .n68(n68), .\d10[69] (d10_adj_2554[69]), 
            .\d10[70] (d10_adj_2554[70]), .n70(n70), .\d10[59] (d10_adj_2554[59]), 
            .\d10[71] (d10_adj_2554[71]), .\d_out_11__N_1819[2] (d_out_11__N_1819_adj_2579[2]), 
            .\d_out_11__N_1819[3] (d_out_11__N_1819_adj_2579[3]), .\d_out_11__N_1819[4] (d_out_11__N_1819_adj_2579[4]), 
            .\d_out_11__N_1819[5] (d_out_11__N_1819_adj_2579[5]), .\d_out_11__N_1819[6] (d_out_11__N_1819_adj_2579[6]), 
            .\d_out_11__N_1819[7] (d_out_11__N_1819_adj_2579[7]), .\d_out_11__N_1819[8] (d_out_11__N_1819_adj_2579[8]), 
            .\d_out_11__N_1819[9] (d_out_11__N_1819_adj_2579[9]), .\d_out_11__N_1819[10] (d_out_11__N_1819_adj_2579[10]), 
            .\d_out_11__N_1819[11] (d_out_11__N_1819_adj_2579[11]), .\CICGain[1] (CICGain[1])) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(180[45] 186[2])
    AMDemodulator AMDemodulator1 (.CIC1_out_clkSin(CIC1_out_clkSin), .\CIC1_outSin[0] (CIC1_outSin[0]), 
            .CIC1_outCos({CIC1_outCos}), .\DataInReg_11__N_1856[0] (DataInReg_11__N_1856[0]), 
            .GND_net(GND_net), .\CIC1_outSin[1] (CIC1_outSin[1]), .\CIC1_outSin[2] (CIC1_outSin[2]), 
            .\CIC1_outSin[3] (CIC1_outSin[3]), .\CIC1_outSin[4] (CIC1_outSin[4]), 
            .\CIC1_outSin[5] (CIC1_outSin[5]), .MYLED_c_0(MYLED_c_0), .MYLED_c_1(MYLED_c_1), 
            .MYLED_c_2(MYLED_c_2), .MYLED_c_3(MYLED_c_3), .MYLED_c_4(MYLED_c_4), 
            .MYLED_c_5(MYLED_c_5), .\DataInReg_11__N_1856[1] (DataInReg_11__N_1856[1]), 
            .\DataInReg_11__N_1856[2] (DataInReg_11__N_1856[2]), .\DataInReg_11__N_1856[3] (DataInReg_11__N_1856[3]), 
            .\DataInReg_11__N_1856[4] (DataInReg_11__N_1856[4]), .\DataInReg_11__N_1856[5] (DataInReg_11__N_1856[5]), 
            .\DataInReg_11__N_1856[6] (DataInReg_11__N_1856[6]), .\DataInReg_11__N_1856[7] (DataInReg_11__N_1856[7]), 
            .\DataInReg_11__N_1856[8] (DataInReg_11__N_1856[8]), .\DemodOut[9] (DemodOut[9]), 
            .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(212[15] 217[10])
    
endmodule
//
// Verilog Description of module PWM
//

module PWM (osc_clk, \DataInReg_11__N_1856[0] , PWMOutP4_c, GND_net, 
            \DemodOut[9] , \DataInReg_11__N_1856[1] , \DataInReg_11__N_1856[2] , 
            \DataInReg_11__N_1856[3] , \DataInReg_11__N_1856[4] , \DataInReg_11__N_1856[5] , 
            \DataInReg_11__N_1856[6] , \DataInReg_11__N_1856[7] , \DataInReg_11__N_1856[8] ) /* synthesis syn_module_defined=1 */ ;
    input osc_clk;
    input \DataInReg_11__N_1856[0] ;
    output PWMOutP4_c;
    input GND_net;
    input \DemodOut[9] ;
    input \DataInReg_11__N_1856[1] ;
    input \DataInReg_11__N_1856[2] ;
    input \DataInReg_11__N_1856[3] ;
    input \DataInReg_11__N_1856[4] ;
    input \DataInReg_11__N_1856[5] ;
    input \DataInReg_11__N_1856[6] ;
    input \DataInReg_11__N_1856[7] ;
    input \DataInReg_11__N_1856[8] ;
    
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(69[8:15])
    wire [9:0]counter;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(7[11:18])
    wire [9:0]n45;
    wire [11:0]DataInReg;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(10[12:21])
    
    wire osc_clk_enable_1406, PWMOut_N_1869, n17, n15, n11, n12, 
        n11509, n11508, n11507, n11506, n11505;
    wire [11:0]n3949;
    
    wire n10974, n10973, n10972, n10971, n10970;
    
    FD1S3AX counter_1006__i0 (.D(n45[0]), .CK(osc_clk), .Q(counter[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_1006__i0.GSR = "ENABLED";
    FD1P3AX DataInReg__i1 (.D(\DataInReg_11__N_1856[0] ), .SP(osc_clk_enable_1406), 
            .CK(osc_clk), .Q(DataInReg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=189, LSE_RLINE=195 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i1.GSR = "ENABLED";
    FD1S3AX PWMOut_15 (.D(PWMOut_N_1869), .CK(osc_clk), .Q(PWMOutP4_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=189, LSE_RLINE=195 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam PWMOut_15.GSR = "ENABLED";
    LUT4 i5384_4_lut (.A(n17), .B(n15), .C(n11), .D(n12), .Z(osc_clk_enable_1406)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(26[7:19])
    defparam i5384_4_lut.init = 16'h0001;
    LUT4 i7_4_lut (.A(counter[1]), .B(counter[4]), .C(counter[6]), .D(counter[8]), 
         .Z(n17)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(26[7:19])
    defparam i7_4_lut.init = 16'hfffe;
    CCU2D counter_1006_add_4_11 (.A0(counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11509), .S0(n45[9]));   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_1006_add_4_11.INIT0 = 16'hfaaa;
    defparam counter_1006_add_4_11.INIT1 = 16'h0000;
    defparam counter_1006_add_4_11.INJECT1_0 = "NO";
    defparam counter_1006_add_4_11.INJECT1_1 = "NO";
    CCU2D counter_1006_add_4_9 (.A0(counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11508), .COUT(n11509), .S0(n45[7]), .S1(n45[8]));   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_1006_add_4_9.INIT0 = 16'hfaaa;
    defparam counter_1006_add_4_9.INIT1 = 16'hfaaa;
    defparam counter_1006_add_4_9.INJECT1_0 = "NO";
    defparam counter_1006_add_4_9.INJECT1_1 = "NO";
    CCU2D counter_1006_add_4_7 (.A0(counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11507), .COUT(n11508), .S0(n45[5]), .S1(n45[6]));   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_1006_add_4_7.INIT0 = 16'hfaaa;
    defparam counter_1006_add_4_7.INIT1 = 16'hfaaa;
    defparam counter_1006_add_4_7.INJECT1_0 = "NO";
    defparam counter_1006_add_4_7.INJECT1_1 = "NO";
    CCU2D counter_1006_add_4_5 (.A0(counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11506), .COUT(n11507), .S0(n45[3]), .S1(n45[4]));   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_1006_add_4_5.INIT0 = 16'hfaaa;
    defparam counter_1006_add_4_5.INIT1 = 16'hfaaa;
    defparam counter_1006_add_4_5.INJECT1_0 = "NO";
    defparam counter_1006_add_4_5.INJECT1_1 = "NO";
    CCU2D counter_1006_add_4_3 (.A0(counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11505), .COUT(n11506), .S0(n45[1]), .S1(n45[2]));   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_1006_add_4_3.INIT0 = 16'hfaaa;
    defparam counter_1006_add_4_3.INIT1 = 16'hfaaa;
    defparam counter_1006_add_4_3.INJECT1_0 = "NO";
    defparam counter_1006_add_4_3.INJECT1_1 = "NO";
    CCU2D counter_1006_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n11505), .S1(n45[0]));   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_1006_add_4_1.INIT0 = 16'hF000;
    defparam counter_1006_add_4_1.INIT1 = 16'h0555;
    defparam counter_1006_add_4_1.INJECT1_0 = "NO";
    defparam counter_1006_add_4_1.INJECT1_1 = "NO";
    LUT4 i1154_1_lut (.A(\DemodOut[9] ), .Z(n3949[9])) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(26[3] 27[35])
    defparam i1154_1_lut.init = 16'h5555;
    FD1S3AX counter_1006__i1 (.D(n45[1]), .CK(osc_clk), .Q(counter[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_1006__i1.GSR = "ENABLED";
    FD1S3AX counter_1006__i2 (.D(n45[2]), .CK(osc_clk), .Q(counter[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_1006__i2.GSR = "ENABLED";
    FD1S3AX counter_1006__i3 (.D(n45[3]), .CK(osc_clk), .Q(counter[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_1006__i3.GSR = "ENABLED";
    FD1S3AX counter_1006__i4 (.D(n45[4]), .CK(osc_clk), .Q(counter[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_1006__i4.GSR = "ENABLED";
    FD1S3AX counter_1006__i5 (.D(n45[5]), .CK(osc_clk), .Q(counter[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_1006__i5.GSR = "ENABLED";
    FD1S3AX counter_1006__i6 (.D(n45[6]), .CK(osc_clk), .Q(counter[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_1006__i6.GSR = "ENABLED";
    FD1S3AX counter_1006__i7 (.D(n45[7]), .CK(osc_clk), .Q(counter[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_1006__i7.GSR = "ENABLED";
    FD1S3AX counter_1006__i8 (.D(n45[8]), .CK(osc_clk), .Q(counter[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_1006__i8.GSR = "ENABLED";
    FD1S3AX counter_1006__i9 (.D(n45[9]), .CK(osc_clk), .Q(counter[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_1006__i9.GSR = "ENABLED";
    FD1P3AX DataInReg__i2 (.D(\DataInReg_11__N_1856[1] ), .SP(osc_clk_enable_1406), 
            .CK(osc_clk), .Q(DataInReg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=189, LSE_RLINE=195 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i2.GSR = "ENABLED";
    FD1P3AX DataInReg__i3 (.D(\DataInReg_11__N_1856[2] ), .SP(osc_clk_enable_1406), 
            .CK(osc_clk), .Q(DataInReg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=189, LSE_RLINE=195 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i3.GSR = "ENABLED";
    FD1P3AX DataInReg__i4 (.D(\DataInReg_11__N_1856[3] ), .SP(osc_clk_enable_1406), 
            .CK(osc_clk), .Q(DataInReg[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=189, LSE_RLINE=195 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i4.GSR = "ENABLED";
    FD1P3AX DataInReg__i5 (.D(\DataInReg_11__N_1856[4] ), .SP(osc_clk_enable_1406), 
            .CK(osc_clk), .Q(DataInReg[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=189, LSE_RLINE=195 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i5.GSR = "ENABLED";
    FD1P3AX DataInReg__i6 (.D(\DataInReg_11__N_1856[5] ), .SP(osc_clk_enable_1406), 
            .CK(osc_clk), .Q(DataInReg[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=189, LSE_RLINE=195 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i6.GSR = "ENABLED";
    FD1P3AX DataInReg__i7 (.D(\DataInReg_11__N_1856[6] ), .SP(osc_clk_enable_1406), 
            .CK(osc_clk), .Q(DataInReg[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=189, LSE_RLINE=195 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i7.GSR = "ENABLED";
    FD1P3AX DataInReg__i8 (.D(\DataInReg_11__N_1856[7] ), .SP(osc_clk_enable_1406), 
            .CK(osc_clk), .Q(DataInReg[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=189, LSE_RLINE=195 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i8.GSR = "ENABLED";
    FD1P3AX DataInReg__i9 (.D(\DataInReg_11__N_1856[8] ), .SP(osc_clk_enable_1406), 
            .CK(osc_clk), .Q(DataInReg[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=189, LSE_RLINE=195 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i9.GSR = "ENABLED";
    FD1P3AX DataInReg__i10 (.D(n3949[9]), .SP(osc_clk_enable_1406), .CK(osc_clk), 
            .Q(DataInReg[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=189, LSE_RLINE=195 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i10.GSR = "ENABLED";
    CCU2D sub_765_add_2_11 (.A0(DataInReg[9]), .B0(counter[9]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n10974), .S1(PWMOut_N_1869));
    defparam sub_765_add_2_11.INIT0 = 16'h5999;
    defparam sub_765_add_2_11.INIT1 = 16'h0000;
    defparam sub_765_add_2_11.INJECT1_0 = "NO";
    defparam sub_765_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_765_add_2_9 (.A0(DataInReg[7]), .B0(counter[7]), .C0(GND_net), 
          .D0(GND_net), .A1(DataInReg[8]), .B1(counter[8]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10973), .COUT(n10974));
    defparam sub_765_add_2_9.INIT0 = 16'h5999;
    defparam sub_765_add_2_9.INIT1 = 16'h5999;
    defparam sub_765_add_2_9.INJECT1_0 = "NO";
    defparam sub_765_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_765_add_2_7 (.A0(DataInReg[5]), .B0(counter[5]), .C0(GND_net), 
          .D0(GND_net), .A1(DataInReg[6]), .B1(counter[6]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10972), .COUT(n10973));
    defparam sub_765_add_2_7.INIT0 = 16'h5999;
    defparam sub_765_add_2_7.INIT1 = 16'h5999;
    defparam sub_765_add_2_7.INJECT1_0 = "NO";
    defparam sub_765_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_765_add_2_5 (.A0(DataInReg[3]), .B0(counter[3]), .C0(GND_net), 
          .D0(GND_net), .A1(DataInReg[4]), .B1(counter[4]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10971), .COUT(n10972));
    defparam sub_765_add_2_5.INIT0 = 16'h5999;
    defparam sub_765_add_2_5.INIT1 = 16'h5999;
    defparam sub_765_add_2_5.INJECT1_0 = "NO";
    defparam sub_765_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_765_add_2_3 (.A0(DataInReg[1]), .B0(counter[1]), .C0(GND_net), 
          .D0(GND_net), .A1(DataInReg[2]), .B1(counter[2]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10970), .COUT(n10971));
    defparam sub_765_add_2_3.INIT0 = 16'h5999;
    defparam sub_765_add_2_3.INIT1 = 16'h5999;
    defparam sub_765_add_2_3.INJECT1_0 = "NO";
    defparam sub_765_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_765_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(DataInReg[0]), .B1(counter[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n10970));
    defparam sub_765_add_2_1.INIT0 = 16'h0000;
    defparam sub_765_add_2_1.INIT1 = 16'h5999;
    defparam sub_765_add_2_1.INJECT1_0 = "NO";
    defparam sub_765_add_2_1.INJECT1_1 = "NO";
    LUT4 i5_2_lut (.A(counter[2]), .B(counter[9]), .Z(n15)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(26[7:19])
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i1_2_lut (.A(counter[0]), .B(counter[5]), .Z(n11)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(26[7:19])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i2_2_lut (.A(counter[7]), .B(counter[3]), .Z(n12)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(26[7:19])
    defparam i2_2_lut.init = 16'heeee;
    
endmodule
//
// Verilog Description of module \uart_rx(CLKS_PER_BIT=87) 
//

module \uart_rx(CLKS_PER_BIT=87)  (osc_clk, i_Rx_Serial_c, o_Rx_Byte1, 
            GND_net, o_Rx_DV1) /* synthesis syn_module_defined=1 */ ;
    input osc_clk;
    input i_Rx_Serial_c;
    output [7:0]o_Rx_Byte1;
    input GND_net;
    output o_Rx_DV1;
    
    wire [7:0]UartClk /* synthesis SET_AS_NETWORK=\uart_rx1/UartClk[2], is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(37[14:21])
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(69[8:15])
    wire [2:0]r_Bit_Index;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(40[17:28])
    
    wire n13055, UartClk_2_enable_1;
    wire [15:0]r_Clock_Count;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(39[18:31])
    
    wire n8811;
    wire [2:0]r_SM_Main;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(43[17:26])
    
    wire n12984, r_Rx_DV_last, r_Rx_DV, n12746, n12748, n12740, 
        n12744, n12501, r_Rx_Data_R, r_Rx_Data;
    wire [7:0]r_Rx_Byte;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(41[17:26])
    
    wire UartClk_2_enable_16, UartClk_2_enable_32, n12642, n12770, n8827, 
        n13058, n13064, UartClk_2_enable_33;
    wire [2:0]n30;
    wire [2:0]n17;
    
    wire UartClk_2_enable_34, n12539, UartClk_2_enable_4, n12226;
    wire [2:0]r_SM_Main_2__N_2424;
    
    wire n12762, UartClk_2_enable_35, n11510, n12983, n12982, UartClk_2_enable_36, 
        n13065, UartClk_2_enable_5, UartClk_2_enable_6, r_Rx_DV_N_2484, 
        UartClk_2_enable_7, n12528, n13062, n8421, r_Rx_DV_last_N_2483, 
        n12973, n12719, n12530, n12651, n13073, UartClk_2_enable_30, 
        n8438;
    wire [15:0]n69;
    
    wire n8789, n12113, n12112, n12111, n12110, n12109, n12108, 
        n12107, n12106, n12758, n12593, n12776, n13071, n13072;
    
    LUT4 i5353_2_lut_3_lut_4_lut (.A(r_Bit_Index[1]), .B(n13055), .C(r_Bit_Index[2]), 
         .D(r_Bit_Index[0]), .Z(UartClk_2_enable_1)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(114[17:39])
    defparam i5353_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i2760_3_lut (.A(r_Clock_Count[1]), .B(r_Clock_Count[3]), .C(r_Clock_Count[2]), 
         .Z(n8811)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i2760_3_lut.init = 16'hecec;
    FD1S3IX r_SM_Main_i0 (.D(n12984), .CK(UartClk[2]), .CD(r_SM_Main[2]), 
            .Q(r_SM_Main[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam r_SM_Main_i0.GSR = "ENABLED";
    FD1S3AX r_Rx_DV_last_60 (.D(r_Rx_DV), .CK(osc_clk), .Q(r_Rx_DV_last)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(47[11] 52[8])
    defparam r_Rx_DV_last_60.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(n12746), .B(n12748), .C(n12740), .D(n12744), .Z(n12501)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(85[17:52])
    defparam i1_4_lut.init = 16'hfffe;
    FD1S3AY r_Rx_Data_R_61 (.D(i_Rx_Serial_c), .CK(UartClk[2]), .Q(r_Rx_Data_R)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(57[11] 62[8])
    defparam r_Rx_Data_R_61.GSR = "ENABLED";
    FD1S3AY r_Rx_Data_62 (.D(r_Rx_Data_R), .CK(UartClk[2]), .Q(r_Rx_Data)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(57[11] 62[8])
    defparam r_Rx_Data_62.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(r_Clock_Count[11]), .B(r_Clock_Count[15]), .Z(n12746)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(85[17:52])
    defparam i1_2_lut.init = 16'heeee;
    FD1P3AX r_Rx_Byte_i4 (.D(r_Rx_Data), .SP(UartClk_2_enable_1), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam r_Rx_Byte_i4.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i0 (.D(r_Rx_Byte[0]), .SP(UartClk_2_enable_16), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam o_Rx_Byte_i0.GSR = "ENABLED";
    FD1P3AX r_Bit_Index_i0 (.D(n12642), .SP(UartClk_2_enable_32), .CK(UartClk[2]), 
            .Q(r_Bit_Index[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam r_Bit_Index_i0.GSR = "ENABLED";
    LUT4 i1_3_lut (.A(r_Clock_Count[13]), .B(r_Clock_Count[8]), .C(r_Clock_Count[7]), 
         .Z(n12748)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(85[17:52])
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_adj_49 (.A(r_Clock_Count[14]), .B(r_Clock_Count[10]), 
         .Z(n12740)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(85[17:52])
    defparam i1_2_lut_adj_49.init = 16'heeee;
    LUT4 i1_2_lut_adj_50 (.A(r_Clock_Count[9]), .B(r_Clock_Count[12]), .Z(n12744)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(85[17:52])
    defparam i1_2_lut_adj_50.init = 16'heeee;
    LUT4 i5338_4_lut (.A(n12770), .B(n12501), .C(n8827), .D(r_SM_Main[1]), 
         .Z(UartClk_2_enable_32)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;
    defparam i5338_4_lut.init = 16'h5455;
    LUT4 i5359_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n13058), .C(n13064), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_33)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(114[17:39])
    defparam i5359_2_lut_3_lut_4_lut.init = 16'h1000;
    FD1S3AX UartClk_1007_1029__i0 (.D(n17[0]), .CK(osc_clk), .Q(n30[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(49[15:29])
    defparam UartClk_1007_1029__i0.GSR = "ENABLED";
    LUT4 i5357_2_lut_3_lut_4_lut (.A(r_Bit_Index[1]), .B(n13055), .C(r_Bit_Index[2]), 
         .D(r_Bit_Index[0]), .Z(UartClk_2_enable_34)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(114[17:39])
    defparam i5357_2_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 i5351_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n13058), .C(n12539), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_4)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(114[17:39])
    defparam i5351_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_adj_51 (.A(r_SM_Main[0]), .B(r_SM_Main[2]), .Z(n12770)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_51.init = 16'heeee;
    LUT4 i1_4_lut_adj_52 (.A(r_Clock_Count[3]), .B(n12226), .C(r_Clock_Count[5]), 
         .D(r_Clock_Count[0]), .Z(r_SM_Main_2__N_2424[0])) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;
    defparam i1_4_lut_adj_52.init = 16'hdfff;
    LUT4 i1_4_lut_adj_53 (.A(r_Clock_Count[1]), .B(n12501), .C(n12762), 
         .D(r_Clock_Count[6]), .Z(n12226)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(85[17:52])
    defparam i1_4_lut_adj_53.init = 16'hfffd;
    LUT4 i5355_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n13058), .C(n13064), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_35)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(114[17:39])
    defparam i5355_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_adj_54 (.A(r_Clock_Count[2]), .B(r_Clock_Count[4]), .Z(n12762)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(85[17:52])
    defparam i1_2_lut_adj_54.init = 16'heeee;
    CCU2D UartClk_1007_1029_add_4_3 (.A0(n30[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(UartClk[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11510), .S0(n17[1]), .S1(n17[2]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(49[15:29])
    defparam UartClk_1007_1029_add_4_3.INIT0 = 16'hfaaa;
    defparam UartClk_1007_1029_add_4_3.INIT1 = 16'hfaaa;
    defparam UartClk_1007_1029_add_4_3.INJECT1_0 = "NO";
    defparam UartClk_1007_1029_add_4_3.INJECT1_1 = "NO";
    CCU2D UartClk_1007_1029_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n30[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n11510), .S1(n17[0]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(49[15:29])
    defparam UartClk_1007_1029_add_4_1.INIT0 = 16'hF000;
    defparam UartClk_1007_1029_add_4_1.INIT1 = 16'h0555;
    defparam UartClk_1007_1029_add_4_1.INJECT1_0 = "NO";
    defparam UartClk_1007_1029_add_4_1.INJECT1_1 = "NO";
    FD1P3AX r_Rx_Byte_i3 (.D(r_Rx_Data), .SP(UartClk_2_enable_4), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam r_Rx_Byte_i3.GSR = "ENABLED";
    PFUMX i5403 (.BLUT(n12983), .ALUT(n12982), .C0(r_SM_Main[1]), .Z(n12984));
    LUT4 i5327_2_lut_3_lut_4_lut (.A(r_Bit_Index[1]), .B(n13055), .C(r_Bit_Index[2]), 
         .D(r_Bit_Index[0]), .Z(UartClk_2_enable_36)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(114[17:39])
    defparam i5327_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i5378_2_lut_3_lut_4_lut (.A(n8827), .B(n12501), .C(r_SM_Main[0]), 
         .D(n13065), .Z(UartClk_2_enable_16)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i5378_2_lut_3_lut_4_lut.init = 16'h00e0;
    FD1P3AX r_Rx_Byte_i2 (.D(r_Rx_Data), .SP(UartClk_2_enable_5), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam r_Rx_Byte_i2.GSR = "ENABLED";
    FD1P3AX r_Rx_DV_64 (.D(r_Rx_DV_N_2484), .SP(UartClk_2_enable_6), .CK(UartClk[2]), 
            .Q(r_Rx_DV)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam r_Rx_DV_64.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i1 (.D(r_Rx_Data), .SP(UartClk_2_enable_7), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam r_Rx_Byte_i1.GSR = "ENABLED";
    FD1S3IX r_SM_Main_i2 (.D(n13062), .CK(UartClk[2]), .CD(n12528), .Q(r_SM_Main[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam r_SM_Main_i2.GSR = "ENABLED";
    LUT4 i2368_1_lut (.A(r_Rx_DV), .Z(n8421)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam i2368_1_lut.init = 16'h5555;
    LUT4 r_Rx_DV_last_I_0_1_lut (.A(r_Rx_DV_last), .Z(r_Rx_DV_last_N_2483)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(50[30:43])
    defparam r_Rx_DV_last_I_0_1_lut.init = 16'h5555;
    LUT4 i1_2_lut_adj_55 (.A(r_Bit_Index[2]), .B(r_Bit_Index[0]), .Z(n12539)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(114[17:39])
    defparam i1_2_lut_adj_55.init = 16'hbbbb;
    LUT4 i4_4_lut (.A(n12973), .B(r_SM_Main[0]), .C(r_SM_Main[1]), .D(n13062), 
         .Z(n12719)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i4_4_lut.init = 16'h2000;
    LUT4 i2_4_lut (.A(r_Bit_Index[0]), .B(n13062), .C(r_Bit_Index[1]), 
         .D(n12530), .Z(n12651)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C (D))))) */ ;
    defparam i2_4_lut.init = 16'h4800;
    LUT4 i5348_2_lut_3_lut_4_lut (.A(r_Bit_Index[1]), .B(n13055), .C(r_Bit_Index[2]), 
         .D(r_Bit_Index[0]), .Z(UartClk_2_enable_5)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(114[17:39])
    defparam i5348_2_lut_3_lut_4_lut.init = 16'h0002;
    FD1S3IX r_SM_Main_i1 (.D(n13073), .CK(UartClk[2]), .CD(r_SM_Main[2]), 
            .Q(r_SM_Main[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam r_SM_Main_i1.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i1 (.D(r_Rx_Byte[1]), .SP(UartClk_2_enable_16), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam o_Rx_Byte_i1.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i0 (.D(n69[0]), .SP(UartClk_2_enable_30), 
            .CD(n8438), .CK(UartClk[2]), .Q(r_Clock_Count[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009__i0.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i15 (.D(n69[15]), .SP(UartClk_2_enable_30), 
            .CD(n8438), .CK(UartClk[2]), .Q(r_Clock_Count[15])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009__i15.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i2 (.D(r_Rx_Byte[2]), .SP(UartClk_2_enable_16), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam o_Rx_Byte_i2.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i3 (.D(r_Rx_Byte[3]), .SP(UartClk_2_enable_16), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam o_Rx_Byte_i3.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i4 (.D(r_Rx_Byte[4]), .SP(UartClk_2_enable_16), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam o_Rx_Byte_i4.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i5 (.D(r_Rx_Byte[5]), .SP(UartClk_2_enable_16), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam o_Rx_Byte_i5.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i6 (.D(r_Rx_Byte[6]), .SP(UartClk_2_enable_16), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam o_Rx_Byte_i6.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i7 (.D(r_Rx_Byte[7]), .SP(UartClk_2_enable_16), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam o_Rx_Byte_i7.GSR = "ENABLED";
    FD1S3AX UartClk_1007_1029__i1 (.D(n17[1]), .CK(osc_clk), .Q(n30[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(49[15:29])
    defparam UartClk_1007_1029__i1.GSR = "ENABLED";
    FD1S3AX UartClk_1007_1029__i2 (.D(n17[2]), .CK(osc_clk), .Q(UartClk[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(49[15:29])
    defparam UartClk_1007_1029__i2.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i14 (.D(n69[14]), .SP(UartClk_2_enable_30), 
            .CD(n8438), .CK(UartClk[2]), .Q(r_Clock_Count[14])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009__i14.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_88 (.A(n8827), .B(n12501), .Z(n13062)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_88.init = 16'heeee;
    LUT4 i5369_2_lut_3_lut_4_lut (.A(n8827), .B(n12501), .C(n13065), .D(r_SM_Main[0]), 
         .Z(r_Rx_DV_N_2484)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;
    defparam i5369_2_lut_3_lut_4_lut.init = 16'h0e00;
    LUT4 r_SM_Main_2__N_2418_2__bdd_3_lut_5402_4_lut (.A(n8827), .B(n12501), 
         .C(r_SM_Main[0]), .D(n8789), .Z(n12982)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C)))) */ ;
    defparam r_SM_Main_2__N_2418_2__bdd_3_lut_5402_4_lut.init = 16'h1e10;
    LUT4 i2_3_lut_4_lut (.A(n8827), .B(n12501), .C(r_Bit_Index[0]), .D(n12530), 
         .Z(n12642)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0e00;
    LUT4 i2776_4_lut (.A(n8811), .B(r_Clock_Count[6]), .C(r_Clock_Count[5]), 
         .D(r_Clock_Count[4]), .Z(n8827)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i2776_4_lut.init = 16'hc8c0;
    CCU2D r_Clock_Count_1009_add_4_17 (.A0(r_Clock_Count[15]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12113), .S0(n69[15]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_17.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_1009_add_4_17.INIT1 = 16'h0000;
    defparam r_Clock_Count_1009_add_4_17.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_17.INJECT1_1 = "NO";
    FD1P3IX r_Clock_Count_1009__i13 (.D(n69[13]), .SP(UartClk_2_enable_30), 
            .CD(n8438), .CK(UartClk[2]), .Q(r_Clock_Count[13])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009__i13.GSR = "ENABLED";
    CCU2D r_Clock_Count_1009_add_4_15 (.A0(r_Clock_Count[13]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[14]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12112), .COUT(n12113), .S0(n69[13]), 
          .S1(n69[14]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_15.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_1009_add_4_15.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_1009_add_4_15.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_15.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_1009_add_4_13 (.A0(r_Clock_Count[11]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[12]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12111), .COUT(n12112), .S0(n69[11]), 
          .S1(n69[12]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_13.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_1009_add_4_13.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_1009_add_4_13.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_13.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_1009_add_4_11 (.A0(r_Clock_Count[9]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[10]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12110), .COUT(n12111), .S0(n69[9]), 
          .S1(n69[10]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_11.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_1009_add_4_11.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_1009_add_4_11.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_11.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_1009_add_4_9 (.A0(r_Clock_Count[7]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[8]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12109), .COUT(n12110), .S0(n69[7]), 
          .S1(n69[8]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_9.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_1009_add_4_9.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_1009_add_4_9.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_9.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_1009_add_4_7 (.A0(r_Clock_Count[5]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[6]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12108), .COUT(n12109), .S0(n69[5]), 
          .S1(n69[6]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_7.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_1009_add_4_7.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_1009_add_4_7.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_7.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_1009_add_4_5 (.A0(r_Clock_Count[3]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[4]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12107), .COUT(n12108), .S0(n69[3]), 
          .S1(n69[4]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_5.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_1009_add_4_5.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_1009_add_4_5.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_5.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_1009_add_4_3 (.A0(r_Clock_Count[1]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[2]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12106), .COUT(n12107), .S0(n69[1]), 
          .S1(n69[2]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_3.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_1009_add_4_3.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_1009_add_4_3.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_3.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_1009_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(r_Clock_Count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n12106), .S1(n69[0]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009_add_4_1.INIT0 = 16'hF000;
    defparam r_Clock_Count_1009_add_4_1.INIT1 = 16'h0555;
    defparam r_Clock_Count_1009_add_4_1.INJECT1_0 = "NO";
    defparam r_Clock_Count_1009_add_4_1.INJECT1_1 = "NO";
    LUT4 i5376_4_lut (.A(r_SM_Main[2]), .B(r_SM_Main[1]), .C(r_SM_Main_2__N_2424[0]), 
         .D(n12758), .Z(UartClk_2_enable_30)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(69[7] 161[14])
    defparam i5376_4_lut.init = 16'h5455;
    LUT4 i1_2_lut_adj_56 (.A(r_Rx_Data), .B(r_SM_Main[0]), .Z(n12758)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_56.init = 16'h8888;
    LUT4 i1_4_lut_adj_57 (.A(r_SM_Main[2]), .B(n12593), .C(n13062), .D(r_SM_Main[1]), 
         .Z(n8438)) /* synthesis lut_function=(!(A+!(B (C (D))+!B (C+!(D))))) */ ;
    defparam i1_4_lut_adj_57.init = 16'h5011;
    LUT4 i5109_3_lut (.A(n12776), .B(r_SM_Main[0]), .C(n12226), .Z(n12593)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i5109_3_lut.init = 16'hc8c8;
    LUT4 i1_4_lut_adj_58 (.A(r_Clock_Count[5]), .B(r_Clock_Count[0]), .C(r_Clock_Count[3]), 
         .D(r_Rx_Data), .Z(n12776)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_4_lut_adj_58.init = 16'hff7f;
    LUT4 r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_else_3_lut (.A(r_SM_Main_2__N_2424[0]), 
         .B(r_Rx_Data), .C(r_SM_Main[0]), .Z(n13071)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(69[7] 161[14])
    defparam r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_else_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_adj_59 (.A(r_SM_Main[1]), .B(r_SM_Main[0]), .Z(n12530)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_59.init = 16'h2222;
    LUT4 i5345_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n13058), .C(n12539), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_7)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(114[17:39])
    defparam i5345_2_lut_3_lut_4_lut.init = 16'h0001;
    FD1P3IX r_Clock_Count_1009__i12 (.D(n69[12]), .SP(UartClk_2_enable_30), 
            .CD(n8438), .CK(UartClk[2]), .Q(r_Clock_Count[12])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009__i12.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i11 (.D(n69[11]), .SP(UartClk_2_enable_30), 
            .CD(n8438), .CK(UartClk[2]), .Q(r_Clock_Count[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009__i11.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i10 (.D(n69[10]), .SP(UartClk_2_enable_30), 
            .CD(n8438), .CK(UartClk[2]), .Q(r_Clock_Count[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009__i10.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i9 (.D(n69[9]), .SP(UartClk_2_enable_30), 
            .CD(n8438), .CK(UartClk[2]), .Q(r_Clock_Count[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009__i9.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i8 (.D(n69[8]), .SP(UartClk_2_enable_30), 
            .CD(n8438), .CK(UartClk[2]), .Q(r_Clock_Count[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009__i8.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i7 (.D(n69[7]), .SP(UartClk_2_enable_30), 
            .CD(n8438), .CK(UartClk[2]), .Q(r_Clock_Count[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009__i7.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i6 (.D(n69[6]), .SP(UartClk_2_enable_30), 
            .CD(n8438), .CK(UartClk[2]), .Q(r_Clock_Count[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009__i6.GSR = "ENABLED";
    LUT4 i21_4_lut_4_lut (.A(r_SM_Main[1]), .B(r_SM_Main[2]), .C(r_SM_Main[0]), 
         .D(n13062), .Z(UartClk_2_enable_6)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(69[7] 161[14])
    defparam i21_4_lut_4_lut.init = 16'h2505;
    LUT4 i5341_2_lut_3_lut (.A(r_SM_Main[1]), .B(r_SM_Main[2]), .C(r_SM_Main[0]), 
         .Z(n12528)) /* synthesis lut_function=((B+!(C))+!A) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(69[7] 161[14])
    defparam i5341_2_lut_3_lut.init = 16'hdfdf;
    FD1S3IX o_Rx_DV_59 (.D(r_Rx_DV_last_N_2483), .CK(osc_clk), .CD(n8421), 
            .Q(o_Rx_DV1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(47[11] 52[8])
    defparam o_Rx_DV_59.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_90 (.A(r_Bit_Index[2]), .B(r_Bit_Index[0]), .Z(n13064)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_90.init = 16'h8888;
    LUT4 r_Bit_Index_2__bdd_3_lut (.A(r_Bit_Index[2]), .B(r_Bit_Index[1]), 
         .C(r_Bit_Index[0]), .Z(n12973)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;
    defparam r_Bit_Index_2__bdd_3_lut.init = 16'h6a6a;
    LUT4 i2_2_lut_3_lut (.A(r_Bit_Index[2]), .B(r_Bit_Index[0]), .C(r_Bit_Index[1]), 
         .Z(n8789)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut.init = 16'h8080;
    FD1P3IX r_Clock_Count_1009__i5 (.D(n69[5]), .SP(UartClk_2_enable_30), 
            .CD(n8438), .CK(UartClk[2]), .Q(r_Clock_Count[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009__i5.GSR = "ENABLED";
    LUT4 r_SM_Main_2__N_2418_2__bdd_3_lut (.A(r_SM_Main_2__N_2424[0]), .B(r_Rx_Data), 
         .C(r_SM_Main[0]), .Z(n12983)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+(C))) */ ;
    defparam r_SM_Main_2__N_2418_2__bdd_3_lut.init = 16'ha3a3;
    FD1P3IX r_Clock_Count_1009__i4 (.D(n69[4]), .SP(UartClk_2_enable_30), 
            .CD(n8438), .CK(UartClk[2]), .Q(r_Clock_Count[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009__i4.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i3 (.D(n69[3]), .SP(UartClk_2_enable_30), 
            .CD(n8438), .CK(UartClk[2]), .Q(r_Clock_Count[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009__i3.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i2 (.D(n69[2]), .SP(UartClk_2_enable_30), 
            .CD(n8438), .CK(UartClk[2]), .Q(r_Clock_Count[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009__i2.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1009__i1 (.D(n69[1]), .SP(UartClk_2_enable_30), 
            .CD(n8438), .CK(UartClk[2]), .Q(r_Clock_Count[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(137[34:54])
    defparam r_Clock_Count_1009__i1.GSR = "ENABLED";
    LUT4 r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_then_3_lut (.A(n12501), .B(n8827), 
         .C(r_SM_Main[0]), .Z(n13072)) /* synthesis lut_function=(!(A (C)+!A (B (C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(69[7] 161[14])
    defparam r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_then_3_lut.init = 16'h1f1f;
    FD1P3AX r_Bit_Index_i2 (.D(n12719), .SP(UartClk_2_enable_32), .CK(UartClk[2]), 
            .Q(r_Bit_Index[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam r_Bit_Index_i2.GSR = "ENABLED";
    FD1P3AX r_Bit_Index_i1 (.D(n12651), .SP(UartClk_2_enable_32), .CK(UartClk[2]), 
            .Q(r_Bit_Index[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam r_Bit_Index_i1.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_91 (.A(r_SM_Main[2]), .B(r_SM_Main[1]), .Z(n13065)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_91.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_84_3_lut_4_lut (.A(r_SM_Main[2]), .B(r_SM_Main[1]), 
         .C(n12501), .D(n8827), .Z(n13058)) /* synthesis lut_function=(A+!(B (C+(D)))) */ ;
    defparam i1_2_lut_rep_84_3_lut_4_lut.init = 16'hbbbf;
    FD1P3AX r_Rx_Byte_i7 (.D(r_Rx_Data), .SP(UartClk_2_enable_33), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam r_Rx_Byte_i7.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i6 (.D(r_Rx_Data), .SP(UartClk_2_enable_34), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam r_Rx_Byte_i6.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i5 (.D(r_Rx_Data), .SP(UartClk_2_enable_35), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam r_Rx_Byte_i5.GSR = "ENABLED";
    PFUMX i5432 (.BLUT(n13071), .ALUT(n13072), .C0(r_SM_Main[1]), .Z(n13073));
    FD1P3AX r_Rx_Byte_i0 (.D(r_Rx_Data), .SP(UartClk_2_enable_36), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=220, LSE_RLINE=225 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(66[10] 162[8])
    defparam r_Rx_Byte_i0.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_81_3_lut_4_lut (.A(n8827), .B(n12501), .C(r_SM_Main[0]), 
         .D(n13065), .Z(n13055)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;
    defparam i1_2_lut_rep_81_3_lut_4_lut.init = 16'hfff1;
    
endmodule
//
// Verilog Description of module Mixer
//

module Mixer (MixerOutSin, osc_clk, DiffOut_c, MixerOutCos, RFIn_c, 
            \LOCosine[12] , GND_net, \LOCosine[10] , \LOCosine[11] , 
            \LOCosine[8] , \LOCosine[9] , \LOCosine[6] , \LOCosine[7] , 
            \LOCosine[4] , \LOCosine[5] , \LOCosine[2] , \LOCosine[3] , 
            \LOCosine[1] , \LOSine[12] , \LOSine[10] , \LOSine[11] , 
            \LOSine[8] , \LOSine[9] , \LOSine[6] , \LOSine[7] , \LOSine[4] , 
            \LOSine[5] , \LOSine[2] , \LOSine[3] , \LOSine[1] ) /* synthesis syn_module_defined=1 */ ;
    output [11:0]MixerOutSin;
    input osc_clk;
    output DiffOut_c;
    output [11:0]MixerOutCos;
    input RFIn_c;
    input \LOCosine[12] ;
    input GND_net;
    input \LOCosine[10] ;
    input \LOCosine[11] ;
    input \LOCosine[8] ;
    input \LOCosine[9] ;
    input \LOCosine[6] ;
    input \LOCosine[7] ;
    input \LOCosine[4] ;
    input \LOCosine[5] ;
    input \LOCosine[2] ;
    input \LOCosine[3] ;
    input \LOCosine[1] ;
    input \LOSine[12] ;
    input \LOSine[10] ;
    input \LOSine[11] ;
    input \LOSine[8] ;
    input \LOSine[9] ;
    input \LOSine[6] ;
    input \LOSine[7] ;
    input \LOSine[4] ;
    input \LOSine[5] ;
    input \LOSine[2] ;
    input \LOSine[3] ;
    input \LOSine[1] ;
    
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(69[8:15])
    wire [11:0]MixerOutSin_11__N_212;
    
    wire RFInR;
    wire [11:0]MixerOutCos_11__N_224;
    
    wire n11054;
    wire [11:0]MixerOutCos_11__N_250;
    
    wire n11053, n11052, n11051, n11050, n11049, n11016;
    wire [11:0]MixerOutSin_11__N_236;
    
    wire n11015, n11014, n11013, n11012, n11011;
    
    FD1S3AX MixerOutSin_i0 (.D(MixerOutSin_11__N_212[0]), .CK(osc_clk), 
            .Q(MixerOutSin[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i0.GSR = "ENABLED";
    FD1S3AY RFInR_14 (.D(DiffOut_c), .CK(osc_clk), .Q(RFInR)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(23[10] 27[8])
    defparam RFInR_14.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i0 (.D(MixerOutCos_11__N_224[0]), .CK(osc_clk), 
            .Q(MixerOutCos[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i0.GSR = "ENABLED";
    FD1S3AY RFInR1_13 (.D(RFIn_c), .CK(osc_clk), .Q(DiffOut_c)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(23[10] 27[8])
    defparam RFInR1_13.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i1 (.D(MixerOutSin_11__N_212[1]), .CK(osc_clk), 
            .Q(MixerOutSin[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i1.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i2 (.D(MixerOutSin_11__N_212[2]), .CK(osc_clk), 
            .Q(MixerOutSin[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i2.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i3 (.D(MixerOutSin_11__N_212[3]), .CK(osc_clk), 
            .Q(MixerOutSin[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i3.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i4 (.D(MixerOutSin_11__N_212[4]), .CK(osc_clk), 
            .Q(MixerOutSin[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i4.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i5 (.D(MixerOutSin_11__N_212[5]), .CK(osc_clk), 
            .Q(MixerOutSin[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i5.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i6 (.D(MixerOutSin_11__N_212[6]), .CK(osc_clk), 
            .Q(MixerOutSin[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i6.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i7 (.D(MixerOutSin_11__N_212[7]), .CK(osc_clk), 
            .Q(MixerOutSin[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i7.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i8 (.D(MixerOutSin_11__N_212[8]), .CK(osc_clk), 
            .Q(MixerOutSin[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i8.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i9 (.D(MixerOutSin_11__N_212[9]), .CK(osc_clk), 
            .Q(MixerOutSin[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i9.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i10 (.D(MixerOutSin_11__N_212[10]), .CK(osc_clk), 
            .Q(MixerOutSin[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i10.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i11 (.D(MixerOutSin_11__N_212[11]), .CK(osc_clk), 
            .Q(MixerOutSin[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i11.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i1 (.D(MixerOutCos_11__N_224[1]), .CK(osc_clk), 
            .Q(MixerOutCos[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i1.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i2 (.D(MixerOutCos_11__N_224[2]), .CK(osc_clk), 
            .Q(MixerOutCos[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i2.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i3 (.D(MixerOutCos_11__N_224[3]), .CK(osc_clk), 
            .Q(MixerOutCos[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i3.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i4 (.D(MixerOutCos_11__N_224[4]), .CK(osc_clk), 
            .Q(MixerOutCos[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i4.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i5 (.D(MixerOutCos_11__N_224[5]), .CK(osc_clk), 
            .Q(MixerOutCos[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i5.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i6 (.D(MixerOutCos_11__N_224[6]), .CK(osc_clk), 
            .Q(MixerOutCos[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i6.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i7 (.D(MixerOutCos_11__N_224[7]), .CK(osc_clk), 
            .Q(MixerOutCos[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i7.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i8 (.D(MixerOutCos_11__N_224[8]), .CK(osc_clk), 
            .Q(MixerOutCos[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i8.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i9 (.D(MixerOutCos_11__N_224[9]), .CK(osc_clk), 
            .Q(MixerOutCos[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i9.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i10 (.D(MixerOutCos_11__N_224[10]), .CK(osc_clk), 
            .Q(MixerOutCos[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i10.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i11 (.D(MixerOutCos_11__N_224[11]), .CK(osc_clk), 
            .Q(MixerOutCos[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=168 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i11.GSR = "ENABLED";
    CCU2D unary_minus_7_add_3_13 (.A0(\LOCosine[12] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11054), .S0(MixerOutCos_11__N_250[11]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(42[26:33])
    defparam unary_minus_7_add_3_13.INIT0 = 16'hf555;
    defparam unary_minus_7_add_3_13.INIT1 = 16'h0000;
    defparam unary_minus_7_add_3_13.INJECT1_0 = "NO";
    defparam unary_minus_7_add_3_13.INJECT1_1 = "NO";
    CCU2D unary_minus_7_add_3_11 (.A0(\LOCosine[10] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOCosine[11] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11053), .COUT(n11054), .S0(MixerOutCos_11__N_250[9]), 
          .S1(MixerOutCos_11__N_250[10]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(42[26:33])
    defparam unary_minus_7_add_3_11.INIT0 = 16'hf555;
    defparam unary_minus_7_add_3_11.INIT1 = 16'hf555;
    defparam unary_minus_7_add_3_11.INJECT1_0 = "NO";
    defparam unary_minus_7_add_3_11.INJECT1_1 = "NO";
    CCU2D unary_minus_7_add_3_9 (.A0(\LOCosine[8] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOCosine[9] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11052), .COUT(n11053), .S0(MixerOutCos_11__N_250[7]), 
          .S1(MixerOutCos_11__N_250[8]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(42[26:33])
    defparam unary_minus_7_add_3_9.INIT0 = 16'hf555;
    defparam unary_minus_7_add_3_9.INIT1 = 16'hf555;
    defparam unary_minus_7_add_3_9.INJECT1_0 = "NO";
    defparam unary_minus_7_add_3_9.INJECT1_1 = "NO";
    CCU2D unary_minus_7_add_3_7 (.A0(\LOCosine[6] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOCosine[7] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11051), .COUT(n11052), .S0(MixerOutCos_11__N_250[5]), 
          .S1(MixerOutCos_11__N_250[6]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(42[26:33])
    defparam unary_minus_7_add_3_7.INIT0 = 16'hf555;
    defparam unary_minus_7_add_3_7.INIT1 = 16'hf555;
    defparam unary_minus_7_add_3_7.INJECT1_0 = "NO";
    defparam unary_minus_7_add_3_7.INJECT1_1 = "NO";
    CCU2D unary_minus_7_add_3_5 (.A0(\LOCosine[4] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOCosine[5] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11050), .COUT(n11051), .S0(MixerOutCos_11__N_250[3]), 
          .S1(MixerOutCos_11__N_250[4]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(42[26:33])
    defparam unary_minus_7_add_3_5.INIT0 = 16'hf555;
    defparam unary_minus_7_add_3_5.INIT1 = 16'hf555;
    defparam unary_minus_7_add_3_5.INJECT1_0 = "NO";
    defparam unary_minus_7_add_3_5.INJECT1_1 = "NO";
    CCU2D unary_minus_7_add_3_3 (.A0(\LOCosine[2] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOCosine[3] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11049), .COUT(n11050), .S0(MixerOutCos_11__N_250[1]), 
          .S1(MixerOutCos_11__N_250[2]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(42[26:33])
    defparam unary_minus_7_add_3_3.INIT0 = 16'hf555;
    defparam unary_minus_7_add_3_3.INIT1 = 16'hf555;
    defparam unary_minus_7_add_3_3.INJECT1_0 = "NO";
    defparam unary_minus_7_add_3_3.INJECT1_1 = "NO";
    CCU2D unary_minus_7_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOCosine[1] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n11049), .S1(MixerOutCos_11__N_250[0]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(42[26:33])
    defparam unary_minus_7_add_3_1.INIT0 = 16'hF000;
    defparam unary_minus_7_add_3_1.INIT1 = 16'h0aaa;
    defparam unary_minus_7_add_3_1.INJECT1_0 = "NO";
    defparam unary_minus_7_add_3_1.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_13 (.A0(\LOSine[12] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11016), .S0(MixerOutSin_11__N_236[11]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(41[26:33])
    defparam unary_minus_6_add_3_13.INIT0 = 16'hf555;
    defparam unary_minus_6_add_3_13.INIT1 = 16'h0000;
    defparam unary_minus_6_add_3_13.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_13.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_11 (.A0(\LOSine[10] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOSine[11] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11015), .COUT(n11016), .S0(MixerOutSin_11__N_236[9]), 
          .S1(MixerOutSin_11__N_236[10]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(41[26:33])
    defparam unary_minus_6_add_3_11.INIT0 = 16'hf555;
    defparam unary_minus_6_add_3_11.INIT1 = 16'hf555;
    defparam unary_minus_6_add_3_11.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_11.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_9 (.A0(\LOSine[8] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOSine[9] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11014), .COUT(n11015), .S0(MixerOutSin_11__N_236[7]), 
          .S1(MixerOutSin_11__N_236[8]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(41[26:33])
    defparam unary_minus_6_add_3_9.INIT0 = 16'hf555;
    defparam unary_minus_6_add_3_9.INIT1 = 16'hf555;
    defparam unary_minus_6_add_3_9.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_9.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_7 (.A0(\LOSine[6] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOSine[7] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11013), .COUT(n11014), .S0(MixerOutSin_11__N_236[5]), 
          .S1(MixerOutSin_11__N_236[6]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(41[26:33])
    defparam unary_minus_6_add_3_7.INIT0 = 16'hf555;
    defparam unary_minus_6_add_3_7.INIT1 = 16'hf555;
    defparam unary_minus_6_add_3_7.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_7.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_5 (.A0(\LOSine[4] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOSine[5] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11012), .COUT(n11013), .S0(MixerOutSin_11__N_236[3]), 
          .S1(MixerOutSin_11__N_236[4]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(41[26:33])
    defparam unary_minus_6_add_3_5.INIT0 = 16'hf555;
    defparam unary_minus_6_add_3_5.INIT1 = 16'hf555;
    defparam unary_minus_6_add_3_5.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_5.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_3 (.A0(\LOSine[2] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOSine[3] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11011), .COUT(n11012), .S0(MixerOutSin_11__N_236[1]), 
          .S1(MixerOutSin_11__N_236[2]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(41[26:33])
    defparam unary_minus_6_add_3_3.INIT0 = 16'hf555;
    defparam unary_minus_6_add_3_3.INIT1 = 16'hf555;
    defparam unary_minus_6_add_3_3.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_3.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOSine[1] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n11011), .S1(MixerOutSin_11__N_236[0]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(41[26:33])
    defparam unary_minus_6_add_3_1.INIT0 = 16'hF000;
    defparam unary_minus_6_add_3_1.INIT1 = 16'h0aaa;
    defparam unary_minus_6_add_3_1.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_1.INJECT1_1 = "NO";
    LUT4 MixerOutCos_11__I_0_i2_3_lut (.A(\LOCosine[2] ), .B(MixerOutCos_11__N_250[1]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i3_3_lut (.A(\LOCosine[3] ), .B(MixerOutCos_11__N_250[2]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i4_3_lut (.A(\LOCosine[4] ), .B(MixerOutCos_11__N_250[3]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i5_3_lut (.A(\LOCosine[5] ), .B(MixerOutCos_11__N_250[4]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i6_3_lut (.A(\LOCosine[6] ), .B(MixerOutCos_11__N_250[5]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i7_3_lut (.A(\LOCosine[7] ), .B(MixerOutCos_11__N_250[6]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i8_3_lut (.A(\LOCosine[8] ), .B(MixerOutCos_11__N_250[7]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i9_3_lut (.A(\LOCosine[9] ), .B(MixerOutCos_11__N_250[8]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i2_3_lut (.A(\LOSine[2] ), .B(MixerOutSin_11__N_236[1]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i3_3_lut (.A(\LOSine[3] ), .B(MixerOutSin_11__N_236[2]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i10_3_lut (.A(\LOCosine[10] ), .B(MixerOutCos_11__N_250[9]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i4_3_lut (.A(\LOSine[4] ), .B(MixerOutSin_11__N_236[3]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i5_3_lut (.A(\LOSine[5] ), .B(MixerOutSin_11__N_236[4]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i6_3_lut (.A(\LOSine[6] ), .B(MixerOutSin_11__N_236[5]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i7_3_lut (.A(\LOSine[7] ), .B(MixerOutSin_11__N_236[6]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i8_3_lut (.A(\LOSine[8] ), .B(MixerOutSin_11__N_236[7]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i9_3_lut (.A(\LOSine[9] ), .B(MixerOutSin_11__N_236[8]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i10_3_lut (.A(\LOSine[10] ), .B(MixerOutSin_11__N_236[9]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i11_3_lut (.A(\LOSine[11] ), .B(MixerOutSin_11__N_236[10]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i11_3_lut (.A(\LOCosine[11] ), .B(MixerOutCos_11__N_250[10]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i12_3_lut (.A(\LOCosine[12] ), .B(MixerOutCos_11__N_250[11]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i12_3_lut (.A(\LOSine[12] ), .B(MixerOutSin_11__N_236[11]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i1_3_lut (.A(\LOSine[1] ), .B(MixerOutSin_11__N_236[0]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i1_3_lut (.A(\LOCosine[1] ), .B(MixerOutCos_11__N_250[0]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i1_3_lut.init = 16'hcaca;
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module SinCos
//

module SinCos (osc_clk, VCC_net, GND_net, \phase_accum[57] , \phase_accum[58] , 
            \phase_accum[59] , \phase_accum[60] , \phase_accum[61] , \phase_accum[62] , 
            \phase_accum[63] , \LOSine[1] , \LOSine[2] , \LOSine[3] , 
            \LOSine[4] , \LOSine[5] , \LOSine[6] , \LOSine[7] , \LOSine[8] , 
            \LOSine[9] , \LOSine[10] , \LOSine[11] , \LOSine[12] , \LOCosine[1] , 
            \LOCosine[2] , \LOCosine[3] , \LOCosine[4] , \LOCosine[5] , 
            \LOCosine[6] , \LOCosine[7] , \LOCosine[8] , \LOCosine[9] , 
            \LOCosine[10] , \LOCosine[11] , \LOCosine[12] , \phase_accum[56] ) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input osc_clk;
    input VCC_net;
    input GND_net;
    input \phase_accum[57] ;
    input \phase_accum[58] ;
    input \phase_accum[59] ;
    input \phase_accum[60] ;
    input \phase_accum[61] ;
    input \phase_accum[62] ;
    input \phase_accum[63] ;
    output \LOSine[1] ;
    output \LOSine[2] ;
    output \LOSine[3] ;
    output \LOSine[4] ;
    output \LOSine[5] ;
    output \LOSine[6] ;
    output \LOSine[7] ;
    output \LOSine[8] ;
    output \LOSine[9] ;
    output \LOSine[10] ;
    output \LOSine[11] ;
    output \LOSine[12] ;
    output \LOCosine[1] ;
    output \LOCosine[2] ;
    output \LOCosine[3] ;
    output \LOCosine[4] ;
    output \LOCosine[5] ;
    output \LOCosine[6] ;
    output \LOCosine[7] ;
    output \LOCosine[8] ;
    output \LOCosine[9] ;
    output \LOCosine[10] ;
    output \LOCosine[11] ;
    output \LOCosine[12] ;
    input \phase_accum[56] ;
    
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(69[8:15])
    
    wire rom_addr0_r_1, rom_addr0_r_1_inv, rom_addr0_r_2, rom_addr0_r_3, 
        rom_addr0_r_4, rom_addr0_r_5, mx_ctrl_r, mx_ctrl_r_1, rom_addr0_r, 
        rom_addr0_r_n, rom_addr0_r_6, rom_dout_11, rom_dout_11_ffin, 
        rom_dout_10, rom_dout_10_ffin, rom_dout_9, rom_dout_9_ffin, 
        rom_dout_8, rom_dout_8_ffin, rom_dout_7, rom_dout_7_ffin, rom_dout_6, 
        rom_dout_6_ffin, rom_dout_5, rom_dout_5_ffin, rom_dout_4, rom_dout_4_ffin, 
        rom_dout_3, rom_dout_3_ffin, rom_dout_2, rom_dout_2_ffin, rom_dout_1, 
        rom_dout_1_ffin, rom_dout, rom_dout_ffin, rom_dout_25, rom_dout_25_ffin, 
        rom_dout_24, rom_dout_24_ffin, rom_dout_23, rom_dout_23_ffin, 
        rom_dout_22, rom_dout_22_ffin, rom_dout_21, rom_dout_21_ffin, 
        rom_dout_20, rom_dout_20_ffin, rom_dout_19, rom_dout_19_ffin, 
        rom_dout_18, rom_dout_18_ffin, rom_dout_17, rom_dout_17_ffin, 
        rom_dout_16, rom_dout_16_ffin, rom_dout_15, rom_dout_15_ffin, 
        rom_dout_14, rom_dout_14_ffin, rom_dout_13, rom_dout_13_ffin, 
        cosromoutsel_i, cosromoutsel, sinromoutsel, sinout_pre_1, sinout_pre_2, 
        sinout_pre_3, sinout_pre_4, sinout_pre_5, sinout_pre_6, sinout_pre_7, 
        sinout_pre_8, sinout_pre_9, sinout_pre_10, sinout_pre_11, sinout_pre_12, 
        cosout_pre_1, cosout_pre_2, cosout_pre_3, cosout_pre_4, cosout_pre_5, 
        cosout_pre_6, cosout_pre_7, cosout_pre_8, cosout_pre_9, cosout_pre_10, 
        cosout_pre_11, cosout_pre_12, rom_addr0_r_inv, co0, rom_addr0_r_n_1, 
        rom_addr0_r_n_2, rom_addr0_r_2_inv, co1, rom_addr0_r_n_3, rom_addr0_r_n_4, 
        rom_addr0_r_3_inv, rom_addr0_r_4_inv, co2, rom_addr0_r_n_5, 
        rom_addr0_r_5_inv, rom_dout_12_ffin, rom_addr0_r_7, rom_addr0_r_8, 
        rom_addr0_r_9, rom_addr0_r_10, rom_addr0_r_11, rom_dout_s_n_1, 
        rom_dout_s_n_2, co0_1, rom_dout_1_inv, rom_dout_2_inv, co1_1, 
        rom_dout_s_n_3, rom_dout_s_n_4, rom_dout_3_inv, rom_dout_4_inv, 
        co2_1, rom_dout_s_n_5, rom_dout_s_n_6, rom_dout_5_inv, rom_dout_6_inv, 
        co3, rom_dout_s_n_7, rom_dout_s_n_8, rom_dout_7_inv, rom_dout_8_inv, 
        co4, rom_dout_s_n_9, rom_dout_s_n_10, rom_dout_9_inv, rom_dout_10_inv, 
        co5, rom_dout_s_n_11, rom_dout_s_n_12, rom_dout_11_inv, rom_dout_12_inv, 
        rom_dout_13_inv, co0_2, rom_dout_c_n_1, rom_dout_c_n_2, rom_dout_14_inv, 
        rom_dout_15_inv, co1_2, rom_dout_c_n_3, rom_dout_c_n_4, rom_dout_16_inv, 
        rom_dout_17_inv, co2_2, rom_dout_c_n_5, rom_dout_c_n_6, rom_dout_18_inv, 
        rom_dout_19_inv, co3_1, rom_dout_c_n_7, rom_dout_c_n_8, rom_dout_20_inv, 
        rom_dout_21_inv, co4_1, rom_dout_c_n_9, rom_dout_c_n_10, rom_dout_22_inv, 
        rom_dout_23_inv, co5_1, rom_dout_c_n_11, rom_dout_c_n_12, rom_dout_24_inv, 
        rom_dout_25_inv, rom_dout_12, rom_dout_inv, func_or_inet, lx_ne0, 
        lx_ne0_inv, out_sel_i, rom_dout_s_1, rom_dout_s_2, rom_dout_s_3, 
        rom_dout_s_4, rom_dout_s_5, rom_dout_s_6, rom_dout_s_7, rom_dout_s_8, 
        rom_dout_s_9, rom_dout_s_10, rom_dout_s_11, rom_dout_s_12, rom_dout_c_1, 
        rom_dout_c_2, rom_dout_c_3, rom_dout_c_4, rom_dout_c_5, rom_dout_c_6, 
        rom_dout_c_7, rom_dout_c_8, rom_dout_c_9, rom_dout_c_10, rom_dout_c_11, 
        rom_dout_c_12, out_sel;
    
    INV INV_29 (.A(rom_addr0_r_1), .Z(rom_addr0_r_1_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    FD1P3DX FF_61 (.D(\phase_accum[57] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(rom_addr0_r_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(312[13:88])
    defparam FF_61.GSR = "ENABLED";
    FD1P3DX FF_60 (.D(\phase_accum[58] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(rom_addr0_r_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(315[13:88])
    defparam FF_60.GSR = "ENABLED";
    FD1P3DX FF_59 (.D(\phase_accum[59] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(rom_addr0_r_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(318[13:88])
    defparam FF_59.GSR = "ENABLED";
    FD1P3DX FF_58 (.D(\phase_accum[60] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(rom_addr0_r_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(321[13:88])
    defparam FF_58.GSR = "ENABLED";
    FD1P3DX FF_57 (.D(\phase_accum[61] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(rom_addr0_r_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(324[13:88])
    defparam FF_57.GSR = "ENABLED";
    FD1P3DX FF_56 (.D(\phase_accum[62] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(mx_ctrl_r)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(327[13:84])
    defparam FF_56.GSR = "ENABLED";
    FD1P3DX FF_55 (.D(\phase_accum[63] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(mx_ctrl_r_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(330[13:86])
    defparam FF_55.GSR = "ENABLED";
    MUX21 muxb_57 (.D0(rom_addr0_r), .D1(rom_addr0_r_n), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    FD1P3DX FF_53 (.D(rom_dout_11_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(355[13] 356[25])
    defparam FF_53.GSR = "ENABLED";
    FD1P3DX FF_52 (.D(rom_dout_10_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(359[13] 360[25])
    defparam FF_52.GSR = "ENABLED";
    FD1P3DX FF_51 (.D(rom_dout_9_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(363[13] 364[24])
    defparam FF_51.GSR = "ENABLED";
    FD1P3DX FF_50 (.D(rom_dout_8_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(367[13] 368[24])
    defparam FF_50.GSR = "ENABLED";
    FD1P3DX FF_49 (.D(rom_dout_7_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(371[13] 372[24])
    defparam FF_49.GSR = "ENABLED";
    FD1P3DX FF_48 (.D(rom_dout_6_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(375[13] 376[24])
    defparam FF_48.GSR = "ENABLED";
    FD1P3DX FF_47 (.D(rom_dout_5_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(379[13] 380[24])
    defparam FF_47.GSR = "ENABLED";
    FD1P3DX FF_46 (.D(rom_dout_4_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(383[13] 384[24])
    defparam FF_46.GSR = "ENABLED";
    FD1P3DX FF_45 (.D(rom_dout_3_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(387[13] 388[24])
    defparam FF_45.GSR = "ENABLED";
    FD1P3DX FF_44 (.D(rom_dout_2_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(391[13] 392[24])
    defparam FF_44.GSR = "ENABLED";
    FD1P3DX FF_43 (.D(rom_dout_1_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(395[13] 396[24])
    defparam FF_43.GSR = "ENABLED";
    FD1P3DX FF_42 (.D(rom_dout_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(399[13] 400[22])
    defparam FF_42.GSR = "ENABLED";
    FD1P3DX FF_41 (.D(rom_dout_25_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_25)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(403[13] 404[25])
    defparam FF_41.GSR = "ENABLED";
    FD1P3DX FF_40 (.D(rom_dout_24_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_24)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(407[13] 408[25])
    defparam FF_40.GSR = "ENABLED";
    FD1P3DX FF_39 (.D(rom_dout_23_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_23)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(411[13] 412[25])
    defparam FF_39.GSR = "ENABLED";
    FD1P3DX FF_38 (.D(rom_dout_22_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_22)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(415[13] 416[25])
    defparam FF_38.GSR = "ENABLED";
    FD1P3DX FF_37 (.D(rom_dout_21_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(419[13] 420[25])
    defparam FF_37.GSR = "ENABLED";
    FD1P3DX FF_36 (.D(rom_dout_20_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(423[13] 424[25])
    defparam FF_36.GSR = "ENABLED";
    FD1P3DX FF_35 (.D(rom_dout_19_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(427[13] 428[25])
    defparam FF_35.GSR = "ENABLED";
    FD1P3DX FF_34 (.D(rom_dout_18_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(431[13] 432[25])
    defparam FF_34.GSR = "ENABLED";
    FD1P3DX FF_33 (.D(rom_dout_17_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(435[13] 436[25])
    defparam FF_33.GSR = "ENABLED";
    FD1P3DX FF_32 (.D(rom_dout_16_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(439[13] 440[25])
    defparam FF_32.GSR = "ENABLED";
    FD1P3DX FF_31 (.D(rom_dout_15_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(443[13] 444[25])
    defparam FF_31.GSR = "ENABLED";
    FD1P3DX FF_30 (.D(rom_dout_14_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(447[13] 448[25])
    defparam FF_30.GSR = "ENABLED";
    FD1P3DX FF_29 (.D(rom_dout_13_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(451[13] 452[25])
    defparam FF_29.GSR = "ENABLED";
    FD1P3DX FF_28 (.D(cosromoutsel_i), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(cosromoutsel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(455[13] 456[26])
    defparam FF_28.GSR = "ENABLED";
    FD1P3DX FF_27 (.D(mx_ctrl_r_1), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(sinromoutsel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(459[13] 460[26])
    defparam FF_27.GSR = "ENABLED";
    FD1P3DX FF_24 (.D(sinout_pre_1), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[1] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(599[13] 600[21])
    defparam FF_24.GSR = "ENABLED";
    FD1P3DX FF_23 (.D(sinout_pre_2), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[2] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(603[13] 604[21])
    defparam FF_23.GSR = "ENABLED";
    FD1P3DX FF_22 (.D(sinout_pre_3), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[3] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(607[13] 608[21])
    defparam FF_22.GSR = "ENABLED";
    FD1P3DX FF_21 (.D(sinout_pre_4), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[4] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(611[13] 612[21])
    defparam FF_21.GSR = "ENABLED";
    FD1P3DX FF_20 (.D(sinout_pre_5), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[5] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(615[13] 616[21])
    defparam FF_20.GSR = "ENABLED";
    FD1P3DX FF_19 (.D(sinout_pre_6), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[6] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(619[13] 620[21])
    defparam FF_19.GSR = "ENABLED";
    FD1P3DX FF_18 (.D(sinout_pre_7), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[7] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(623[13] 624[21])
    defparam FF_18.GSR = "ENABLED";
    FD1P3DX FF_17 (.D(sinout_pre_8), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[8] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(627[13] 628[21])
    defparam FF_17.GSR = "ENABLED";
    FD1P3DX FF_16 (.D(sinout_pre_9), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[9] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(631[13] 632[21])
    defparam FF_16.GSR = "ENABLED";
    FD1P3DX FF_15 (.D(sinout_pre_10), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[10] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(635[13] 636[22])
    defparam FF_15.GSR = "ENABLED";
    FD1P3DX FF_14 (.D(sinout_pre_11), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[11] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(639[13] 640[22])
    defparam FF_14.GSR = "ENABLED";
    FD1P3DX FF_13 (.D(sinout_pre_12), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[12] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(643[13] 644[22])
    defparam FF_13.GSR = "ENABLED";
    FD1P3DX FF_11 (.D(cosout_pre_1), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[1] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(650[13] 651[23])
    defparam FF_11.GSR = "ENABLED";
    FD1P3DX FF_10 (.D(cosout_pre_2), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[2] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(654[13] 655[23])
    defparam FF_10.GSR = "ENABLED";
    FD1P3DX FF_9 (.D(cosout_pre_3), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[3] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(658[13] 659[23])
    defparam FF_9.GSR = "ENABLED";
    FD1P3DX FF_8 (.D(cosout_pre_4), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[4] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(662[13] 663[23])
    defparam FF_8.GSR = "ENABLED";
    FD1P3DX FF_7 (.D(cosout_pre_5), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[5] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(666[13] 667[23])
    defparam FF_7.GSR = "ENABLED";
    FD1P3DX FF_6 (.D(cosout_pre_6), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[6] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(670[13] 671[23])
    defparam FF_6.GSR = "ENABLED";
    FD1P3DX FF_5 (.D(cosout_pre_7), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[7] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(674[13] 675[23])
    defparam FF_5.GSR = "ENABLED";
    FD1P3DX FF_4 (.D(cosout_pre_8), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[8] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(678[13] 679[23])
    defparam FF_4.GSR = "ENABLED";
    FD1P3DX FF_3 (.D(cosout_pre_9), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[9] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(682[13] 683[23])
    defparam FF_3.GSR = "ENABLED";
    FD1P3DX FF_2 (.D(cosout_pre_10), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[10] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(686[13] 687[24])
    defparam FF_2.GSR = "ENABLED";
    FD1P3DX FF_1 (.D(cosout_pre_11), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[11] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(690[13] 691[24])
    defparam FF_1.GSR = "ENABLED";
    FD1P3DX FF_0 (.D(cosout_pre_12), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[12] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(694[13] 695[24])
    defparam FF_0.GSR = "ENABLED";
    FADD2B neg_rom_addr0_r_n_0 (.A0(GND_net), .A1(rom_addr0_r_inv), .B0(GND_net), 
           .B1(VCC_net), .CI(GND_net), .COUT(co0), .S1(rom_addr0_r_n)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    FADD2B neg_rom_addr0_r_n_1 (.A0(rom_addr0_r_1_inv), .A1(rom_addr0_r_2_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co0), .COUT(co1), .S0(rom_addr0_r_n_1), 
           .S1(rom_addr0_r_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    FADD2B neg_rom_addr0_r_n_2 (.A0(rom_addr0_r_3_inv), .A1(rom_addr0_r_4_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co1), .COUT(co2), .S0(rom_addr0_r_n_3), 
           .S1(rom_addr0_r_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    FADD2B neg_rom_addr0_r_n_3 (.A0(rom_addr0_r_5_inv), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co2), .S0(rom_addr0_r_n_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    ROM64X1A triglut_1_0_25 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_12_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_25.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    FADD2B neg_rom_dout_s_n_1 (.A0(rom_dout_1_inv), .A1(rom_dout_2_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co0_1), .COUT(co1_1), .S0(rom_dout_s_n_1), 
           .S1(rom_dout_s_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    FADD2B neg_rom_dout_s_n_2 (.A0(rom_dout_3_inv), .A1(rom_dout_4_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co1_1), .COUT(co2_1), .S0(rom_dout_s_n_3), 
           .S1(rom_dout_s_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    FADD2B neg_rom_dout_s_n_3 (.A0(rom_dout_5_inv), .A1(rom_dout_6_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co2_1), .COUT(co3), .S0(rom_dout_s_n_5), 
           .S1(rom_dout_s_n_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    FADD2B neg_rom_dout_s_n_4 (.A0(rom_dout_7_inv), .A1(rom_dout_8_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co3), .COUT(co4), .S0(rom_dout_s_n_7), 
           .S1(rom_dout_s_n_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    FADD2B neg_rom_dout_s_n_5 (.A0(rom_dout_9_inv), .A1(rom_dout_10_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co4), .COUT(co5), .S0(rom_dout_s_n_9), 
           .S1(rom_dout_s_n_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    FADD2B neg_rom_dout_s_n_6 (.A0(rom_dout_11_inv), .A1(rom_dout_12_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co5), .S0(rom_dout_s_n_11), 
           .S1(rom_dout_s_n_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_30 (.A(rom_addr0_r_2), .Z(rom_addr0_r_2_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    FADD2B neg_rom_dout_c_n_0 (.A0(GND_net), .A1(rom_dout_13_inv), .B0(GND_net), 
           .B1(VCC_net), .CI(GND_net), .COUT(co0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    FADD2B neg_rom_dout_c_n_1 (.A0(rom_dout_14_inv), .A1(rom_dout_15_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co0_2), .COUT(co1_2), .S0(rom_dout_c_n_1), 
           .S1(rom_dout_c_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    FADD2B neg_rom_dout_c_n_2 (.A0(rom_dout_16_inv), .A1(rom_dout_17_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co1_2), .COUT(co2_2), .S0(rom_dout_c_n_3), 
           .S1(rom_dout_c_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    FADD2B neg_rom_dout_c_n_3 (.A0(rom_dout_18_inv), .A1(rom_dout_19_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co2_2), .COUT(co3_1), .S0(rom_dout_c_n_5), 
           .S1(rom_dout_c_n_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    FADD2B neg_rom_dout_c_n_4 (.A0(rom_dout_20_inv), .A1(rom_dout_21_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co3_1), .COUT(co4_1), .S0(rom_dout_c_n_7), 
           .S1(rom_dout_c_n_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    FADD2B neg_rom_dout_c_n_5 (.A0(rom_dout_22_inv), .A1(rom_dout_23_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co4_1), .COUT(co5_1), .S0(rom_dout_c_n_9), 
           .S1(rom_dout_c_n_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    FADD2B neg_rom_dout_c_n_6 (.A0(rom_dout_24_inv), .A1(rom_dout_25_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co5_1), .S0(rom_dout_c_n_11), 
           .S1(rom_dout_c_n_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_31 (.A(rom_addr0_r_3), .Z(rom_addr0_r_3_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_32 (.A(rom_addr0_r_4), .Z(rom_addr0_r_4_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_33 (.A(rom_addr0_r_5), .Z(rom_addr0_r_5_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_28 (.A(rom_addr0_r), .Z(rom_addr0_r_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    XOR2 XOR2_t1 (.A(mx_ctrl_r), .B(mx_ctrl_r_1), .Z(cosromoutsel_i)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(241[10:70])
    INV INV_27 (.A(rom_dout_12), .Z(rom_dout_12_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_26 (.A(rom_dout_11), .Z(rom_dout_11_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_25 (.A(rom_dout_10), .Z(rom_dout_10_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_24 (.A(rom_dout_9), .Z(rom_dout_9_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_23 (.A(rom_dout_8), .Z(rom_dout_8_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_22 (.A(rom_dout_7), .Z(rom_dout_7_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_21 (.A(rom_dout_6), .Z(rom_dout_6_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_20 (.A(rom_dout_5), .Z(rom_dout_5_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_19 (.A(rom_dout_4), .Z(rom_dout_4_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_18 (.A(rom_dout_3), .Z(rom_dout_3_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_17 (.A(rom_dout_2), .Z(rom_dout_2_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_16 (.A(rom_dout_1), .Z(rom_dout_1_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_15 (.A(rom_dout), .Z(rom_dout_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_14 (.A(rom_dout_25), .Z(rom_dout_25_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_13 (.A(rom_dout_24), .Z(rom_dout_24_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_12 (.A(rom_dout_23), .Z(rom_dout_23_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_11 (.A(rom_dout_22), .Z(rom_dout_22_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_10 (.A(rom_dout_21), .Z(rom_dout_21_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_9 (.A(rom_dout_20), .Z(rom_dout_20_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_8 (.A(rom_dout_19), .Z(rom_dout_19_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_7 (.A(rom_dout_18), .Z(rom_dout_18_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_6 (.A(rom_dout_17), .Z(rom_dout_17_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_5 (.A(rom_dout_16), .Z(rom_dout_16_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_4 (.A(rom_dout_15), .Z(rom_dout_15_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_3 (.A(rom_dout_14), .Z(rom_dout_14_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    INV INV_2 (.A(rom_dout_13), .Z(rom_dout_13_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    ROM16X1A LUT4_1 (.AD0(rom_addr0_r_9), .AD1(rom_addr0_r_8), .AD2(rom_addr0_r_7), 
            .AD3(rom_addr0_r_6), .DO0(func_or_inet)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam LUT4_1.initval = 16'b1111111111111110;
    ROM16X1A LUT4_0 (.AD0(GND_net), .AD1(rom_addr0_r_11), .AD2(rom_addr0_r_10), 
            .AD3(func_or_inet), .DO0(lx_ne0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam LUT4_0.initval = 16'b1111111111111110;
    INV INV_1 (.A(lx_ne0), .Z(lx_ne0_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    AND2 AND2_t0 (.A(mx_ctrl_r), .B(lx_ne0_inv), .Z(out_sel_i)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(305[10:64])
    FD1P3DX FF_62 (.D(\phase_accum[56] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(rom_addr0_r)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(309[13:86])
    defparam FF_62.GSR = "ENABLED";
    MUX21 muxb_56 (.D0(rom_addr0_r_1), .D1(rom_addr0_r_n_1), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_55 (.D0(rom_addr0_r_2), .D1(rom_addr0_r_n_2), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_54 (.D0(rom_addr0_r_3), .D1(rom_addr0_r_n_3), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_53 (.D0(rom_addr0_r_4), .D1(rom_addr0_r_n_4), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_52 (.D0(rom_addr0_r_5), .D1(rom_addr0_r_n_5), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    FD1P3DX FF_54 (.D(rom_dout_12_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(351[13] 352[25])
    defparam FF_54.GSR = "ENABLED";
    MUX21 muxb_50 (.D0(rom_dout_1), .D1(rom_dout_s_n_1), .SD(sinromoutsel), 
          .Z(rom_dout_s_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_49 (.D0(rom_dout_2), .D1(rom_dout_s_n_2), .SD(sinromoutsel), 
          .Z(rom_dout_s_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_48 (.D0(rom_dout_3), .D1(rom_dout_s_n_3), .SD(sinromoutsel), 
          .Z(rom_dout_s_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_47 (.D0(rom_dout_4), .D1(rom_dout_s_n_4), .SD(sinromoutsel), 
          .Z(rom_dout_s_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_46 (.D0(rom_dout_5), .D1(rom_dout_s_n_5), .SD(sinromoutsel), 
          .Z(rom_dout_s_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_45 (.D0(rom_dout_6), .D1(rom_dout_s_n_6), .SD(sinromoutsel), 
          .Z(rom_dout_s_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_44 (.D0(rom_dout_7), .D1(rom_dout_s_n_7), .SD(sinromoutsel), 
          .Z(rom_dout_s_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_43 (.D0(rom_dout_8), .D1(rom_dout_s_n_8), .SD(sinromoutsel), 
          .Z(rom_dout_s_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_42 (.D0(rom_dout_9), .D1(rom_dout_s_n_9), .SD(sinromoutsel), 
          .Z(rom_dout_s_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_41 (.D0(rom_dout_10), .D1(rom_dout_s_n_10), .SD(sinromoutsel), 
          .Z(rom_dout_s_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_40 (.D0(rom_dout_11), .D1(rom_dout_s_n_11), .SD(sinromoutsel), 
          .Z(rom_dout_s_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_39 (.D0(rom_dout_12), .D1(rom_dout_s_n_12), .SD(sinromoutsel), 
          .Z(rom_dout_s_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_37 (.D0(rom_dout_14), .D1(rom_dout_c_n_1), .SD(cosromoutsel), 
          .Z(rom_dout_c_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_36 (.D0(rom_dout_15), .D1(rom_dout_c_n_2), .SD(cosromoutsel), 
          .Z(rom_dout_c_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_35 (.D0(rom_dout_16), .D1(rom_dout_c_n_3), .SD(cosromoutsel), 
          .Z(rom_dout_c_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_34 (.D0(rom_dout_17), .D1(rom_dout_c_n_4), .SD(cosromoutsel), 
          .Z(rom_dout_c_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_33 (.D0(rom_dout_18), .D1(rom_dout_c_n_5), .SD(cosromoutsel), 
          .Z(rom_dout_c_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_32 (.D0(rom_dout_19), .D1(rom_dout_c_n_6), .SD(cosromoutsel), 
          .Z(rom_dout_c_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_31 (.D0(rom_dout_20), .D1(rom_dout_c_n_7), .SD(cosromoutsel), 
          .Z(rom_dout_c_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_30 (.D0(rom_dout_21), .D1(rom_dout_c_n_8), .SD(cosromoutsel), 
          .Z(rom_dout_c_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_29 (.D0(rom_dout_22), .D1(rom_dout_c_n_9), .SD(cosromoutsel), 
          .Z(rom_dout_c_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_28 (.D0(rom_dout_23), .D1(rom_dout_c_n_10), .SD(cosromoutsel), 
          .Z(rom_dout_c_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_27 (.D0(rom_dout_24), .D1(rom_dout_c_n_11), .SD(cosromoutsel), 
          .Z(rom_dout_c_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_26 (.D0(rom_dout_25), .D1(rom_dout_c_n_12), .SD(cosromoutsel), 
          .Z(rom_dout_c_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    FD1P3DX FF_26 (.D(out_sel_i), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(out_sel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(541[13:83])
    defparam FF_26.GSR = "ENABLED";
    MUX21 muxb_24 (.D0(rom_dout_s_1), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_23 (.D0(rom_dout_s_2), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_22 (.D0(rom_dout_s_3), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_21 (.D0(rom_dout_s_4), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_20 (.D0(rom_dout_s_5), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_19 (.D0(rom_dout_s_6), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_18 (.D0(rom_dout_s_7), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_17 (.D0(rom_dout_s_8), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_16 (.D0(rom_dout_s_9), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_15 (.D0(rom_dout_s_10), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_14 (.D0(rom_dout_s_11), .D1(VCC_net), .SD(out_sel), .Z(sinout_pre_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_13 (.D0(rom_dout_s_12), .D1(mx_ctrl_r_1), .SD(out_sel), 
          .Z(sinout_pre_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_11 (.D0(rom_dout_c_1), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_10 (.D0(rom_dout_c_2), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_9 (.D0(rom_dout_c_3), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_8 (.D0(rom_dout_c_4), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_7 (.D0(rom_dout_c_5), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_6 (.D0(rom_dout_c_6), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_5 (.D0(rom_dout_c_7), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_4 (.D0(rom_dout_c_8), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_3 (.D0(rom_dout_c_9), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_2 (.D0(rom_dout_c_10), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_1 (.D0(rom_dout_c_11), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    MUX21 muxb_0 (.D0(rom_dout_c_12), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    ROM64X1A triglut_1_0_24 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_11_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_24.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    ROM64X1A triglut_1_0_23 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_10_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_23.initval = 64'b1111111111111111111111111111111111111111110000000000000000000000;
    ROM64X1A triglut_1_0_22 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_9_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_22.initval = 64'b1111111111111111111111111111100000000000001111111111100000000000;
    ROM64X1A triglut_1_0_21 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_8_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_21.initval = 64'b1111111111111111111100000000011111110000001111110000011111000000;
    ROM64X1A triglut_1_0_20 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_7_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_20.initval = 64'b1111111111111100000011111000011110001110001110001110011100111000;
    ROM64X1A triglut_1_0_19 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_6_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_19.initval = 64'b1111111111000011100011100110011001001101101101001001011010110100;
    ROM64X1A triglut_1_0_18 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_5_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_18.initval = 64'b1111111000110011011010010101010100101001001001101100110001100110;
    ROM64X1A triglut_1_0_17 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_4_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_17.initval = 64'b1111100100101010110011000000000001110011011010110101010110101010;
    ROM64X1A triglut_1_0_16 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_3_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_16.initval = 64'b1110010110011100010101001111111101101010110011100000000011110000;
    ROM64X1A triglut_1_0_15 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_2_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_15.initval = 64'b1101000010100011001111010111110011001100010101100000000011001100;
    ROM64X1A triglut_1_0_14 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_1_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_14.initval = 64'b1111011011100010010110111011101001110011000000100111110010101010;
    ROM64X1A triglut_1_0_13 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_13.initval = 64'b1000100101001010011001010111111001010010011110001001001001111000;
    ROM64X1A triglut_1_0_12 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_25_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_12.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    ROM64X1A triglut_1_0_11 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_24_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_11.initval = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    ROM64X1A triglut_1_0_10 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_23_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_10.initval = 64'b0000000000000000000001111111111111111111111111111111111111111110;
    ROM64X1A triglut_1_0_9 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_22_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_9.initval = 64'b0000000000111111111110000000000000111111111111111111111111111110;
    ROM64X1A triglut_1_0_8 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_21_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_8.initval = 64'b0000011111000001111110000001111111000000000111111111111111111110;
    ROM64X1A triglut_1_0_7 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_20_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_7.initval = 64'b0011100111001110001110001110001111000011111000000111111111111110;
    ROM64X1A triglut_1_0_6 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_19_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_6.initval = 64'b0101101011010010010110110110010011001100111000111000011111111110;
    ROM64X1A triglut_1_0_5 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_18_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_5.initval = 64'b1100110001100110110010010010100101010101001011011001100011111110;
    ROM64X1A triglut_1_0_4 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_17_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_4.initval = 64'b1010101101010101101011011001110000000000011001101010100100111110;
    ROM64X1A triglut_1_0_3 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_16_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_3.initval = 64'b0001111000000000111001101010110111111110010101000111001101001110;
    ROM64X1A triglut_1_0_2 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_15_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_2.initval = 64'b0110011000000000110101000110011001111101011110011000101000010110;
    ROM64X1A triglut_1_0_1 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_14_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_1.initval = 64'b1010101001111100100000011001110010111011101101001000111011011110;
    ROM64X1A triglut_1_0_0 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_13_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    defparam triglut_1_0_0.initval = 64'b0011110010010010001111001001010011111101010011001010010100100010;
    FADD2B neg_rom_dout_s_n_0 (.A0(GND_net), .A1(rom_dout_inv), .B0(GND_net), 
           .B1(VCC_net), .CI(GND_net), .COUT(co0_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=148 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(141[8] 148[2])
    
endmodule
//
// Verilog Description of module \CIC(width=72,decimation_ratio=4096) 
//

module \CIC(width=72,decimation_ratio=4096)  (MixerOutSin, osc_clk, GND_net, 
            CIC1_out_clkSin, \CIC1_outSin[0] , \CICGain[0] , \CICGain[1] , 
            n62, \d10[60] , n63, \d_out_11__N_1819[2] , n64, \d_out_11__N_1819[3] , 
            n65, \d_out_11__N_1819[4] , n66, \d_out_11__N_1819[5] , 
            n67, \d_out_11__N_1819[6] , n68, \d_out_11__N_1819[7] , 
            \d10[68] , \d_out_11__N_1819[8] , n70, \d_out_11__N_1819[9] , 
            \d10[71] , \d_out_11__N_1819[11] , \CIC1_outSin[1] , \CIC1_outSin[2] , 
            \CIC1_outSin[3] , \CIC1_outSin[4] , \CIC1_outSin[5] , MYLED_c_0, 
            MYLED_c_1, MYLED_c_2, MYLED_c_3, MYLED_c_4, MYLED_c_5, 
            \d10[67] , \d10[69] , \d10[70] , \d10[65] , \d10[66] , 
            \d10[63] , \d_out_11__N_1819[10] , \d10[64] , \d10[61] , 
            \d10[62] , n61, \d10[59] ) /* synthesis syn_module_defined=1 */ ;
    input [11:0]MixerOutSin;
    input osc_clk;
    input GND_net;
    output CIC1_out_clkSin;
    output \CIC1_outSin[0] ;
    input \CICGain[0] ;
    input \CICGain[1] ;
    input n62;
    input \d10[60] ;
    input n63;
    output \d_out_11__N_1819[2] ;
    input n64;
    output \d_out_11__N_1819[3] ;
    input n65;
    output \d_out_11__N_1819[4] ;
    input n66;
    output \d_out_11__N_1819[5] ;
    input n67;
    output \d_out_11__N_1819[6] ;
    input n68;
    output \d_out_11__N_1819[7] ;
    input \d10[68] ;
    output \d_out_11__N_1819[8] ;
    input n70;
    output \d_out_11__N_1819[9] ;
    input \d10[71] ;
    output \d_out_11__N_1819[11] ;
    output \CIC1_outSin[1] ;
    output \CIC1_outSin[2] ;
    output \CIC1_outSin[3] ;
    output \CIC1_outSin[4] ;
    output \CIC1_outSin[5] ;
    output MYLED_c_0;
    output MYLED_c_1;
    output MYLED_c_2;
    output MYLED_c_3;
    output MYLED_c_4;
    output MYLED_c_5;
    input \d10[67] ;
    input \d10[69] ;
    input \d10[70] ;
    input \d10[65] ;
    input \d10[66] ;
    input \d10[63] ;
    output \d_out_11__N_1819[10] ;
    input \d10[64] ;
    input \d10[61] ;
    input \d10[62] ;
    input n61;
    input \d10[59] ;
    
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(69[8:15])
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(85[6:21])
    
    wire n11965;
    wire [71:0]d1;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(35[26:28])
    
    wire n4299;
    wire [35:0]n4300;
    wire [71:0]d1_71__N_418;
    
    wire n11966;
    wire [71:0]d_tmp;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(30[26:31])
    
    wire osc_clk_enable_141;
    wire [71:0]d5;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(39[26:28])
    wire [71:0]d_d_tmp;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(30[33:40])
    
    wire osc_clk_enable_69;
    wire [71:0]d2;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(36[26:28])
    wire [71:0]d2_71__N_490;
    
    wire n11540;
    wire [71:0]d9;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(46[26:28])
    wire [71:0]d_d9;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(46[30:34])
    wire [35:0]n5972;
    
    wire n11541;
    wire [71:0]d3;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(37[26:28])
    wire [71:0]d3_71__N_562;
    wire [71:0]d4;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(38[26:28])
    wire [71:0]d4_71__N_634;
    wire [71:0]d5_71__N_706;
    wire [71:0]d6;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(43[26:28])
    wire [71:0]d6_71__N_1459;
    wire [71:0]d_d6;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(43[30:34])
    
    wire n11532, n11533, d_clk_tmp, n8403, v_comb;
    wire [71:0]d7;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(44[26:28])
    wire [71:0]d7_71__N_1531;
    wire [71:0]d_d7;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(44[30:34])
    wire [71:0]d8;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(45[26:28])
    wire [71:0]d8_71__N_1603;
    wire [71:0]d_d8;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(45[30:34])
    wire [71:0]d9_71__N_1675;
    wire [71:0]d_out_11__N_1819;
    wire [15:0]count;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(50[14:19])
    wire [15:0]count_15__N_1442;
    wire [71:0]d10;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(47[26:29])
    
    wire n62_c, n16, n13069, n13070, n23, n132, n63_c, n11335, 
        n11336, n65_c, n135, n11964, n11963, n11962, n11961, n11960, 
        n11955;
    wire [35:0]n4452;
    
    wire n11954, n11953, n11952, n64_c, n11334, n11333, n11332, 
        n11331, n134, n17, n61_c, n131, n66_c, n19, osc_clk_enable_410, 
        n70_c, n140, osc_clk_enable_460, osc_clk_enable_310, n11587;
    wire [35:0]n5820;
    
    wire n11586, n11585, n11584, n11583, n11582, n11581, n11580, 
        n11579, n11578, n11577, n11576, n11575, n11574, n11573, 
        n11572, n11571, n11570, n11951, n132_adj_2488, osc_clk_enable_160, 
        n20, n11531, n11530, n68_c, n11529;
    wire [35:0]n6010;
    
    wire n11528, n11527, n11526, n11525, n11524, n11523, n11522, 
        n11521, n11520, n11539, n133, n24, n11519, n11518, n11517, 
        n13176, n11516, n136, n137, n11568, n5819, n11515, n21, 
        n16_adj_2489, n138, n11567, n11566, n11565, n11514, n131_adj_2491, 
        n11564, n11563, n11562, n11561, n11560, n11559, n11558, 
        n11557, n11513, n11556, n11512, n11555, n11554, n11553, 
        n11552, n11551, n11547, n11546, n11545, n11544, n21_adj_2495, 
        n26, n15, d_clk_tmp_N_1831, n11950, n133_adj_2497, n134_adj_2500, 
        n135_adj_2502, n136_adj_2505, n137_adj_2507, n11538, n138_adj_2511, 
        n11537, n8425;
    wire [15:0]n375;
    
    wire n140_adj_2514;
    wire [35:0]n4604;
    wire [35:0]n4756;
    
    wire osc_clk_enable_660, n11949, n11948, n11947, n11946, n11945, 
        n11944, n11943, n11942, n11941, n11940, n11939, osc_clk_enable_210, 
        osc_clk_enable_260, osc_clk_enable_360, osc_clk_enable_510, osc_clk_enable_560, 
        osc_clk_enable_610, osc_clk_enable_710;
    wire [71:0]d10_71__N_1747;
    
    wire n11936, n4451, n11935, n11934, n11933, n11932, n11931, 
        n11930, n11929, n11928, n11927, n11926, n11925, n11924, 
        n11923, n11922, n11536, n11921, n11920, n11919, n11914, 
        n11913, n11912, n11911, n11535, n11910, n11534, n11909, 
        n11908;
    wire [35:0]n4908;
    
    wire n11134;
    wire [35:0]n6884;
    
    wire n11133, n11132, n11131, n11130, n11129, n11128, n11127, 
        n11126, n11125, n11124, n11123, n11122, n11121, n11120, 
        n11119, n11118, n11117, n11115, n6883, n11114, n11113, 
        n11112, n11111, n11110, n11109, n11108, n11107, n11106, 
        n11105, n11104, n11103, n11102, n11101, n11100, n11099, 
        n11098, n11094;
    wire [35:0]n7036;
    
    wire n11093, n11092, n11091, n11090, n11089, n11088, n11087, 
        n11086, n11085, n11084, n11083, n11082, n11081, n11080, 
        n11079, n11078, n11077, n11075, n7035, n11074, n11073, 
        n11072, n11071, n11070, n11069, n11068, n11067, n11066, 
        n11065, n11064, n11063, n11062, n11061, n11060, n11059, 
        n11058, n10969, n4147, n10968, n10967, n10966, n10965, 
        n10964, n10963, n10962, n10961, n10960, n10959, n10958, 
        n10957, n10956, n10955, n10954, n10953, n10952, n10930, 
        n10929, n10928, n10927, n10926, n10925, n10924, n10923, 
        n10922, n10921, n10920, n10919, n10918, n10917, n10916, 
        n10915, n10914, n10913, n10806, n10805, n10804, n10803, 
        n10802, n10801, n10800, n10799, n10779, n4907, n10778, 
        n10777, n10776, n10775, n10774, n10773, n10772, n10771, 
        n10770, n10769, n10768, n10767, n10766, n10765, n10764, 
        n10763, n10762, n10760, n4755, n10759, n10758, n10757, 
        n10756, n10755, n10754, n10753, n10752, n10751, n10750, 
        n10749, n10748, n10747, n10746, n10745, n10744, n10743, 
        n10741, n4603, n10740, n10739, n10738, n10737, n10736, 
        n10735, n10734, n10733, n10732, n10731, n10730, n10729, 
        n10728, n10727, n10726, n10725, n10724, n10722, n10721, 
        n10720, n10719, n10718, n10717, n10716, n10715, n10714, 
        n10713, n10712, n10711, n10710, n10709, n10708, n10707, 
        n10706, n10705, n10660, n10659, n10658, n10657, n10656, 
        n10655, n10654, n10653, n10652, n10651, n10650, n10649, 
        n10648, n10647, n10646, n10645, n10644, n10643, n12131, 
        n12130, n12129, n12128, n12127, n12126, n12125, n12124, 
        n11484, n11483, n11482, n11481, n11480, n11479, n11478, 
        n11477, n11476, n11475, n11474, n11473, n11472, n11471, 
        n11470, n11469, n11468, n11467, n11348, n5971, n11347, 
        n11346, n11345, n11344, n11343, n11342, n11341, n11340, 
        n11339, n11338, n11337, n54, n12123, n12122, n12121, n12120, 
        n12119, n12118, n12117, n12116, n12115, n12114, n11907, 
        n11906, n11905, n11904, n11903, n11902, n11901, n11900, 
        n11899, n11898, n11895, n11894, n11893, n11892, n11891, 
        n11890, n11889, n11888, n11887, n11886, n11885, n11884, 
        n11883, n11882, n11881, n11880, n11879, n11878, n11873, 
        n11872, n11871, n11870, n11869, n11868, n11867, n11866, 
        n11865, n11864, n11863, n11862, n11861, n11860, n11859, 
        n11858, n11857, n11854, n11853, n11852, n11851, n13180, 
        n13075, n12037;
    wire [35:0]n4148;
    
    wire n11850, n13074, n12036, n12035, n12034, n11849, n11848, 
        n12033, n12032, n12031, n11847, n12030, n12029, n12028, 
        n11846, n11845, n12027, n12026, n12025, n11844, n12024, 
        n12023, n12022, n11843, n11842, n12021, n12020, n12018, 
        n12017, n12016, n12015, n12014, n12013, n12012, n12011, 
        n12010, n12009, n12008, n12007, n12006, n12005, n11841, 
        n12004, n12003, n12002, n12001, n11996, n11840, n11995, 
        n11994, n11993, n11992, n11991, n11839, n11990, n11989, 
        n11988, n11987, n13077, n11543, n11542, n13081, n13080, 
        n11986, n11985, n11984, n11983, n11982, n11981, n11980, 
        n11838, n13084, n11837, n13083, n11832, n13078, n11831, 
        n11830, n11829, n11828, n11827, n11826, n11825, n11824, 
        n11823, n11822, n25, n11821, n11820, n11819, n11818, n11817, 
        n11816, n11813, n11812, n11811, n11977, n11810, n11809, 
        n11976, n11975, n11808, n11807, n11806, n11805, n11804, 
        n11803, n11802, n11801, n11800, n11799, n11798, n11797, 
        n11796, n11974, n11973, n11972, n11971, n11970, n11969, 
        n11968, n11967;
    
    CCU2D add_1052_13 (.A0(d1[46]), .B0(n4299), .C0(n4300[10]), .D0(MixerOutSin[11]), 
          .A1(d1[47]), .B1(n4299), .C1(n4300[11]), .D1(MixerOutSin[11]), 
          .CIN(n11965), .COUT(n11966), .S0(d1_71__N_418[46]), .S1(d1_71__N_418[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1052_13.INIT0 = 16'h74b8;
    defparam add_1052_13.INIT1 = 16'h74b8;
    defparam add_1052_13.INJECT1_0 = "NO";
    defparam add_1052_13.INJECT1_1 = "NO";
    FD1P3AX d_tmp_i0_i0 (.D(d5[0]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i0 (.D(d_tmp[0]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i0.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i3 (.D(d5[3]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i2 (.D(d5[2]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i2.GSR = "ENABLED";
    FD1S3AX d2_i0 (.D(d2_71__N_490[0]), .CK(osc_clk), .Q(d2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i0.GSR = "ENABLED";
    CCU2D add_1106_23 (.A0(d9[57]), .B0(d_d9[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[58]), .B1(d_d9[58]), .C1(GND_net), .D1(GND_net), .CIN(n11540), 
          .COUT(n11541), .S0(n5972[21]), .S1(n5972[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1106_23.INIT0 = 16'h5999;
    defparam add_1106_23.INIT1 = 16'h5999;
    defparam add_1106_23.INJECT1_0 = "NO";
    defparam add_1106_23.INJECT1_1 = "NO";
    FD1S3AX d3_i0 (.D(d3_71__N_562[0]), .CK(osc_clk), .Q(d3[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i0.GSR = "ENABLED";
    FD1S3AX d4_i0 (.D(d4_71__N_634[0]), .CK(osc_clk), .Q(d4[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i0.GSR = "ENABLED";
    FD1S3AX d5_i0 (.D(d5_71__N_706[0]), .CK(osc_clk), .Q(d5[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i0.GSR = "ENABLED";
    FD1P3AX d6_i0_i0 (.D(d6_71__N_1459[0]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i0 (.D(d6[0]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i0.GSR = "ENABLED";
    CCU2D add_1106_7 (.A0(d9[41]), .B0(d_d9[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[42]), .B1(d_d9[42]), .C1(GND_net), .D1(GND_net), .CIN(n11532), 
          .COUT(n11533));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1106_7.INIT0 = 16'h5999;
    defparam add_1106_7.INIT1 = 16'h5999;
    defparam add_1106_7.INJECT1_0 = "NO";
    defparam add_1106_7.INJECT1_1 = "NO";
    FD1S3JX d_clk_tmp_65 (.D(n8403), .CK(osc_clk), .PD(osc_clk_enable_141), 
            .Q(d_clk_tmp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_clk_tmp_65.GSR = "ENABLED";
    FD1S3AX v_comb_66 (.D(osc_clk_enable_141), .CK(osc_clk), .Q(v_comb)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66.GSR = "ENABLED";
    FD1S3AX d_clk_67 (.D(d_clk_tmp), .CK(osc_clk), .Q(CIC1_out_clkSin)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_clk_67.GSR = "ENABLED";
    FD1P3AX d7_i0_i0 (.D(d7_71__N_1531[0]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i0 (.D(d7[0]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d8_i0_i0 (.D(d8_71__N_1603[0]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i0 (.D(d8[0]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d9_i0_i0 (.D(d9_71__N_1675[0]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i0 (.D(d9[0]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_out_i0_i0 (.D(d_out_11__N_1819[0]), .SP(osc_clk_enable_69), 
            .CK(osc_clk), .Q(\CIC1_outSin[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i0.GSR = "ENABLED";
    FD1S3AX d1_i0 (.D(d1_71__N_418[0]), .CK(osc_clk), .Q(d1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i0.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i1 (.D(d5[1]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i1.GSR = "ENABLED";
    FD1S3IX count__i0 (.D(count_15__N_1442[0]), .CK(osc_clk), .CD(osc_clk_enable_141), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i0.GSR = "ENABLED";
    LUT4 shift_right_31_i62_3_lut (.A(d10[61]), .B(d10[62]), .C(\CICGain[0] ), 
         .Z(n62_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i62_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut (.A(count[5]), .B(count[4]), .Z(n16)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i9_4_lut (.A(n13069), .B(count[6]), .C(n13070), .D(count[2]), 
         .Z(n23)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 shift_right_31_i132_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n62), .D(\d10[60] ), .Z(n132)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i132_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i63_3_lut (.A(d10[62]), .B(d10[63]), .C(\CICGain[0] ), 
         .Z(n63_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i63_3_lut.init = 16'hcaca;
    CCU2D add_1105_11 (.A0(d9[9]), .B0(d_d9[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[10]), .B1(d_d9[10]), .C1(GND_net), .D1(GND_net), .CIN(n11335), 
          .COUT(n11336));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1105_11.INIT0 = 16'h5999;
    defparam add_1105_11.INIT1 = 16'h5999;
    defparam add_1105_11.INJECT1_0 = "NO";
    defparam add_1105_11.INJECT1_1 = "NO";
    LUT4 shift_right_31_i135_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65_c), .D(d10[63]), .Z(n135)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i135_3_lut_4_lut.init = 16'hf960;
    CCU2D add_1052_11 (.A0(d1[44]), .B0(n4299), .C0(n4300[8]), .D0(MixerOutSin[11]), 
          .A1(d1[45]), .B1(n4299), .C1(n4300[9]), .D1(MixerOutSin[11]), 
          .CIN(n11964), .COUT(n11965), .S0(d1_71__N_418[44]), .S1(d1_71__N_418[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1052_11.INIT0 = 16'h74b8;
    defparam add_1052_11.INIT1 = 16'h74b8;
    defparam add_1052_11.INJECT1_0 = "NO";
    defparam add_1052_11.INJECT1_1 = "NO";
    CCU2D add_1052_9 (.A0(d1[42]), .B0(n4299), .C0(n4300[6]), .D0(MixerOutSin[11]), 
          .A1(d1[43]), .B1(n4299), .C1(n4300[7]), .D1(MixerOutSin[11]), 
          .CIN(n11963), .COUT(n11964), .S0(d1_71__N_418[42]), .S1(d1_71__N_418[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1052_9.INIT0 = 16'h74b8;
    defparam add_1052_9.INIT1 = 16'h74b8;
    defparam add_1052_9.INJECT1_0 = "NO";
    defparam add_1052_9.INJECT1_1 = "NO";
    CCU2D add_1052_7 (.A0(d1[40]), .B0(n4299), .C0(n4300[4]), .D0(MixerOutSin[11]), 
          .A1(d1[41]), .B1(n4299), .C1(n4300[5]), .D1(MixerOutSin[11]), 
          .CIN(n11962), .COUT(n11963), .S0(d1_71__N_418[40]), .S1(d1_71__N_418[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1052_7.INIT0 = 16'h74b8;
    defparam add_1052_7.INIT1 = 16'h74b8;
    defparam add_1052_7.INJECT1_0 = "NO";
    defparam add_1052_7.INJECT1_1 = "NO";
    CCU2D add_1052_5 (.A0(d1[38]), .B0(n4299), .C0(n4300[2]), .D0(MixerOutSin[11]), 
          .A1(d1[39]), .B1(n4299), .C1(n4300[3]), .D1(MixerOutSin[11]), 
          .CIN(n11961), .COUT(n11962), .S0(d1_71__N_418[38]), .S1(d1_71__N_418[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1052_5.INIT0 = 16'h74b8;
    defparam add_1052_5.INIT1 = 16'h74b8;
    defparam add_1052_5.INJECT1_0 = "NO";
    defparam add_1052_5.INJECT1_1 = "NO";
    CCU2D add_1052_3 (.A0(d1[36]), .B0(n4299), .C0(n4300[0]), .D0(MixerOutSin[11]), 
          .A1(d1[37]), .B1(n4299), .C1(n4300[1]), .D1(MixerOutSin[11]), 
          .CIN(n11960), .COUT(n11961), .S0(d1_71__N_418[36]), .S1(d1_71__N_418[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1052_3.INIT0 = 16'h74b8;
    defparam add_1052_3.INIT1 = 16'h74b8;
    defparam add_1052_3.INJECT1_0 = "NO";
    defparam add_1052_3.INJECT1_1 = "NO";
    CCU2D add_1052_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n4299), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11960));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1052_1.INIT0 = 16'hF000;
    defparam add_1052_1.INIT1 = 16'h0555;
    defparam add_1052_1.INJECT1_0 = "NO";
    defparam add_1052_1.INJECT1_1 = "NO";
    CCU2D add_1056_36 (.A0(d1[70]), .B0(d2[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[71]), .B1(d2[71]), .C1(GND_net), .D1(GND_net), .CIN(n11955), 
          .S0(n4452[34]), .S1(n4452[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1056_36.INIT0 = 16'h5666;
    defparam add_1056_36.INIT1 = 16'h5666;
    defparam add_1056_36.INJECT1_0 = "NO";
    defparam add_1056_36.INJECT1_1 = "NO";
    CCU2D add_1056_34 (.A0(d1[68]), .B0(d2[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[69]), .B1(d2[69]), .C1(GND_net), .D1(GND_net), .CIN(n11954), 
          .COUT(n11955), .S0(n4452[32]), .S1(n4452[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1056_34.INIT0 = 16'h5666;
    defparam add_1056_34.INIT1 = 16'h5666;
    defparam add_1056_34.INJECT1_0 = "NO";
    defparam add_1056_34.INJECT1_1 = "NO";
    CCU2D add_1056_32 (.A0(d1[66]), .B0(d2[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[67]), .B1(d2[67]), .C1(GND_net), .D1(GND_net), .CIN(n11953), 
          .COUT(n11954), .S0(n4452[30]), .S1(n4452[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1056_32.INIT0 = 16'h5666;
    defparam add_1056_32.INIT1 = 16'h5666;
    defparam add_1056_32.INJECT1_0 = "NO";
    defparam add_1056_32.INJECT1_1 = "NO";
    CCU2D add_1056_30 (.A0(d1[64]), .B0(d2[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[65]), .B1(d2[65]), .C1(GND_net), .D1(GND_net), .CIN(n11952), 
          .COUT(n11953), .S0(n4452[28]), .S1(n4452[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1056_30.INIT0 = 16'h5666;
    defparam add_1056_30.INIT1 = 16'h5666;
    defparam add_1056_30.INJECT1_0 = "NO";
    defparam add_1056_30.INJECT1_1 = "NO";
    LUT4 shift_right_31_i64_3_lut (.A(d10[63]), .B(d10[64]), .C(\CICGain[0] ), 
         .Z(n64_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i64_3_lut.init = 16'hcaca;
    CCU2D add_1105_9 (.A0(d9[7]), .B0(d_d9[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[8]), .B1(d_d9[8]), .C1(GND_net), .D1(GND_net), .CIN(n11334), 
          .COUT(n11335));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1105_9.INIT0 = 16'h5999;
    defparam add_1105_9.INIT1 = 16'h5999;
    defparam add_1105_9.INJECT1_0 = "NO";
    defparam add_1105_9.INJECT1_1 = "NO";
    CCU2D add_1105_7 (.A0(d9[5]), .B0(d_d9[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[6]), .B1(d_d9[6]), .C1(GND_net), .D1(GND_net), .CIN(n11333), 
          .COUT(n11334));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1105_7.INIT0 = 16'h5999;
    defparam add_1105_7.INIT1 = 16'h5999;
    defparam add_1105_7.INJECT1_0 = "NO";
    defparam add_1105_7.INJECT1_1 = "NO";
    CCU2D add_1105_5 (.A0(d9[3]), .B0(d_d9[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[4]), .B1(d_d9[4]), .C1(GND_net), .D1(GND_net), .CIN(n11332), 
          .COUT(n11333));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1105_5.INIT0 = 16'h5999;
    defparam add_1105_5.INIT1 = 16'h5999;
    defparam add_1105_5.INJECT1_0 = "NO";
    defparam add_1105_5.INJECT1_1 = "NO";
    CCU2D add_1105_3 (.A0(d9[1]), .B0(d_d9[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[2]), .B1(d_d9[2]), .C1(GND_net), .D1(GND_net), .CIN(n11331), 
          .COUT(n11332));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1105_3.INIT0 = 16'h5999;
    defparam add_1105_3.INIT1 = 16'h5999;
    defparam add_1105_3.INJECT1_0 = "NO";
    defparam add_1105_3.INJECT1_1 = "NO";
    LUT4 shift_right_31_i65_3_lut (.A(d10[64]), .B(d10[65]), .C(\CICGain[0] ), 
         .Z(n65_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i65_3_lut.init = 16'hcaca;
    CCU2D add_1105_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d9[0]), .B1(d_d9[0]), .C1(GND_net), .D1(GND_net), .COUT(n11331));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1105_1.INIT0 = 16'h0000;
    defparam add_1105_1.INIT1 = 16'h5999;
    defparam add_1105_1.INJECT1_0 = "NO";
    defparam add_1105_1.INJECT1_1 = "NO";
    LUT4 shift_right_31_i134_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64_c), .D(d10[62]), .Z(n134)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i134_3_lut_4_lut.init = 16'hf960;
    LUT4 i3_2_lut (.A(count[10]), .B(count[0]), .Z(n17)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    LUT4 shift_right_31_i131_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n61_c), .D(d10[59]), .Z(n131)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i131_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i66_3_lut (.A(d10[65]), .B(d10[66]), .C(\CICGain[0] ), 
         .Z(n66_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i66_3_lut.init = 16'hcaca;
    LUT4 i5_2_lut (.A(count[4]), .B(count[11]), .Z(n19)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i5_2_lut.init = 16'hbbbb;
    LUT4 i4658_2_lut (.A(MixerOutSin[11]), .B(d1[36]), .Z(n4300[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4658_2_lut.init = 16'h6666;
    FD1S3AX v_comb_66_rep_108 (.D(osc_clk_enable_141), .CK(osc_clk), .Q(osc_clk_enable_410)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_108.GSR = "ENABLED";
    LUT4 shift_right_31_i140_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n70_c), .D(d10[68]), .Z(n140)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i140_3_lut_4_lut.init = 16'hf960;
    FD1P3AX d_tmp_i0_i4 (.D(d5[4]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i15 (.D(d5[15]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i15.GSR = "ENABLED";
    LUT4 shift_right_31_i203_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63_c), .D(n131), .Z(d_out_11__N_1819[2])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i203_3_lut_4_lut.init = 16'hfe10;
    FD1S3AX v_comb_66_rep_109 (.D(osc_clk_enable_141), .CK(osc_clk), .Q(osc_clk_enable_460)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_109.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_106 (.D(osc_clk_enable_141), .CK(osc_clk), .Q(osc_clk_enable_310)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_106.GSR = "ENABLED";
    CCU2D add_1101_37 (.A0(d8[71]), .B0(d_d8[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11587), 
          .S0(n5820[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1101_37.INIT0 = 16'h5999;
    defparam add_1101_37.INIT1 = 16'h0000;
    defparam add_1101_37.INJECT1_0 = "NO";
    defparam add_1101_37.INJECT1_1 = "NO";
    CCU2D add_1101_35 (.A0(d8[69]), .B0(d_d8[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[70]), .B1(d_d8[70]), .C1(GND_net), .D1(GND_net), .CIN(n11586), 
          .COUT(n11587), .S0(n5820[33]), .S1(n5820[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1101_35.INIT0 = 16'h5999;
    defparam add_1101_35.INIT1 = 16'h5999;
    defparam add_1101_35.INJECT1_0 = "NO";
    defparam add_1101_35.INJECT1_1 = "NO";
    CCU2D add_1101_33 (.A0(d8[67]), .B0(d_d8[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[68]), .B1(d_d8[68]), .C1(GND_net), .D1(GND_net), .CIN(n11585), 
          .COUT(n11586), .S0(n5820[31]), .S1(n5820[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1101_33.INIT0 = 16'h5999;
    defparam add_1101_33.INIT1 = 16'h5999;
    defparam add_1101_33.INJECT1_0 = "NO";
    defparam add_1101_33.INJECT1_1 = "NO";
    CCU2D add_1101_31 (.A0(d8[65]), .B0(d_d8[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[66]), .B1(d_d8[66]), .C1(GND_net), .D1(GND_net), .CIN(n11584), 
          .COUT(n11585), .S0(n5820[29]), .S1(n5820[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1101_31.INIT0 = 16'h5999;
    defparam add_1101_31.INIT1 = 16'h5999;
    defparam add_1101_31.INJECT1_0 = "NO";
    defparam add_1101_31.INJECT1_1 = "NO";
    CCU2D add_1101_29 (.A0(d8[63]), .B0(d_d8[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[64]), .B1(d_d8[64]), .C1(GND_net), .D1(GND_net), .CIN(n11583), 
          .COUT(n11584), .S0(n5820[27]), .S1(n5820[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1101_29.INIT0 = 16'h5999;
    defparam add_1101_29.INIT1 = 16'h5999;
    defparam add_1101_29.INJECT1_0 = "NO";
    defparam add_1101_29.INJECT1_1 = "NO";
    CCU2D add_1101_27 (.A0(d8[61]), .B0(d_d8[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[62]), .B1(d_d8[62]), .C1(GND_net), .D1(GND_net), .CIN(n11582), 
          .COUT(n11583), .S0(n5820[25]), .S1(n5820[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1101_27.INIT0 = 16'h5999;
    defparam add_1101_27.INIT1 = 16'h5999;
    defparam add_1101_27.INJECT1_0 = "NO";
    defparam add_1101_27.INJECT1_1 = "NO";
    CCU2D add_1101_25 (.A0(d8[59]), .B0(d_d8[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[60]), .B1(d_d8[60]), .C1(GND_net), .D1(GND_net), .CIN(n11581), 
          .COUT(n11582), .S0(n5820[23]), .S1(n5820[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1101_25.INIT0 = 16'h5999;
    defparam add_1101_25.INIT1 = 16'h5999;
    defparam add_1101_25.INJECT1_0 = "NO";
    defparam add_1101_25.INJECT1_1 = "NO";
    CCU2D add_1101_23 (.A0(d8[57]), .B0(d_d8[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[58]), .B1(d_d8[58]), .C1(GND_net), .D1(GND_net), .CIN(n11580), 
          .COUT(n11581), .S0(n5820[21]), .S1(n5820[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1101_23.INIT0 = 16'h5999;
    defparam add_1101_23.INIT1 = 16'h5999;
    defparam add_1101_23.INJECT1_0 = "NO";
    defparam add_1101_23.INJECT1_1 = "NO";
    CCU2D add_1101_21 (.A0(d8[55]), .B0(d_d8[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[56]), .B1(d_d8[56]), .C1(GND_net), .D1(GND_net), .CIN(n11579), 
          .COUT(n11580), .S0(n5820[19]), .S1(n5820[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1101_21.INIT0 = 16'h5999;
    defparam add_1101_21.INIT1 = 16'h5999;
    defparam add_1101_21.INJECT1_0 = "NO";
    defparam add_1101_21.INJECT1_1 = "NO";
    CCU2D add_1101_19 (.A0(d8[53]), .B0(d_d8[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[54]), .B1(d_d8[54]), .C1(GND_net), .D1(GND_net), .CIN(n11578), 
          .COUT(n11579), .S0(n5820[17]), .S1(n5820[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1101_19.INIT0 = 16'h5999;
    defparam add_1101_19.INIT1 = 16'h5999;
    defparam add_1101_19.INJECT1_0 = "NO";
    defparam add_1101_19.INJECT1_1 = "NO";
    CCU2D add_1101_17 (.A0(d8[51]), .B0(d_d8[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[52]), .B1(d_d8[52]), .C1(GND_net), .D1(GND_net), .CIN(n11577), 
          .COUT(n11578), .S0(n5820[15]), .S1(n5820[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1101_17.INIT0 = 16'h5999;
    defparam add_1101_17.INIT1 = 16'h5999;
    defparam add_1101_17.INJECT1_0 = "NO";
    defparam add_1101_17.INJECT1_1 = "NO";
    CCU2D add_1101_15 (.A0(d8[49]), .B0(d_d8[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[50]), .B1(d_d8[50]), .C1(GND_net), .D1(GND_net), .CIN(n11576), 
          .COUT(n11577), .S0(n5820[13]), .S1(n5820[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1101_15.INIT0 = 16'h5999;
    defparam add_1101_15.INIT1 = 16'h5999;
    defparam add_1101_15.INJECT1_0 = "NO";
    defparam add_1101_15.INJECT1_1 = "NO";
    CCU2D add_1101_13 (.A0(d8[47]), .B0(d_d8[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[48]), .B1(d_d8[48]), .C1(GND_net), .D1(GND_net), .CIN(n11575), 
          .COUT(n11576), .S0(n5820[11]), .S1(n5820[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1101_13.INIT0 = 16'h5999;
    defparam add_1101_13.INIT1 = 16'h5999;
    defparam add_1101_13.INJECT1_0 = "NO";
    defparam add_1101_13.INJECT1_1 = "NO";
    CCU2D add_1101_11 (.A0(d8[45]), .B0(d_d8[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[46]), .B1(d_d8[46]), .C1(GND_net), .D1(GND_net), .CIN(n11574), 
          .COUT(n11575), .S0(n5820[9]), .S1(n5820[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1101_11.INIT0 = 16'h5999;
    defparam add_1101_11.INIT1 = 16'h5999;
    defparam add_1101_11.INJECT1_0 = "NO";
    defparam add_1101_11.INJECT1_1 = "NO";
    CCU2D add_1101_9 (.A0(d8[43]), .B0(d_d8[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[44]), .B1(d_d8[44]), .C1(GND_net), .D1(GND_net), .CIN(n11573), 
          .COUT(n11574), .S0(n5820[7]), .S1(n5820[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1101_9.INIT0 = 16'h5999;
    defparam add_1101_9.INIT1 = 16'h5999;
    defparam add_1101_9.INJECT1_0 = "NO";
    defparam add_1101_9.INJECT1_1 = "NO";
    CCU2D add_1101_7 (.A0(d8[41]), .B0(d_d8[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[42]), .B1(d_d8[42]), .C1(GND_net), .D1(GND_net), .CIN(n11572), 
          .COUT(n11573), .S0(n5820[5]), .S1(n5820[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1101_7.INIT0 = 16'h5999;
    defparam add_1101_7.INIT1 = 16'h5999;
    defparam add_1101_7.INJECT1_0 = "NO";
    defparam add_1101_7.INJECT1_1 = "NO";
    CCU2D add_1101_5 (.A0(d8[39]), .B0(d_d8[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[40]), .B1(d_d8[40]), .C1(GND_net), .D1(GND_net), .CIN(n11571), 
          .COUT(n11572), .S0(n5820[3]), .S1(n5820[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1101_5.INIT0 = 16'h5999;
    defparam add_1101_5.INIT1 = 16'h5999;
    defparam add_1101_5.INJECT1_0 = "NO";
    defparam add_1101_5.INJECT1_1 = "NO";
    CCU2D add_1101_3 (.A0(d8[37]), .B0(d_d8[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[38]), .B1(d_d8[38]), .C1(GND_net), .D1(GND_net), .CIN(n11570), 
          .COUT(n11571), .S0(n5820[1]), .S1(n5820[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1101_3.INIT0 = 16'h5999;
    defparam add_1101_3.INIT1 = 16'h5999;
    defparam add_1101_3.INJECT1_0 = "NO";
    defparam add_1101_3.INJECT1_1 = "NO";
    CCU2D add_1056_28 (.A0(d1[62]), .B0(d2[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[63]), .B1(d2[63]), .C1(GND_net), .D1(GND_net), .CIN(n11951), 
          .COUT(n11952), .S0(n4452[26]), .S1(n4452[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1056_28.INIT0 = 16'h5666;
    defparam add_1056_28.INIT1 = 16'h5666;
    defparam add_1056_28.INJECT1_0 = "NO";
    defparam add_1056_28.INJECT1_1 = "NO";
    LUT4 shift_right_31_i204_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64_c), .D(n132_adj_2488), .Z(d_out_11__N_1819[3])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i204_3_lut_4_lut.init = 16'hfe10;
    FD1P3AX d_d_tmp_i0_i71 (.D(d_tmp[71]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i70 (.D(d_tmp[70]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i69 (.D(d_tmp[69]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i68 (.D(d_tmp[68]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i67 (.D(d_tmp[67]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i66 (.D(d_tmp[66]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i65 (.D(d_tmp[65]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i64 (.D(d_tmp[64]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i63 (.D(d_tmp[63]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i62 (.D(d_tmp[62]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i61 (.D(d_tmp[61]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i60 (.D(d_tmp[60]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i59 (.D(d_tmp[59]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i58 (.D(d_tmp[58]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i57 (.D(d_tmp[57]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i56 (.D(d_tmp[56]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i55 (.D(d_tmp[55]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i54 (.D(d_tmp[54]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i53 (.D(d_tmp[53]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i52 (.D(d_tmp[52]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i51 (.D(d_tmp[51]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i50 (.D(d_tmp[50]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i49 (.D(d_tmp[49]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i48 (.D(d_tmp[48]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i47 (.D(d_tmp[47]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i46 (.D(d_tmp[46]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i45 (.D(d_tmp[45]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i44 (.D(d_tmp[44]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i43 (.D(d_tmp[43]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i42 (.D(d_tmp[42]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i41 (.D(d_tmp[41]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i40 (.D(d_tmp[40]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i39 (.D(d_tmp[39]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i38 (.D(d_tmp[38]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i37 (.D(d_tmp[37]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i36 (.D(d_tmp[36]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i35 (.D(d_tmp[35]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i34 (.D(d_tmp[34]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i33 (.D(d_tmp[33]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i32 (.D(d_tmp[32]), .SP(osc_clk_enable_69), .CK(osc_clk), 
            .Q(d_d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i25 (.D(d_tmp[25]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i24 (.D(d_tmp[24]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i23 (.D(d_tmp[23]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i22 (.D(d_tmp[22]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i21 (.D(d_tmp[21]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i20 (.D(d_tmp[20]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i19 (.D(d_tmp[19]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i26 (.D(d_tmp[26]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i27 (.D(d_tmp[27]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i27.GSR = "ENABLED";
    LUT4 i6_2_lut (.A(count[1]), .B(count[10]), .Z(n20)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    CCU2D add_1106_5 (.A0(d9[39]), .B0(d_d9[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[40]), .B1(d_d9[40]), .C1(GND_net), .D1(GND_net), .CIN(n11531), 
          .COUT(n11532));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1106_5.INIT0 = 16'h5999;
    defparam add_1106_5.INIT1 = 16'h5999;
    defparam add_1106_5.INJECT1_0 = "NO";
    defparam add_1106_5.INJECT1_1 = "NO";
    CCU2D add_1106_3 (.A0(d9[37]), .B0(d_d9[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[38]), .B1(d_d9[38]), .C1(GND_net), .D1(GND_net), .CIN(n11530), 
          .COUT(n11531));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1106_3.INIT0 = 16'h5999;
    defparam add_1106_3.INIT1 = 16'h5999;
    defparam add_1106_3.INJECT1_0 = "NO";
    defparam add_1106_3.INJECT1_1 = "NO";
    FD1P3AX d_d_tmp_i0_i28 (.D(d_tmp[28]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i28.GSR = "ENABLED";
    CCU2D add_1106_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d9[36]), .B1(d_d9[36]), .C1(GND_net), .D1(GND_net), .COUT(n11530));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1106_1.INIT0 = 16'hF000;
    defparam add_1106_1.INIT1 = 16'h5999;
    defparam add_1106_1.INJECT1_0 = "NO";
    defparam add_1106_1.INJECT1_1 = "NO";
    LUT4 shift_right_31_i68_3_lut (.A(d10[67]), .B(d10[68]), .C(\CICGain[0] ), 
         .Z(n68_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i68_3_lut.init = 16'hcaca;
    CCU2D add_1107_37 (.A0(d9[71]), .B0(d_d9[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11529), 
          .S0(n6010[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1107_37.INIT0 = 16'h5999;
    defparam add_1107_37.INIT1 = 16'h0000;
    defparam add_1107_37.INJECT1_0 = "NO";
    defparam add_1107_37.INJECT1_1 = "NO";
    CCU2D add_1107_35 (.A0(d9[69]), .B0(d_d9[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[70]), .B1(d_d9[70]), .C1(GND_net), .D1(GND_net), .CIN(n11528), 
          .COUT(n11529), .S0(n6010[33]), .S1(n6010[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1107_35.INIT0 = 16'h5999;
    defparam add_1107_35.INIT1 = 16'h5999;
    defparam add_1107_35.INJECT1_0 = "NO";
    defparam add_1107_35.INJECT1_1 = "NO";
    CCU2D add_1107_33 (.A0(d9[67]), .B0(d_d9[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[68]), .B1(d_d9[68]), .C1(GND_net), .D1(GND_net), .CIN(n11527), 
          .COUT(n11528), .S0(n6010[31]), .S1(n6010[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1107_33.INIT0 = 16'h5999;
    defparam add_1107_33.INIT1 = 16'h5999;
    defparam add_1107_33.INJECT1_0 = "NO";
    defparam add_1107_33.INJECT1_1 = "NO";
    CCU2D add_1107_31 (.A0(d9[65]), .B0(d_d9[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[66]), .B1(d_d9[66]), .C1(GND_net), .D1(GND_net), .CIN(n11526), 
          .COUT(n11527), .S0(n6010[29]), .S1(n6010[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1107_31.INIT0 = 16'h5999;
    defparam add_1107_31.INIT1 = 16'h5999;
    defparam add_1107_31.INJECT1_0 = "NO";
    defparam add_1107_31.INJECT1_1 = "NO";
    CCU2D add_1107_29 (.A0(d9[63]), .B0(d_d9[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[64]), .B1(d_d9[64]), .C1(GND_net), .D1(GND_net), .CIN(n11525), 
          .COUT(n11526), .S0(n6010[27]), .S1(n6010[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1107_29.INIT0 = 16'h5999;
    defparam add_1107_29.INIT1 = 16'h5999;
    defparam add_1107_29.INJECT1_0 = "NO";
    defparam add_1107_29.INJECT1_1 = "NO";
    CCU2D add_1107_27 (.A0(d9[61]), .B0(d_d9[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[62]), .B1(d_d9[62]), .C1(GND_net), .D1(GND_net), .CIN(n11524), 
          .COUT(n11525), .S0(n6010[25]), .S1(n6010[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1107_27.INIT0 = 16'h5999;
    defparam add_1107_27.INIT1 = 16'h5999;
    defparam add_1107_27.INJECT1_0 = "NO";
    defparam add_1107_27.INJECT1_1 = "NO";
    CCU2D add_1107_25 (.A0(d9[59]), .B0(d_d9[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[60]), .B1(d_d9[60]), .C1(GND_net), .D1(GND_net), .CIN(n11523), 
          .COUT(n11524), .S0(n6010[23]), .S1(n6010[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1107_25.INIT0 = 16'h5999;
    defparam add_1107_25.INIT1 = 16'h5999;
    defparam add_1107_25.INJECT1_0 = "NO";
    defparam add_1107_25.INJECT1_1 = "NO";
    CCU2D add_1107_23 (.A0(d9[57]), .B0(d_d9[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[58]), .B1(d_d9[58]), .C1(GND_net), .D1(GND_net), .CIN(n11522), 
          .COUT(n11523), .S0(n6010[21]), .S1(n6010[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1107_23.INIT0 = 16'h5999;
    defparam add_1107_23.INIT1 = 16'h5999;
    defparam add_1107_23.INJECT1_0 = "NO";
    defparam add_1107_23.INJECT1_1 = "NO";
    CCU2D add_1107_21 (.A0(d9[55]), .B0(d_d9[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[56]), .B1(d_d9[56]), .C1(GND_net), .D1(GND_net), .CIN(n11521), 
          .COUT(n11522));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1107_21.INIT0 = 16'h5999;
    defparam add_1107_21.INIT1 = 16'h5999;
    defparam add_1107_21.INJECT1_0 = "NO";
    defparam add_1107_21.INJECT1_1 = "NO";
    CCU2D add_1107_19 (.A0(d9[53]), .B0(d_d9[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[54]), .B1(d_d9[54]), .C1(GND_net), .D1(GND_net), .CIN(n11520), 
          .COUT(n11521));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1107_19.INIT0 = 16'h5999;
    defparam add_1107_19.INIT1 = 16'h5999;
    defparam add_1107_19.INJECT1_0 = "NO";
    defparam add_1107_19.INJECT1_1 = "NO";
    CCU2D add_1106_21 (.A0(d9[55]), .B0(d_d9[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[56]), .B1(d_d9[56]), .C1(GND_net), .D1(GND_net), .CIN(n11539), 
          .COUT(n11540));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1106_21.INIT0 = 16'h5999;
    defparam add_1106_21.INIT1 = 16'h5999;
    defparam add_1106_21.INJECT1_0 = "NO";
    defparam add_1106_21.INJECT1_1 = "NO";
    LUT4 shift_right_31_i205_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65_c), .D(n133), .Z(d_out_11__N_1819[4])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i205_3_lut_4_lut.init = 16'hfe10;
    LUT4 i10_4_lut (.A(count[8]), .B(count[9]), .C(count[1]), .D(count[7]), 
         .Z(n24)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i10_4_lut.init = 16'h8000;
    CCU2D add_1107_17 (.A0(d9[51]), .B0(d_d9[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[52]), .B1(d_d9[52]), .C1(GND_net), .D1(GND_net), .CIN(n11519), 
          .COUT(n11520));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1107_17.INIT0 = 16'h5999;
    defparam add_1107_17.INIT1 = 16'h5999;
    defparam add_1107_17.INJECT1_0 = "NO";
    defparam add_1107_17.INJECT1_1 = "NO";
    CCU2D add_1107_15 (.A0(d9[49]), .B0(d_d9[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[50]), .B1(d_d9[50]), .C1(GND_net), .D1(GND_net), .CIN(n11518), 
          .COUT(n11519));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1107_15.INIT0 = 16'h5999;
    defparam add_1107_15.INIT1 = 16'h5999;
    defparam add_1107_15.INJECT1_0 = "NO";
    defparam add_1107_15.INJECT1_1 = "NO";
    LUT4 shift_right_31_i206_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66_c), .D(n134), .Z(d_out_11__N_1819[5])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i206_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_1107_13 (.A0(d9[47]), .B0(d_d9[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[48]), .B1(d_d9[48]), .C1(GND_net), .D1(GND_net), .CIN(n11517), 
          .COUT(n11518));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1107_13.INIT0 = 16'h5999;
    defparam add_1107_13.INIT1 = 16'h5999;
    defparam add_1107_13.INJECT1_0 = "NO";
    defparam add_1107_13.INJECT1_1 = "NO";
    LUT4 shift_right_31_i207_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n13176), .D(n135), .Z(d_out_11__N_1819[6])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i207_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_1101_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d8[36]), .B1(d_d8[36]), .C1(GND_net), .D1(GND_net), .COUT(n11570), 
          .S1(n5820[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1101_1.INIT0 = 16'hF000;
    defparam add_1101_1.INIT1 = 16'h5999;
    defparam add_1101_1.INJECT1_0 = "NO";
    defparam add_1101_1.INJECT1_1 = "NO";
    CCU2D add_1107_11 (.A0(d9[45]), .B0(d_d9[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[46]), .B1(d_d9[46]), .C1(GND_net), .D1(GND_net), .CIN(n11516), 
          .COUT(n11517));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1107_11.INIT0 = 16'h5999;
    defparam add_1107_11.INIT1 = 16'h5999;
    defparam add_1107_11.INJECT1_0 = "NO";
    defparam add_1107_11.INJECT1_1 = "NO";
    LUT4 shift_right_31_i208_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n68_c), .D(n136), .Z(d_out_11__N_1819[7])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i208_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i141_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n137), .D(d10[68]), .Z(d_out_11__N_1819[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i141_3_lut_4_lut.init = 16'hf1e0;
    CCU2D add_1102_37 (.A0(d_d8[70]), .B0(n5819), .C0(n5820[34]), .D0(d8[70]), 
          .A1(d_d8[71]), .B1(n5819), .C1(n5820[35]), .D1(d8[71]), .CIN(n11568), 
          .S0(d9_71__N_1675[70]), .S1(d9_71__N_1675[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1102_37.INIT0 = 16'hb874;
    defparam add_1102_37.INIT1 = 16'hb874;
    defparam add_1102_37.INJECT1_0 = "NO";
    defparam add_1102_37.INJECT1_1 = "NO";
    CCU2D add_1107_9 (.A0(d9[43]), .B0(d_d9[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[44]), .B1(d_d9[44]), .C1(GND_net), .D1(GND_net), .CIN(n11515), 
          .COUT(n11516));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1107_9.INIT0 = 16'h5999;
    defparam add_1107_9.INIT1 = 16'h5999;
    defparam add_1107_9.INJECT1_0 = "NO";
    defparam add_1107_9.INJECT1_1 = "NO";
    LUT4 i7_2_lut (.A(count[9]), .B(count[7]), .Z(n21)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i2_2_lut_adj_25 (.A(count[0]), .B(count[5]), .Z(n16_adj_2489)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_25.init = 16'heeee;
    FD1P3AX d_d_tmp_i0_i29 (.D(d_tmp[29]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i29.GSR = "ENABLED";
    LUT4 shift_right_31_i210_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n70_c), .D(n138), .Z(d_out_11__N_1819[9])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i210_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_1102_35 (.A0(d_d8[68]), .B0(n5819), .C0(n5820[32]), .D0(d8[68]), 
          .A1(d_d8[69]), .B1(n5819), .C1(n5820[33]), .D1(d8[69]), .CIN(n11567), 
          .COUT(n11568), .S0(d9_71__N_1675[68]), .S1(d9_71__N_1675[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1102_35.INIT0 = 16'hb874;
    defparam add_1102_35.INIT1 = 16'hb874;
    defparam add_1102_35.INJECT1_0 = "NO";
    defparam add_1102_35.INJECT1_1 = "NO";
    CCU2D add_1102_33 (.A0(d_d8[66]), .B0(n5819), .C0(n5820[30]), .D0(d8[66]), 
          .A1(d_d8[67]), .B1(n5819), .C1(n5820[31]), .D1(d8[67]), .CIN(n11566), 
          .COUT(n11567), .S0(d9_71__N_1675[66]), .S1(d9_71__N_1675[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1102_33.INIT0 = 16'hb874;
    defparam add_1102_33.INIT1 = 16'hb874;
    defparam add_1102_33.INJECT1_0 = "NO";
    defparam add_1102_33.INJECT1_1 = "NO";
    CCU2D add_1102_31 (.A0(d_d8[64]), .B0(n5819), .C0(n5820[28]), .D0(d8[64]), 
          .A1(d_d8[65]), .B1(n5819), .C1(n5820[29]), .D1(d8[65]), .CIN(n11565), 
          .COUT(n11566), .S0(d9_71__N_1675[64]), .S1(d9_71__N_1675[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1102_31.INIT0 = 16'hb874;
    defparam add_1102_31.INIT1 = 16'hb874;
    defparam add_1102_31.INJECT1_0 = "NO";
    defparam add_1102_31.INJECT1_1 = "NO";
    LUT4 shift_right_31_i70_3_lut (.A(d10[69]), .B(d10[70]), .C(\CICGain[0] ), 
         .Z(n70_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i70_3_lut.init = 16'hcaca;
    CCU2D add_1107_7 (.A0(d9[41]), .B0(d_d9[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[42]), .B1(d_d9[42]), .C1(GND_net), .D1(GND_net), .CIN(n11514), 
          .COUT(n11515));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1107_7.INIT0 = 16'h5999;
    defparam add_1107_7.INIT1 = 16'h5999;
    defparam add_1107_7.INJECT1_0 = "NO";
    defparam add_1107_7.INJECT1_1 = "NO";
    LUT4 shift_right_31_i212_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(d10[71]), .D(n140), .Z(d_out_11__N_1819[11])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i212_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i203_3_lut_4_lut_adj_26 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63), .D(n131_adj_2491), .Z(\d_out_11__N_1819[2] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i203_3_lut_4_lut_adj_26.init = 16'hfe10;
    LUT4 shift_right_31_i204_3_lut_4_lut_adj_27 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64), .D(n132), .Z(\d_out_11__N_1819[3] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i204_3_lut_4_lut_adj_27.init = 16'hfe10;
    CCU2D add_1102_29 (.A0(d_d8[62]), .B0(n5819), .C0(n5820[26]), .D0(d8[62]), 
          .A1(d_d8[63]), .B1(n5819), .C1(n5820[27]), .D1(d8[63]), .CIN(n11564), 
          .COUT(n11565), .S0(d9_71__N_1675[62]), .S1(d9_71__N_1675[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1102_29.INIT0 = 16'hb874;
    defparam add_1102_29.INIT1 = 16'hb874;
    defparam add_1102_29.INJECT1_0 = "NO";
    defparam add_1102_29.INJECT1_1 = "NO";
    CCU2D add_1102_27 (.A0(d_d8[60]), .B0(n5819), .C0(n5820[24]), .D0(d8[60]), 
          .A1(d_d8[61]), .B1(n5819), .C1(n5820[25]), .D1(d8[61]), .CIN(n11563), 
          .COUT(n11564), .S0(d9_71__N_1675[60]), .S1(d9_71__N_1675[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1102_27.INIT0 = 16'hb874;
    defparam add_1102_27.INIT1 = 16'hb874;
    defparam add_1102_27.INJECT1_0 = "NO";
    defparam add_1102_27.INJECT1_1 = "NO";
    CCU2D add_1102_25 (.A0(d_d8[58]), .B0(n5819), .C0(n5820[22]), .D0(d8[58]), 
          .A1(d_d8[59]), .B1(n5819), .C1(n5820[23]), .D1(d8[59]), .CIN(n11562), 
          .COUT(n11563), .S0(d9_71__N_1675[58]), .S1(d9_71__N_1675[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1102_25.INIT0 = 16'hb874;
    defparam add_1102_25.INIT1 = 16'hb874;
    defparam add_1102_25.INJECT1_0 = "NO";
    defparam add_1102_25.INJECT1_1 = "NO";
    CCU2D add_1102_23 (.A0(d_d8[56]), .B0(n5819), .C0(n5820[20]), .D0(d8[56]), 
          .A1(d_d8[57]), .B1(n5819), .C1(n5820[21]), .D1(d8[57]), .CIN(n11561), 
          .COUT(n11562), .S0(d9_71__N_1675[56]), .S1(d9_71__N_1675[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1102_23.INIT0 = 16'hb874;
    defparam add_1102_23.INIT1 = 16'hb874;
    defparam add_1102_23.INJECT1_0 = "NO";
    defparam add_1102_23.INJECT1_1 = "NO";
    CCU2D add_1102_21 (.A0(d_d8[54]), .B0(n5819), .C0(n5820[18]), .D0(d8[54]), 
          .A1(d_d8[55]), .B1(n5819), .C1(n5820[19]), .D1(d8[55]), .CIN(n11560), 
          .COUT(n11561), .S0(d9_71__N_1675[54]), .S1(d9_71__N_1675[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1102_21.INIT0 = 16'hb874;
    defparam add_1102_21.INIT1 = 16'hb874;
    defparam add_1102_21.INJECT1_0 = "NO";
    defparam add_1102_21.INJECT1_1 = "NO";
    CCU2D add_1102_19 (.A0(d_d8[52]), .B0(n5819), .C0(n5820[16]), .D0(d8[52]), 
          .A1(d_d8[53]), .B1(n5819), .C1(n5820[17]), .D1(d8[53]), .CIN(n11559), 
          .COUT(n11560), .S0(d9_71__N_1675[52]), .S1(d9_71__N_1675[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1102_19.INIT0 = 16'hb874;
    defparam add_1102_19.INIT1 = 16'hb874;
    defparam add_1102_19.INJECT1_0 = "NO";
    defparam add_1102_19.INJECT1_1 = "NO";
    CCU2D add_1102_17 (.A0(d_d8[50]), .B0(n5819), .C0(n5820[14]), .D0(d8[50]), 
          .A1(d_d8[51]), .B1(n5819), .C1(n5820[15]), .D1(d8[51]), .CIN(n11558), 
          .COUT(n11559), .S0(d9_71__N_1675[50]), .S1(d9_71__N_1675[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1102_17.INIT0 = 16'hb874;
    defparam add_1102_17.INIT1 = 16'hb874;
    defparam add_1102_17.INJECT1_0 = "NO";
    defparam add_1102_17.INJECT1_1 = "NO";
    CCU2D add_1102_15 (.A0(d_d8[48]), .B0(n5819), .C0(n5820[12]), .D0(d8[48]), 
          .A1(d_d8[49]), .B1(n5819), .C1(n5820[13]), .D1(d8[49]), .CIN(n11557), 
          .COUT(n11558), .S0(d9_71__N_1675[48]), .S1(d9_71__N_1675[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1102_15.INIT0 = 16'hb874;
    defparam add_1102_15.INIT1 = 16'hb874;
    defparam add_1102_15.INJECT1_0 = "NO";
    defparam add_1102_15.INJECT1_1 = "NO";
    CCU2D add_1107_5 (.A0(d9[39]), .B0(d_d9[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[40]), .B1(d_d9[40]), .C1(GND_net), .D1(GND_net), .CIN(n11513), 
          .COUT(n11514));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1107_5.INIT0 = 16'h5999;
    defparam add_1107_5.INIT1 = 16'h5999;
    defparam add_1107_5.INJECT1_0 = "NO";
    defparam add_1107_5.INJECT1_1 = "NO";
    CCU2D add_1102_13 (.A0(d_d8[46]), .B0(n5819), .C0(n5820[10]), .D0(d8[46]), 
          .A1(d_d8[47]), .B1(n5819), .C1(n5820[11]), .D1(d8[47]), .CIN(n11556), 
          .COUT(n11557), .S0(d9_71__N_1675[46]), .S1(d9_71__N_1675[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1102_13.INIT0 = 16'hb874;
    defparam add_1102_13.INIT1 = 16'hb874;
    defparam add_1102_13.INJECT1_0 = "NO";
    defparam add_1102_13.INJECT1_1 = "NO";
    CCU2D add_1107_3 (.A0(d9[37]), .B0(d_d9[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[38]), .B1(d_d9[38]), .C1(GND_net), .D1(GND_net), .CIN(n11512), 
          .COUT(n11513));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1107_3.INIT0 = 16'h5999;
    defparam add_1107_3.INIT1 = 16'h5999;
    defparam add_1107_3.INJECT1_0 = "NO";
    defparam add_1107_3.INJECT1_1 = "NO";
    CCU2D add_1102_11 (.A0(d_d8[44]), .B0(n5819), .C0(n5820[8]), .D0(d8[44]), 
          .A1(d_d8[45]), .B1(n5819), .C1(n5820[9]), .D1(d8[45]), .CIN(n11555), 
          .COUT(n11556), .S0(d9_71__N_1675[44]), .S1(d9_71__N_1675[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1102_11.INIT0 = 16'hb874;
    defparam add_1102_11.INIT1 = 16'hb874;
    defparam add_1102_11.INJECT1_0 = "NO";
    defparam add_1102_11.INJECT1_1 = "NO";
    CCU2D add_1102_9 (.A0(d_d8[42]), .B0(n5819), .C0(n5820[6]), .D0(d8[42]), 
          .A1(d_d8[43]), .B1(n5819), .C1(n5820[7]), .D1(d8[43]), .CIN(n11554), 
          .COUT(n11555), .S0(d9_71__N_1675[42]), .S1(d9_71__N_1675[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1102_9.INIT0 = 16'hb874;
    defparam add_1102_9.INIT1 = 16'hb874;
    defparam add_1102_9.INJECT1_0 = "NO";
    defparam add_1102_9.INJECT1_1 = "NO";
    CCU2D add_1102_7 (.A0(d_d8[40]), .B0(n5819), .C0(n5820[4]), .D0(d8[40]), 
          .A1(d_d8[41]), .B1(n5819), .C1(n5820[5]), .D1(d8[41]), .CIN(n11553), 
          .COUT(n11554), .S0(d9_71__N_1675[40]), .S1(d9_71__N_1675[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1102_7.INIT0 = 16'hb874;
    defparam add_1102_7.INIT1 = 16'hb874;
    defparam add_1102_7.INJECT1_0 = "NO";
    defparam add_1102_7.INJECT1_1 = "NO";
    CCU2D add_1102_5 (.A0(d_d8[38]), .B0(n5819), .C0(n5820[2]), .D0(d8[38]), 
          .A1(d_d8[39]), .B1(n5819), .C1(n5820[3]), .D1(d8[39]), .CIN(n11552), 
          .COUT(n11553), .S0(d9_71__N_1675[38]), .S1(d9_71__N_1675[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1102_5.INIT0 = 16'hb874;
    defparam add_1102_5.INIT1 = 16'hb874;
    defparam add_1102_5.INJECT1_0 = "NO";
    defparam add_1102_5.INJECT1_1 = "NO";
    CCU2D add_1102_3 (.A0(d_d8[36]), .B0(n5819), .C0(n5820[0]), .D0(d8[36]), 
          .A1(d_d8[37]), .B1(n5819), .C1(n5820[1]), .D1(d8[37]), .CIN(n11551), 
          .COUT(n11552), .S0(d9_71__N_1675[36]), .S1(d9_71__N_1675[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1102_3.INIT0 = 16'hb874;
    defparam add_1102_3.INIT1 = 16'hb874;
    defparam add_1102_3.INJECT1_0 = "NO";
    defparam add_1102_3.INJECT1_1 = "NO";
    CCU2D add_1102_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5819), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11551));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1102_1.INIT0 = 16'hF000;
    defparam add_1102_1.INIT1 = 16'h0555;
    defparam add_1102_1.INJECT1_0 = "NO";
    defparam add_1102_1.INJECT1_1 = "NO";
    CCU2D add_1106_37 (.A0(d9[71]), .B0(d_d9[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11547), 
          .S0(n5972[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1106_37.INIT0 = 16'h5999;
    defparam add_1106_37.INIT1 = 16'h0000;
    defparam add_1106_37.INJECT1_0 = "NO";
    defparam add_1106_37.INJECT1_1 = "NO";
    CCU2D add_1106_35 (.A0(d9[69]), .B0(d_d9[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[70]), .B1(d_d9[70]), .C1(GND_net), .D1(GND_net), .CIN(n11546), 
          .COUT(n11547), .S0(n5972[33]), .S1(n5972[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1106_35.INIT0 = 16'h5999;
    defparam add_1106_35.INIT1 = 16'h5999;
    defparam add_1106_35.INJECT1_0 = "NO";
    defparam add_1106_35.INJECT1_1 = "NO";
    CCU2D add_1106_33 (.A0(d9[67]), .B0(d_d9[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[68]), .B1(d_d9[68]), .C1(GND_net), .D1(GND_net), .CIN(n11545), 
          .COUT(n11546), .S0(n5972[31]), .S1(n5972[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1106_33.INIT0 = 16'h5999;
    defparam add_1106_33.INIT1 = 16'h5999;
    defparam add_1106_33.INJECT1_0 = "NO";
    defparam add_1106_33.INJECT1_1 = "NO";
    CCU2D add_1106_31 (.A0(d9[65]), .B0(d_d9[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[66]), .B1(d_d9[66]), .C1(GND_net), .D1(GND_net), .CIN(n11544), 
          .COUT(n11545), .S0(n5972[29]), .S1(n5972[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1106_31.INIT0 = 16'h5999;
    defparam add_1106_31.INIT1 = 16'h5999;
    defparam add_1106_31.INJECT1_0 = "NO";
    defparam add_1106_31.INJECT1_1 = "NO";
    CCU2D add_1107_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d9[36]), .B1(d_d9[36]), .C1(GND_net), .D1(GND_net), .COUT(n11512));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1107_1.INIT0 = 16'h0000;
    defparam add_1107_1.INIT1 = 16'h5999;
    defparam add_1107_1.INJECT1_0 = "NO";
    defparam add_1107_1.INJECT1_1 = "NO";
    LUT4 i13_4_lut (.A(n21_adj_2495), .B(n26), .C(n15), .D(n16), .Z(d_clk_tmp_N_1831)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i13_4_lut.init = 16'h8000;
    FD1P3AX d_d_tmp_i0_i30 (.D(d_tmp[30]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i31 (.D(d_tmp[31]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i31.GSR = "ENABLED";
    CCU2D add_1056_26 (.A0(d1[60]), .B0(d2[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[61]), .B1(d2[61]), .C1(GND_net), .D1(GND_net), .CIN(n11950), 
          .COUT(n11951), .S0(n4452[24]), .S1(n4452[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1056_26.INIT0 = 16'h5666;
    defparam add_1056_26.INIT1 = 16'h5666;
    defparam add_1056_26.INJECT1_0 = "NO";
    defparam add_1056_26.INJECT1_1 = "NO";
    LUT4 shift_right_31_i205_3_lut_4_lut_adj_28 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65), .D(n133_adj_2497), .Z(\d_out_11__N_1819[4] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i205_3_lut_4_lut_adj_28.init = 16'hfe10;
    LUT4 shift_right_31_i206_3_lut_4_lut_adj_29 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66), .D(n134_adj_2500), .Z(\d_out_11__N_1819[5] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i206_3_lut_4_lut_adj_29.init = 16'hfe10;
    LUT4 shift_right_31_i207_3_lut_4_lut_adj_30 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n67), .D(n135_adj_2502), .Z(\d_out_11__N_1819[6] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i207_3_lut_4_lut_adj_30.init = 16'hfe10;
    LUT4 shift_right_31_i208_3_lut_4_lut_adj_31 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n68), .D(n136_adj_2505), .Z(\d_out_11__N_1819[7] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i208_3_lut_4_lut_adj_31.init = 16'hfe10;
    LUT4 shift_right_31_i141_3_lut_4_lut_adj_32 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n137_adj_2507), .D(\d10[68] ), .Z(\d_out_11__N_1819[8] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i141_3_lut_4_lut_adj_32.init = 16'hf1e0;
    LUT4 i12_4_lut (.A(n17), .B(n24), .C(count[6]), .D(count[11]), .Z(n26)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i12_4_lut.init = 16'h8000;
    FD1P3AX d_tmp_i0_i14 (.D(d5[14]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i18 (.D(d_tmp[18]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i17 (.D(d_tmp[17]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i16 (.D(d_tmp[16]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i16.GSR = "ENABLED";
    CCU2D add_1106_19 (.A0(d9[53]), .B0(d_d9[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[54]), .B1(d_d9[54]), .C1(GND_net), .D1(GND_net), .CIN(n11538), 
          .COUT(n11539));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1106_19.INIT0 = 16'h5999;
    defparam add_1106_19.INIT1 = 16'h5999;
    defparam add_1106_19.INJECT1_0 = "NO";
    defparam add_1106_19.INJECT1_1 = "NO";
    FD1P3AX d_d_tmp_i0_i15 (.D(d_tmp[15]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i15.GSR = "ENABLED";
    LUT4 shift_right_31_i210_3_lut_4_lut_adj_33 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n70), .D(n138_adj_2511), .Z(\d_out_11__N_1819[9] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i210_3_lut_4_lut_adj_33.init = 16'hfe10;
    FD1P3AX d_d_tmp_i0_i14 (.D(d_tmp[14]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i13 (.D(d_tmp[13]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i12 (.D(d_tmp[12]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i11 (.D(d_tmp[11]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i10 (.D(d_tmp[10]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i9 (.D(d_tmp[9]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i8 (.D(d_tmp[8]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i7 (.D(d_tmp[7]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i6 (.D(d_tmp[6]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i5 (.D(d_tmp[5]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i4 (.D(d_tmp[4]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i4.GSR = "ENABLED";
    CCU2D add_1106_17 (.A0(d9[51]), .B0(d_d9[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[52]), .B1(d_d9[52]), .C1(GND_net), .D1(GND_net), .CIN(n11537), 
          .COUT(n11538));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1106_17.INIT0 = 16'h5999;
    defparam add_1106_17.INIT1 = 16'h5999;
    defparam add_1106_17.INJECT1_0 = "NO";
    defparam add_1106_17.INJECT1_1 = "NO";
    FD1S3IX count__i1 (.D(n375[1]), .CK(osc_clk), .CD(n8425), .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i1.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i3 (.D(d_tmp[3]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i2 (.D(d_tmp[2]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i1 (.D(d_tmp[1]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d_d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i71 (.D(d5[71]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i70 (.D(d5[70]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i69 (.D(d5[69]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i68 (.D(d5[68]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i67 (.D(d5[67]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i66 (.D(d5[66]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i65 (.D(d5[65]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i64 (.D(d5[64]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i63 (.D(d5[63]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i62 (.D(d5[62]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i61 (.D(d5[61]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i60 (.D(d5[60]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i59 (.D(d5[59]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i58 (.D(d5[58]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i57 (.D(d5[57]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i56 (.D(d5[56]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i55 (.D(d5[55]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i54 (.D(d5[54]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i53 (.D(d5[53]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i52 (.D(d5[52]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i51 (.D(d5[51]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i50 (.D(d5[50]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i49 (.D(d5[49]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i48 (.D(d5[48]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i47 (.D(d5[47]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i46 (.D(d5[46]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i45 (.D(d5[45]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i44 (.D(d5[44]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i43 (.D(d5[43]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i42 (.D(d5[42]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i41 (.D(d5[41]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i40 (.D(d5[40]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i39 (.D(d5[39]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i38 (.D(d5[38]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i37 (.D(d5[37]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i36 (.D(d5[36]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i35 (.D(d5[35]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i34 (.D(d5[34]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i33 (.D(d5[33]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i32 (.D(d5[32]), .SP(osc_clk_enable_141), .CK(osc_clk), 
            .Q(d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i31 (.D(d5[31]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i30 (.D(d5[30]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i29 (.D(d5[29]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i28 (.D(d5[28]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i27 (.D(d5[27]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i26 (.D(d5[26]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i25 (.D(d5[25]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i24 (.D(d5[24]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i23 (.D(d5[23]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i22 (.D(d5[22]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i21 (.D(d5[21]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i20 (.D(d5[20]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i19 (.D(d5[19]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i18 (.D(d5[18]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i17 (.D(d5[17]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i13 (.D(d5[13]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i12 (.D(d5[12]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i12.GSR = "ENABLED";
    LUT4 shift_right_31_i212_3_lut_4_lut_adj_34 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(\d10[71] ), .D(n140_adj_2514), .Z(\d_out_11__N_1819[11] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i212_3_lut_4_lut_adj_34.init = 16'hfe10;
    FD1P3AX d_tmp_i0_i16 (.D(d5[16]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i11 (.D(d5[11]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i11.GSR = "ENABLED";
    LUT4 i4652_2_lut (.A(d2[36]), .B(d3[36]), .Z(n4604[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4652_2_lut.init = 16'h6666;
    FD1P3AX d_tmp_i0_i10 (.D(d5[10]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i10.GSR = "ENABLED";
    LUT4 i4649_2_lut (.A(d3[36]), .B(d4[36]), .Z(n4756[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4649_2_lut.init = 16'h6666;
    FD1S3AX v_comb_66_rep_113 (.D(osc_clk_enable_141), .CK(osc_clk), .Q(osc_clk_enable_660)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_113.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i9 (.D(d5[9]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i8 (.D(d5[8]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i7 (.D(d5[7]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i6 (.D(d5[6]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i5 (.D(d5[5]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i5.GSR = "ENABLED";
    LUT4 i73_2_lut_rep_95 (.A(count[13]), .B(count[15]), .Z(n13069)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i73_2_lut_rep_95.init = 16'heeee;
    FD1S3AX d2_i1 (.D(d2_71__N_490[1]), .CK(osc_clk), .Q(d2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i1.GSR = "ENABLED";
    CCU2D add_1056_24 (.A0(d1[58]), .B0(d2[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[59]), .B1(d2[59]), .C1(GND_net), .D1(GND_net), .CIN(n11949), 
          .COUT(n11950), .S0(n4452[22]), .S1(n4452[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1056_24.INIT0 = 16'h5666;
    defparam add_1056_24.INIT1 = 16'h5666;
    defparam add_1056_24.INJECT1_0 = "NO";
    defparam add_1056_24.INJECT1_1 = "NO";
    CCU2D add_1056_22 (.A0(d1[56]), .B0(d2[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[57]), .B1(d2[57]), .C1(GND_net), .D1(GND_net), .CIN(n11948), 
          .COUT(n11949), .S0(n4452[20]), .S1(n4452[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1056_22.INIT0 = 16'h5666;
    defparam add_1056_22.INIT1 = 16'h5666;
    defparam add_1056_22.INJECT1_0 = "NO";
    defparam add_1056_22.INJECT1_1 = "NO";
    CCU2D add_1056_20 (.A0(d1[54]), .B0(d2[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[55]), .B1(d2[55]), .C1(GND_net), .D1(GND_net), .CIN(n11947), 
          .COUT(n11948), .S0(n4452[18]), .S1(n4452[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1056_20.INIT0 = 16'h5666;
    defparam add_1056_20.INIT1 = 16'h5666;
    defparam add_1056_20.INJECT1_0 = "NO";
    defparam add_1056_20.INJECT1_1 = "NO";
    CCU2D add_1056_18 (.A0(d1[52]), .B0(d2[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[53]), .B1(d2[53]), .C1(GND_net), .D1(GND_net), .CIN(n11946), 
          .COUT(n11947), .S0(n4452[16]), .S1(n4452[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1056_18.INIT0 = 16'h5666;
    defparam add_1056_18.INIT1 = 16'h5666;
    defparam add_1056_18.INJECT1_0 = "NO";
    defparam add_1056_18.INJECT1_1 = "NO";
    CCU2D add_1056_16 (.A0(d1[50]), .B0(d2[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[51]), .B1(d2[51]), .C1(GND_net), .D1(GND_net), .CIN(n11945), 
          .COUT(n11946), .S0(n4452[14]), .S1(n4452[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1056_16.INIT0 = 16'h5666;
    defparam add_1056_16.INIT1 = 16'h5666;
    defparam add_1056_16.INJECT1_0 = "NO";
    defparam add_1056_16.INJECT1_1 = "NO";
    CCU2D add_1056_14 (.A0(d1[48]), .B0(d2[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[49]), .B1(d2[49]), .C1(GND_net), .D1(GND_net), .CIN(n11944), 
          .COUT(n11945), .S0(n4452[12]), .S1(n4452[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1056_14.INIT0 = 16'h5666;
    defparam add_1056_14.INIT1 = 16'h5666;
    defparam add_1056_14.INJECT1_0 = "NO";
    defparam add_1056_14.INJECT1_1 = "NO";
    CCU2D add_1056_12 (.A0(d1[46]), .B0(d2[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[47]), .B1(d2[47]), .C1(GND_net), .D1(GND_net), .CIN(n11943), 
          .COUT(n11944), .S0(n4452[10]), .S1(n4452[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1056_12.INIT0 = 16'h5666;
    defparam add_1056_12.INIT1 = 16'h5666;
    defparam add_1056_12.INJECT1_0 = "NO";
    defparam add_1056_12.INJECT1_1 = "NO";
    CCU2D add_1056_10 (.A0(d1[44]), .B0(d2[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[45]), .B1(d2[45]), .C1(GND_net), .D1(GND_net), .CIN(n11942), 
          .COUT(n11943), .S0(n4452[8]), .S1(n4452[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1056_10.INIT0 = 16'h5666;
    defparam add_1056_10.INIT1 = 16'h5666;
    defparam add_1056_10.INJECT1_0 = "NO";
    defparam add_1056_10.INJECT1_1 = "NO";
    CCU2D add_1056_8 (.A0(d1[42]), .B0(d2[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[43]), .B1(d2[43]), .C1(GND_net), .D1(GND_net), .CIN(n11941), 
          .COUT(n11942), .S0(n4452[6]), .S1(n4452[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1056_8.INIT0 = 16'h5666;
    defparam add_1056_8.INIT1 = 16'h5666;
    defparam add_1056_8.INJECT1_0 = "NO";
    defparam add_1056_8.INJECT1_1 = "NO";
    CCU2D add_1056_6 (.A0(d1[40]), .B0(d2[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[41]), .B1(d2[41]), .C1(GND_net), .D1(GND_net), .CIN(n11940), 
          .COUT(n11941), .S0(n4452[4]), .S1(n4452[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1056_6.INIT0 = 16'h5666;
    defparam add_1056_6.INIT1 = 16'h5666;
    defparam add_1056_6.INJECT1_0 = "NO";
    defparam add_1056_6.INJECT1_1 = "NO";
    CCU2D add_1056_4 (.A0(d1[38]), .B0(d2[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[39]), .B1(d2[39]), .C1(GND_net), .D1(GND_net), .CIN(n11939), 
          .COUT(n11940), .S0(n4452[2]), .S1(n4452[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1056_4.INIT0 = 16'h5666;
    defparam add_1056_4.INIT1 = 16'h5666;
    defparam add_1056_4.INJECT1_0 = "NO";
    defparam add_1056_4.INJECT1_1 = "NO";
    CCU2D add_1056_2 (.A0(d1[36]), .B0(d2[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[37]), .B1(d2[37]), .C1(GND_net), .D1(GND_net), .COUT(n11939), 
          .S1(n4452[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1056_2.INIT0 = 16'h7000;
    defparam add_1056_2.INIT1 = 16'h5666;
    defparam add_1056_2.INJECT1_0 = "NO";
    defparam add_1056_2.INJECT1_1 = "NO";
    FD1S3AX d2_i2 (.D(d2_71__N_490[2]), .CK(osc_clk), .Q(d2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i2.GSR = "ENABLED";
    FD1S3AX d2_i3 (.D(d2_71__N_490[3]), .CK(osc_clk), .Q(d2[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i3.GSR = "ENABLED";
    FD1S3AX d2_i4 (.D(d2_71__N_490[4]), .CK(osc_clk), .Q(d2[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i4.GSR = "ENABLED";
    FD1S3AX d2_i5 (.D(d2_71__N_490[5]), .CK(osc_clk), .Q(d2[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i5.GSR = "ENABLED";
    FD1S3AX d2_i6 (.D(d2_71__N_490[6]), .CK(osc_clk), .Q(d2[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i6.GSR = "ENABLED";
    FD1S3AX d2_i7 (.D(d2_71__N_490[7]), .CK(osc_clk), .Q(d2[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i7.GSR = "ENABLED";
    FD1S3AX d2_i8 (.D(d2_71__N_490[8]), .CK(osc_clk), .Q(d2[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i8.GSR = "ENABLED";
    FD1S3AX d2_i9 (.D(d2_71__N_490[9]), .CK(osc_clk), .Q(d2[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i9.GSR = "ENABLED";
    FD1S3AX d2_i10 (.D(d2_71__N_490[10]), .CK(osc_clk), .Q(d2[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i10.GSR = "ENABLED";
    FD1S3AX d2_i11 (.D(d2_71__N_490[11]), .CK(osc_clk), .Q(d2[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i11.GSR = "ENABLED";
    FD1S3AX d2_i12 (.D(d2_71__N_490[12]), .CK(osc_clk), .Q(d2[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i12.GSR = "ENABLED";
    FD1S3AX d2_i13 (.D(d2_71__N_490[13]), .CK(osc_clk), .Q(d2[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i13.GSR = "ENABLED";
    FD1S3AX d2_i14 (.D(d2_71__N_490[14]), .CK(osc_clk), .Q(d2[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i14.GSR = "ENABLED";
    FD1S3AX d2_i15 (.D(d2_71__N_490[15]), .CK(osc_clk), .Q(d2[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i15.GSR = "ENABLED";
    FD1S3AX d2_i16 (.D(d2_71__N_490[16]), .CK(osc_clk), .Q(d2[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i16.GSR = "ENABLED";
    FD1S3AX d2_i17 (.D(d2_71__N_490[17]), .CK(osc_clk), .Q(d2[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i17.GSR = "ENABLED";
    FD1S3AX d2_i18 (.D(d2_71__N_490[18]), .CK(osc_clk), .Q(d2[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i18.GSR = "ENABLED";
    FD1S3AX d2_i19 (.D(d2_71__N_490[19]), .CK(osc_clk), .Q(d2[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i19.GSR = "ENABLED";
    FD1S3AX d2_i20 (.D(d2_71__N_490[20]), .CK(osc_clk), .Q(d2[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i20.GSR = "ENABLED";
    FD1S3AX d2_i21 (.D(d2_71__N_490[21]), .CK(osc_clk), .Q(d2[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i21.GSR = "ENABLED";
    FD1S3AX d2_i22 (.D(d2_71__N_490[22]), .CK(osc_clk), .Q(d2[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i22.GSR = "ENABLED";
    FD1S3AX d2_i23 (.D(d2_71__N_490[23]), .CK(osc_clk), .Q(d2[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i23.GSR = "ENABLED";
    FD1S3AX d2_i24 (.D(d2_71__N_490[24]), .CK(osc_clk), .Q(d2[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i24.GSR = "ENABLED";
    FD1S3AX d2_i25 (.D(d2_71__N_490[25]), .CK(osc_clk), .Q(d2[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i25.GSR = "ENABLED";
    FD1S3AX d2_i26 (.D(d2_71__N_490[26]), .CK(osc_clk), .Q(d2[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i26.GSR = "ENABLED";
    FD1S3AX d2_i27 (.D(d2_71__N_490[27]), .CK(osc_clk), .Q(d2[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i27.GSR = "ENABLED";
    FD1S3AX d2_i28 (.D(d2_71__N_490[28]), .CK(osc_clk), .Q(d2[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i28.GSR = "ENABLED";
    FD1S3AX d2_i29 (.D(d2_71__N_490[29]), .CK(osc_clk), .Q(d2[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i29.GSR = "ENABLED";
    FD1S3AX d2_i30 (.D(d2_71__N_490[30]), .CK(osc_clk), .Q(d2[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i30.GSR = "ENABLED";
    FD1S3AX d2_i31 (.D(d2_71__N_490[31]), .CK(osc_clk), .Q(d2[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i31.GSR = "ENABLED";
    FD1S3AX d2_i32 (.D(d2_71__N_490[32]), .CK(osc_clk), .Q(d2[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i32.GSR = "ENABLED";
    FD1S3AX d2_i33 (.D(d2_71__N_490[33]), .CK(osc_clk), .Q(d2[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i33.GSR = "ENABLED";
    FD1S3AX d2_i34 (.D(d2_71__N_490[34]), .CK(osc_clk), .Q(d2[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i34.GSR = "ENABLED";
    FD1S3AX d2_i35 (.D(d2_71__N_490[35]), .CK(osc_clk), .Q(d2[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i35.GSR = "ENABLED";
    FD1S3AX d2_i36 (.D(d2_71__N_490[36]), .CK(osc_clk), .Q(d2[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i36.GSR = "ENABLED";
    FD1S3AX d2_i37 (.D(d2_71__N_490[37]), .CK(osc_clk), .Q(d2[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i37.GSR = "ENABLED";
    FD1S3AX d2_i38 (.D(d2_71__N_490[38]), .CK(osc_clk), .Q(d2[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i38.GSR = "ENABLED";
    FD1S3AX d2_i39 (.D(d2_71__N_490[39]), .CK(osc_clk), .Q(d2[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i39.GSR = "ENABLED";
    FD1S3AX d2_i40 (.D(d2_71__N_490[40]), .CK(osc_clk), .Q(d2[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i40.GSR = "ENABLED";
    FD1S3AX d2_i41 (.D(d2_71__N_490[41]), .CK(osc_clk), .Q(d2[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i41.GSR = "ENABLED";
    FD1S3AX d2_i42 (.D(d2_71__N_490[42]), .CK(osc_clk), .Q(d2[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i42.GSR = "ENABLED";
    FD1S3AX d2_i43 (.D(d2_71__N_490[43]), .CK(osc_clk), .Q(d2[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i43.GSR = "ENABLED";
    FD1S3AX d2_i44 (.D(d2_71__N_490[44]), .CK(osc_clk), .Q(d2[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i44.GSR = "ENABLED";
    FD1S3AX d2_i45 (.D(d2_71__N_490[45]), .CK(osc_clk), .Q(d2[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i45.GSR = "ENABLED";
    FD1S3AX d2_i46 (.D(d2_71__N_490[46]), .CK(osc_clk), .Q(d2[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i46.GSR = "ENABLED";
    FD1S3AX d2_i47 (.D(d2_71__N_490[47]), .CK(osc_clk), .Q(d2[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i47.GSR = "ENABLED";
    FD1S3AX d2_i48 (.D(d2_71__N_490[48]), .CK(osc_clk), .Q(d2[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i48.GSR = "ENABLED";
    FD1S3AX d2_i49 (.D(d2_71__N_490[49]), .CK(osc_clk), .Q(d2[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i49.GSR = "ENABLED";
    FD1S3AX d2_i50 (.D(d2_71__N_490[50]), .CK(osc_clk), .Q(d2[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i50.GSR = "ENABLED";
    FD1S3AX d2_i51 (.D(d2_71__N_490[51]), .CK(osc_clk), .Q(d2[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i51.GSR = "ENABLED";
    FD1S3AX d2_i52 (.D(d2_71__N_490[52]), .CK(osc_clk), .Q(d2[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i52.GSR = "ENABLED";
    FD1S3AX d2_i53 (.D(d2_71__N_490[53]), .CK(osc_clk), .Q(d2[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i53.GSR = "ENABLED";
    FD1S3AX d2_i54 (.D(d2_71__N_490[54]), .CK(osc_clk), .Q(d2[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i54.GSR = "ENABLED";
    FD1S3AX d2_i55 (.D(d2_71__N_490[55]), .CK(osc_clk), .Q(d2[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i55.GSR = "ENABLED";
    FD1S3AX d2_i56 (.D(d2_71__N_490[56]), .CK(osc_clk), .Q(d2[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i56.GSR = "ENABLED";
    FD1S3AX d2_i57 (.D(d2_71__N_490[57]), .CK(osc_clk), .Q(d2[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i57.GSR = "ENABLED";
    FD1S3AX d2_i58 (.D(d2_71__N_490[58]), .CK(osc_clk), .Q(d2[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i58.GSR = "ENABLED";
    FD1S3AX d2_i59 (.D(d2_71__N_490[59]), .CK(osc_clk), .Q(d2[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i59.GSR = "ENABLED";
    FD1S3AX d2_i60 (.D(d2_71__N_490[60]), .CK(osc_clk), .Q(d2[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i60.GSR = "ENABLED";
    FD1S3AX d2_i61 (.D(d2_71__N_490[61]), .CK(osc_clk), .Q(d2[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i61.GSR = "ENABLED";
    FD1S3AX d2_i62 (.D(d2_71__N_490[62]), .CK(osc_clk), .Q(d2[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i62.GSR = "ENABLED";
    FD1S3AX d2_i63 (.D(d2_71__N_490[63]), .CK(osc_clk), .Q(d2[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i63.GSR = "ENABLED";
    FD1S3AX d2_i64 (.D(d2_71__N_490[64]), .CK(osc_clk), .Q(d2[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i64.GSR = "ENABLED";
    FD1S3AX d2_i65 (.D(d2_71__N_490[65]), .CK(osc_clk), .Q(d2[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i65.GSR = "ENABLED";
    FD1S3AX d2_i66 (.D(d2_71__N_490[66]), .CK(osc_clk), .Q(d2[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i66.GSR = "ENABLED";
    FD1S3AX d2_i67 (.D(d2_71__N_490[67]), .CK(osc_clk), .Q(d2[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i67.GSR = "ENABLED";
    FD1S3AX d2_i68 (.D(d2_71__N_490[68]), .CK(osc_clk), .Q(d2[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i68.GSR = "ENABLED";
    FD1S3AX d2_i69 (.D(d2_71__N_490[69]), .CK(osc_clk), .Q(d2[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i69.GSR = "ENABLED";
    FD1S3AX d2_i70 (.D(d2_71__N_490[70]), .CK(osc_clk), .Q(d2[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i70.GSR = "ENABLED";
    FD1S3AX d2_i71 (.D(d2_71__N_490[71]), .CK(osc_clk), .Q(d2[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i71.GSR = "ENABLED";
    FD1S3AX d3_i1 (.D(d3_71__N_562[1]), .CK(osc_clk), .Q(d3[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i1.GSR = "ENABLED";
    FD1S3AX d3_i2 (.D(d3_71__N_562[2]), .CK(osc_clk), .Q(d3[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i2.GSR = "ENABLED";
    FD1S3AX d3_i3 (.D(d3_71__N_562[3]), .CK(osc_clk), .Q(d3[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i3.GSR = "ENABLED";
    FD1S3AX d3_i4 (.D(d3_71__N_562[4]), .CK(osc_clk), .Q(d3[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i4.GSR = "ENABLED";
    FD1S3AX d3_i5 (.D(d3_71__N_562[5]), .CK(osc_clk), .Q(d3[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i5.GSR = "ENABLED";
    FD1S3AX d3_i6 (.D(d3_71__N_562[6]), .CK(osc_clk), .Q(d3[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i6.GSR = "ENABLED";
    FD1S3AX d3_i7 (.D(d3_71__N_562[7]), .CK(osc_clk), .Q(d3[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i7.GSR = "ENABLED";
    FD1S3AX d3_i8 (.D(d3_71__N_562[8]), .CK(osc_clk), .Q(d3[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i8.GSR = "ENABLED";
    FD1S3AX d3_i9 (.D(d3_71__N_562[9]), .CK(osc_clk), .Q(d3[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i9.GSR = "ENABLED";
    FD1S3AX d3_i10 (.D(d3_71__N_562[10]), .CK(osc_clk), .Q(d3[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i10.GSR = "ENABLED";
    FD1S3AX d3_i11 (.D(d3_71__N_562[11]), .CK(osc_clk), .Q(d3[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i11.GSR = "ENABLED";
    FD1S3AX d3_i12 (.D(d3_71__N_562[12]), .CK(osc_clk), .Q(d3[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i12.GSR = "ENABLED";
    FD1S3AX d3_i13 (.D(d3_71__N_562[13]), .CK(osc_clk), .Q(d3[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i13.GSR = "ENABLED";
    FD1S3AX d3_i14 (.D(d3_71__N_562[14]), .CK(osc_clk), .Q(d3[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i14.GSR = "ENABLED";
    FD1S3AX d3_i15 (.D(d3_71__N_562[15]), .CK(osc_clk), .Q(d3[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i15.GSR = "ENABLED";
    FD1S3AX d3_i16 (.D(d3_71__N_562[16]), .CK(osc_clk), .Q(d3[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i16.GSR = "ENABLED";
    FD1S3AX d3_i17 (.D(d3_71__N_562[17]), .CK(osc_clk), .Q(d3[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i17.GSR = "ENABLED";
    FD1S3AX d3_i18 (.D(d3_71__N_562[18]), .CK(osc_clk), .Q(d3[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i18.GSR = "ENABLED";
    FD1S3AX d3_i19 (.D(d3_71__N_562[19]), .CK(osc_clk), .Q(d3[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i19.GSR = "ENABLED";
    FD1S3AX d3_i20 (.D(d3_71__N_562[20]), .CK(osc_clk), .Q(d3[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i20.GSR = "ENABLED";
    FD1S3AX d3_i21 (.D(d3_71__N_562[21]), .CK(osc_clk), .Q(d3[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i21.GSR = "ENABLED";
    FD1S3AX d3_i22 (.D(d3_71__N_562[22]), .CK(osc_clk), .Q(d3[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i22.GSR = "ENABLED";
    FD1S3AX d3_i23 (.D(d3_71__N_562[23]), .CK(osc_clk), .Q(d3[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i23.GSR = "ENABLED";
    FD1S3AX d3_i24 (.D(d3_71__N_562[24]), .CK(osc_clk), .Q(d3[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i24.GSR = "ENABLED";
    FD1S3AX d3_i25 (.D(d3_71__N_562[25]), .CK(osc_clk), .Q(d3[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i25.GSR = "ENABLED";
    FD1S3AX d3_i26 (.D(d3_71__N_562[26]), .CK(osc_clk), .Q(d3[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i26.GSR = "ENABLED";
    FD1S3AX d3_i27 (.D(d3_71__N_562[27]), .CK(osc_clk), .Q(d3[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i27.GSR = "ENABLED";
    FD1S3AX d3_i28 (.D(d3_71__N_562[28]), .CK(osc_clk), .Q(d3[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i28.GSR = "ENABLED";
    FD1S3AX d3_i29 (.D(d3_71__N_562[29]), .CK(osc_clk), .Q(d3[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i29.GSR = "ENABLED";
    FD1S3AX d3_i30 (.D(d3_71__N_562[30]), .CK(osc_clk), .Q(d3[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i30.GSR = "ENABLED";
    FD1S3AX d3_i31 (.D(d3_71__N_562[31]), .CK(osc_clk), .Q(d3[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i31.GSR = "ENABLED";
    FD1S3AX d3_i32 (.D(d3_71__N_562[32]), .CK(osc_clk), .Q(d3[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i32.GSR = "ENABLED";
    FD1S3AX d3_i33 (.D(d3_71__N_562[33]), .CK(osc_clk), .Q(d3[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i33.GSR = "ENABLED";
    FD1S3AX d3_i34 (.D(d3_71__N_562[34]), .CK(osc_clk), .Q(d3[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i34.GSR = "ENABLED";
    FD1S3AX d3_i35 (.D(d3_71__N_562[35]), .CK(osc_clk), .Q(d3[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i35.GSR = "ENABLED";
    FD1S3AX d3_i36 (.D(d3_71__N_562[36]), .CK(osc_clk), .Q(d3[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i36.GSR = "ENABLED";
    FD1S3AX d3_i37 (.D(d3_71__N_562[37]), .CK(osc_clk), .Q(d3[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i37.GSR = "ENABLED";
    FD1S3AX d3_i38 (.D(d3_71__N_562[38]), .CK(osc_clk), .Q(d3[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i38.GSR = "ENABLED";
    FD1S3AX d3_i39 (.D(d3_71__N_562[39]), .CK(osc_clk), .Q(d3[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i39.GSR = "ENABLED";
    FD1S3AX d3_i40 (.D(d3_71__N_562[40]), .CK(osc_clk), .Q(d3[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i40.GSR = "ENABLED";
    FD1S3AX d3_i41 (.D(d3_71__N_562[41]), .CK(osc_clk), .Q(d3[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i41.GSR = "ENABLED";
    FD1S3AX d3_i42 (.D(d3_71__N_562[42]), .CK(osc_clk), .Q(d3[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i42.GSR = "ENABLED";
    FD1S3AX d3_i43 (.D(d3_71__N_562[43]), .CK(osc_clk), .Q(d3[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i43.GSR = "ENABLED";
    FD1S3AX d3_i44 (.D(d3_71__N_562[44]), .CK(osc_clk), .Q(d3[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i44.GSR = "ENABLED";
    FD1S3AX d3_i45 (.D(d3_71__N_562[45]), .CK(osc_clk), .Q(d3[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i45.GSR = "ENABLED";
    FD1S3AX d3_i46 (.D(d3_71__N_562[46]), .CK(osc_clk), .Q(d3[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i46.GSR = "ENABLED";
    FD1S3AX d3_i47 (.D(d3_71__N_562[47]), .CK(osc_clk), .Q(d3[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i47.GSR = "ENABLED";
    FD1S3AX d3_i48 (.D(d3_71__N_562[48]), .CK(osc_clk), .Q(d3[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i48.GSR = "ENABLED";
    FD1S3AX d3_i49 (.D(d3_71__N_562[49]), .CK(osc_clk), .Q(d3[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i49.GSR = "ENABLED";
    FD1S3AX d3_i50 (.D(d3_71__N_562[50]), .CK(osc_clk), .Q(d3[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i50.GSR = "ENABLED";
    FD1S3AX d3_i51 (.D(d3_71__N_562[51]), .CK(osc_clk), .Q(d3[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i51.GSR = "ENABLED";
    FD1S3AX d3_i52 (.D(d3_71__N_562[52]), .CK(osc_clk), .Q(d3[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i52.GSR = "ENABLED";
    FD1S3AX d3_i53 (.D(d3_71__N_562[53]), .CK(osc_clk), .Q(d3[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i53.GSR = "ENABLED";
    FD1S3AX d3_i54 (.D(d3_71__N_562[54]), .CK(osc_clk), .Q(d3[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i54.GSR = "ENABLED";
    FD1S3AX d3_i55 (.D(d3_71__N_562[55]), .CK(osc_clk), .Q(d3[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i55.GSR = "ENABLED";
    FD1S3AX d3_i56 (.D(d3_71__N_562[56]), .CK(osc_clk), .Q(d3[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i56.GSR = "ENABLED";
    FD1S3AX d3_i57 (.D(d3_71__N_562[57]), .CK(osc_clk), .Q(d3[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i57.GSR = "ENABLED";
    FD1S3AX d3_i58 (.D(d3_71__N_562[58]), .CK(osc_clk), .Q(d3[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i58.GSR = "ENABLED";
    FD1S3AX d3_i59 (.D(d3_71__N_562[59]), .CK(osc_clk), .Q(d3[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i59.GSR = "ENABLED";
    FD1S3AX d3_i60 (.D(d3_71__N_562[60]), .CK(osc_clk), .Q(d3[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i60.GSR = "ENABLED";
    FD1S3AX d3_i61 (.D(d3_71__N_562[61]), .CK(osc_clk), .Q(d3[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i61.GSR = "ENABLED";
    FD1S3AX d3_i62 (.D(d3_71__N_562[62]), .CK(osc_clk), .Q(d3[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i62.GSR = "ENABLED";
    FD1S3AX d3_i63 (.D(d3_71__N_562[63]), .CK(osc_clk), .Q(d3[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i63.GSR = "ENABLED";
    FD1S3AX d3_i64 (.D(d3_71__N_562[64]), .CK(osc_clk), .Q(d3[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i64.GSR = "ENABLED";
    FD1S3AX d3_i65 (.D(d3_71__N_562[65]), .CK(osc_clk), .Q(d3[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i65.GSR = "ENABLED";
    FD1S3AX d3_i66 (.D(d3_71__N_562[66]), .CK(osc_clk), .Q(d3[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i66.GSR = "ENABLED";
    FD1S3AX d3_i67 (.D(d3_71__N_562[67]), .CK(osc_clk), .Q(d3[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i67.GSR = "ENABLED";
    FD1S3AX d3_i68 (.D(d3_71__N_562[68]), .CK(osc_clk), .Q(d3[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i68.GSR = "ENABLED";
    FD1S3AX d3_i69 (.D(d3_71__N_562[69]), .CK(osc_clk), .Q(d3[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i69.GSR = "ENABLED";
    FD1S3AX d3_i70 (.D(d3_71__N_562[70]), .CK(osc_clk), .Q(d3[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i70.GSR = "ENABLED";
    FD1S3AX d3_i71 (.D(d3_71__N_562[71]), .CK(osc_clk), .Q(d3[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i71.GSR = "ENABLED";
    FD1S3AX d4_i1 (.D(d4_71__N_634[1]), .CK(osc_clk), .Q(d4[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i1.GSR = "ENABLED";
    FD1S3AX d4_i2 (.D(d4_71__N_634[2]), .CK(osc_clk), .Q(d4[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i2.GSR = "ENABLED";
    FD1S3AX d4_i3 (.D(d4_71__N_634[3]), .CK(osc_clk), .Q(d4[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i3.GSR = "ENABLED";
    FD1S3AX d4_i4 (.D(d4_71__N_634[4]), .CK(osc_clk), .Q(d4[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i4.GSR = "ENABLED";
    FD1S3AX d4_i5 (.D(d4_71__N_634[5]), .CK(osc_clk), .Q(d4[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i5.GSR = "ENABLED";
    FD1S3AX d4_i6 (.D(d4_71__N_634[6]), .CK(osc_clk), .Q(d4[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i6.GSR = "ENABLED";
    FD1S3AX d4_i7 (.D(d4_71__N_634[7]), .CK(osc_clk), .Q(d4[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i7.GSR = "ENABLED";
    FD1S3AX d4_i8 (.D(d4_71__N_634[8]), .CK(osc_clk), .Q(d4[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i8.GSR = "ENABLED";
    FD1S3AX d4_i9 (.D(d4_71__N_634[9]), .CK(osc_clk), .Q(d4[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i9.GSR = "ENABLED";
    FD1S3AX d4_i10 (.D(d4_71__N_634[10]), .CK(osc_clk), .Q(d4[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i10.GSR = "ENABLED";
    FD1S3AX d4_i11 (.D(d4_71__N_634[11]), .CK(osc_clk), .Q(d4[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i11.GSR = "ENABLED";
    FD1S3AX d4_i12 (.D(d4_71__N_634[12]), .CK(osc_clk), .Q(d4[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i12.GSR = "ENABLED";
    FD1S3AX d4_i13 (.D(d4_71__N_634[13]), .CK(osc_clk), .Q(d4[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i13.GSR = "ENABLED";
    FD1S3AX d4_i14 (.D(d4_71__N_634[14]), .CK(osc_clk), .Q(d4[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i14.GSR = "ENABLED";
    FD1S3AX d4_i15 (.D(d4_71__N_634[15]), .CK(osc_clk), .Q(d4[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i15.GSR = "ENABLED";
    FD1S3AX d4_i16 (.D(d4_71__N_634[16]), .CK(osc_clk), .Q(d4[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i16.GSR = "ENABLED";
    FD1S3AX d4_i17 (.D(d4_71__N_634[17]), .CK(osc_clk), .Q(d4[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i17.GSR = "ENABLED";
    FD1S3AX d4_i18 (.D(d4_71__N_634[18]), .CK(osc_clk), .Q(d4[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i18.GSR = "ENABLED";
    FD1S3AX d4_i19 (.D(d4_71__N_634[19]), .CK(osc_clk), .Q(d4[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i19.GSR = "ENABLED";
    FD1S3AX d4_i20 (.D(d4_71__N_634[20]), .CK(osc_clk), .Q(d4[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i20.GSR = "ENABLED";
    FD1S3AX d4_i21 (.D(d4_71__N_634[21]), .CK(osc_clk), .Q(d4[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i21.GSR = "ENABLED";
    FD1S3AX d4_i22 (.D(d4_71__N_634[22]), .CK(osc_clk), .Q(d4[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i22.GSR = "ENABLED";
    FD1S3AX d4_i23 (.D(d4_71__N_634[23]), .CK(osc_clk), .Q(d4[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i23.GSR = "ENABLED";
    FD1S3AX d4_i24 (.D(d4_71__N_634[24]), .CK(osc_clk), .Q(d4[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i24.GSR = "ENABLED";
    FD1S3AX d4_i25 (.D(d4_71__N_634[25]), .CK(osc_clk), .Q(d4[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i25.GSR = "ENABLED";
    FD1S3AX d4_i26 (.D(d4_71__N_634[26]), .CK(osc_clk), .Q(d4[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i26.GSR = "ENABLED";
    FD1S3AX d4_i27 (.D(d4_71__N_634[27]), .CK(osc_clk), .Q(d4[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i27.GSR = "ENABLED";
    FD1S3AX d4_i28 (.D(d4_71__N_634[28]), .CK(osc_clk), .Q(d4[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i28.GSR = "ENABLED";
    FD1S3AX d4_i29 (.D(d4_71__N_634[29]), .CK(osc_clk), .Q(d4[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i29.GSR = "ENABLED";
    FD1S3AX d4_i30 (.D(d4_71__N_634[30]), .CK(osc_clk), .Q(d4[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i30.GSR = "ENABLED";
    FD1S3AX d4_i31 (.D(d4_71__N_634[31]), .CK(osc_clk), .Q(d4[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i31.GSR = "ENABLED";
    FD1S3AX d4_i32 (.D(d4_71__N_634[32]), .CK(osc_clk), .Q(d4[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i32.GSR = "ENABLED";
    FD1S3AX d4_i33 (.D(d4_71__N_634[33]), .CK(osc_clk), .Q(d4[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i33.GSR = "ENABLED";
    FD1S3AX d4_i34 (.D(d4_71__N_634[34]), .CK(osc_clk), .Q(d4[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i34.GSR = "ENABLED";
    FD1S3AX d4_i35 (.D(d4_71__N_634[35]), .CK(osc_clk), .Q(d4[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i35.GSR = "ENABLED";
    FD1S3AX d4_i36 (.D(d4_71__N_634[36]), .CK(osc_clk), .Q(d4[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i36.GSR = "ENABLED";
    FD1S3AX d4_i37 (.D(d4_71__N_634[37]), .CK(osc_clk), .Q(d4[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i37.GSR = "ENABLED";
    FD1S3AX d4_i38 (.D(d4_71__N_634[38]), .CK(osc_clk), .Q(d4[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i38.GSR = "ENABLED";
    FD1S3AX d4_i39 (.D(d4_71__N_634[39]), .CK(osc_clk), .Q(d4[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i39.GSR = "ENABLED";
    FD1S3AX d4_i40 (.D(d4_71__N_634[40]), .CK(osc_clk), .Q(d4[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i40.GSR = "ENABLED";
    FD1S3AX d4_i41 (.D(d4_71__N_634[41]), .CK(osc_clk), .Q(d4[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i41.GSR = "ENABLED";
    FD1S3AX d4_i42 (.D(d4_71__N_634[42]), .CK(osc_clk), .Q(d4[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i42.GSR = "ENABLED";
    FD1S3AX d4_i43 (.D(d4_71__N_634[43]), .CK(osc_clk), .Q(d4[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i43.GSR = "ENABLED";
    FD1S3AX d4_i44 (.D(d4_71__N_634[44]), .CK(osc_clk), .Q(d4[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i44.GSR = "ENABLED";
    FD1S3AX d4_i45 (.D(d4_71__N_634[45]), .CK(osc_clk), .Q(d4[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i45.GSR = "ENABLED";
    FD1S3AX d4_i46 (.D(d4_71__N_634[46]), .CK(osc_clk), .Q(d4[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i46.GSR = "ENABLED";
    FD1S3AX d4_i47 (.D(d4_71__N_634[47]), .CK(osc_clk), .Q(d4[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i47.GSR = "ENABLED";
    FD1S3AX d4_i48 (.D(d4_71__N_634[48]), .CK(osc_clk), .Q(d4[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i48.GSR = "ENABLED";
    FD1S3AX d4_i49 (.D(d4_71__N_634[49]), .CK(osc_clk), .Q(d4[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i49.GSR = "ENABLED";
    FD1S3AX d4_i50 (.D(d4_71__N_634[50]), .CK(osc_clk), .Q(d4[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i50.GSR = "ENABLED";
    FD1S3AX d4_i51 (.D(d4_71__N_634[51]), .CK(osc_clk), .Q(d4[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i51.GSR = "ENABLED";
    FD1S3AX d4_i52 (.D(d4_71__N_634[52]), .CK(osc_clk), .Q(d4[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i52.GSR = "ENABLED";
    FD1S3AX d4_i53 (.D(d4_71__N_634[53]), .CK(osc_clk), .Q(d4[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i53.GSR = "ENABLED";
    FD1S3AX d4_i54 (.D(d4_71__N_634[54]), .CK(osc_clk), .Q(d4[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i54.GSR = "ENABLED";
    FD1S3AX d4_i55 (.D(d4_71__N_634[55]), .CK(osc_clk), .Q(d4[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i55.GSR = "ENABLED";
    FD1S3AX d4_i56 (.D(d4_71__N_634[56]), .CK(osc_clk), .Q(d4[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i56.GSR = "ENABLED";
    FD1S3AX d4_i57 (.D(d4_71__N_634[57]), .CK(osc_clk), .Q(d4[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i57.GSR = "ENABLED";
    FD1S3AX d4_i58 (.D(d4_71__N_634[58]), .CK(osc_clk), .Q(d4[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i58.GSR = "ENABLED";
    FD1S3AX d4_i59 (.D(d4_71__N_634[59]), .CK(osc_clk), .Q(d4[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i59.GSR = "ENABLED";
    FD1S3AX d4_i60 (.D(d4_71__N_634[60]), .CK(osc_clk), .Q(d4[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i60.GSR = "ENABLED";
    FD1S3AX d4_i61 (.D(d4_71__N_634[61]), .CK(osc_clk), .Q(d4[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i61.GSR = "ENABLED";
    FD1S3AX d4_i62 (.D(d4_71__N_634[62]), .CK(osc_clk), .Q(d4[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i62.GSR = "ENABLED";
    FD1S3AX d4_i63 (.D(d4_71__N_634[63]), .CK(osc_clk), .Q(d4[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i63.GSR = "ENABLED";
    FD1S3AX d4_i64 (.D(d4_71__N_634[64]), .CK(osc_clk), .Q(d4[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i64.GSR = "ENABLED";
    FD1S3AX d4_i65 (.D(d4_71__N_634[65]), .CK(osc_clk), .Q(d4[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i65.GSR = "ENABLED";
    FD1S3AX d4_i66 (.D(d4_71__N_634[66]), .CK(osc_clk), .Q(d4[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i66.GSR = "ENABLED";
    FD1S3AX d4_i67 (.D(d4_71__N_634[67]), .CK(osc_clk), .Q(d4[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i67.GSR = "ENABLED";
    FD1S3AX d4_i68 (.D(d4_71__N_634[68]), .CK(osc_clk), .Q(d4[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i68.GSR = "ENABLED";
    FD1S3AX d4_i69 (.D(d4_71__N_634[69]), .CK(osc_clk), .Q(d4[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i69.GSR = "ENABLED";
    FD1S3AX d4_i70 (.D(d4_71__N_634[70]), .CK(osc_clk), .Q(d4[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i70.GSR = "ENABLED";
    FD1S3AX d4_i71 (.D(d4_71__N_634[71]), .CK(osc_clk), .Q(d4[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i71.GSR = "ENABLED";
    FD1S3AX d5_i1 (.D(d5_71__N_706[1]), .CK(osc_clk), .Q(d5[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i1.GSR = "ENABLED";
    FD1S3AX d5_i2 (.D(d5_71__N_706[2]), .CK(osc_clk), .Q(d5[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i2.GSR = "ENABLED";
    FD1S3AX d5_i3 (.D(d5_71__N_706[3]), .CK(osc_clk), .Q(d5[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i3.GSR = "ENABLED";
    FD1S3AX d5_i4 (.D(d5_71__N_706[4]), .CK(osc_clk), .Q(d5[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i4.GSR = "ENABLED";
    FD1S3AX d5_i5 (.D(d5_71__N_706[5]), .CK(osc_clk), .Q(d5[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i5.GSR = "ENABLED";
    FD1S3AX d5_i6 (.D(d5_71__N_706[6]), .CK(osc_clk), .Q(d5[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i6.GSR = "ENABLED";
    FD1S3AX d5_i7 (.D(d5_71__N_706[7]), .CK(osc_clk), .Q(d5[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i7.GSR = "ENABLED";
    FD1S3AX d5_i8 (.D(d5_71__N_706[8]), .CK(osc_clk), .Q(d5[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i8.GSR = "ENABLED";
    FD1S3AX d5_i9 (.D(d5_71__N_706[9]), .CK(osc_clk), .Q(d5[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i9.GSR = "ENABLED";
    FD1S3AX d5_i10 (.D(d5_71__N_706[10]), .CK(osc_clk), .Q(d5[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i10.GSR = "ENABLED";
    FD1S3AX d5_i11 (.D(d5_71__N_706[11]), .CK(osc_clk), .Q(d5[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i11.GSR = "ENABLED";
    FD1S3AX d5_i12 (.D(d5_71__N_706[12]), .CK(osc_clk), .Q(d5[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i12.GSR = "ENABLED";
    FD1S3AX d5_i13 (.D(d5_71__N_706[13]), .CK(osc_clk), .Q(d5[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i13.GSR = "ENABLED";
    FD1S3AX d5_i14 (.D(d5_71__N_706[14]), .CK(osc_clk), .Q(d5[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i14.GSR = "ENABLED";
    FD1S3AX d5_i15 (.D(d5_71__N_706[15]), .CK(osc_clk), .Q(d5[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i15.GSR = "ENABLED";
    FD1S3AX d5_i16 (.D(d5_71__N_706[16]), .CK(osc_clk), .Q(d5[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i16.GSR = "ENABLED";
    FD1S3AX d5_i17 (.D(d5_71__N_706[17]), .CK(osc_clk), .Q(d5[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i17.GSR = "ENABLED";
    FD1S3AX d5_i18 (.D(d5_71__N_706[18]), .CK(osc_clk), .Q(d5[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i18.GSR = "ENABLED";
    FD1S3AX d5_i19 (.D(d5_71__N_706[19]), .CK(osc_clk), .Q(d5[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i19.GSR = "ENABLED";
    FD1S3AX d5_i20 (.D(d5_71__N_706[20]), .CK(osc_clk), .Q(d5[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i20.GSR = "ENABLED";
    FD1S3AX d5_i21 (.D(d5_71__N_706[21]), .CK(osc_clk), .Q(d5[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i21.GSR = "ENABLED";
    FD1S3AX d5_i22 (.D(d5_71__N_706[22]), .CK(osc_clk), .Q(d5[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i22.GSR = "ENABLED";
    FD1S3AX d5_i23 (.D(d5_71__N_706[23]), .CK(osc_clk), .Q(d5[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i23.GSR = "ENABLED";
    FD1S3AX d5_i24 (.D(d5_71__N_706[24]), .CK(osc_clk), .Q(d5[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i24.GSR = "ENABLED";
    FD1S3AX d5_i25 (.D(d5_71__N_706[25]), .CK(osc_clk), .Q(d5[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i25.GSR = "ENABLED";
    FD1S3AX d5_i26 (.D(d5_71__N_706[26]), .CK(osc_clk), .Q(d5[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i26.GSR = "ENABLED";
    FD1S3AX d5_i27 (.D(d5_71__N_706[27]), .CK(osc_clk), .Q(d5[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i27.GSR = "ENABLED";
    FD1S3AX d5_i28 (.D(d5_71__N_706[28]), .CK(osc_clk), .Q(d5[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i28.GSR = "ENABLED";
    FD1S3AX d5_i29 (.D(d5_71__N_706[29]), .CK(osc_clk), .Q(d5[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i29.GSR = "ENABLED";
    FD1S3AX d5_i30 (.D(d5_71__N_706[30]), .CK(osc_clk), .Q(d5[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i30.GSR = "ENABLED";
    FD1S3AX d5_i31 (.D(d5_71__N_706[31]), .CK(osc_clk), .Q(d5[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i31.GSR = "ENABLED";
    FD1S3AX d5_i32 (.D(d5_71__N_706[32]), .CK(osc_clk), .Q(d5[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i32.GSR = "ENABLED";
    FD1S3AX d5_i33 (.D(d5_71__N_706[33]), .CK(osc_clk), .Q(d5[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i33.GSR = "ENABLED";
    FD1S3AX d5_i34 (.D(d5_71__N_706[34]), .CK(osc_clk), .Q(d5[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i34.GSR = "ENABLED";
    FD1S3AX d5_i35 (.D(d5_71__N_706[35]), .CK(osc_clk), .Q(d5[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i35.GSR = "ENABLED";
    FD1S3AX d5_i36 (.D(d5_71__N_706[36]), .CK(osc_clk), .Q(d5[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i36.GSR = "ENABLED";
    FD1S3AX d5_i37 (.D(d5_71__N_706[37]), .CK(osc_clk), .Q(d5[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i37.GSR = "ENABLED";
    FD1S3AX d5_i38 (.D(d5_71__N_706[38]), .CK(osc_clk), .Q(d5[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i38.GSR = "ENABLED";
    FD1S3AX d5_i39 (.D(d5_71__N_706[39]), .CK(osc_clk), .Q(d5[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i39.GSR = "ENABLED";
    FD1S3AX d5_i40 (.D(d5_71__N_706[40]), .CK(osc_clk), .Q(d5[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i40.GSR = "ENABLED";
    FD1S3AX d5_i41 (.D(d5_71__N_706[41]), .CK(osc_clk), .Q(d5[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i41.GSR = "ENABLED";
    FD1S3AX d5_i42 (.D(d5_71__N_706[42]), .CK(osc_clk), .Q(d5[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i42.GSR = "ENABLED";
    FD1S3AX d5_i43 (.D(d5_71__N_706[43]), .CK(osc_clk), .Q(d5[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i43.GSR = "ENABLED";
    FD1S3AX d5_i44 (.D(d5_71__N_706[44]), .CK(osc_clk), .Q(d5[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i44.GSR = "ENABLED";
    FD1S3AX d5_i45 (.D(d5_71__N_706[45]), .CK(osc_clk), .Q(d5[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i45.GSR = "ENABLED";
    FD1S3AX d5_i46 (.D(d5_71__N_706[46]), .CK(osc_clk), .Q(d5[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i46.GSR = "ENABLED";
    FD1S3AX d5_i47 (.D(d5_71__N_706[47]), .CK(osc_clk), .Q(d5[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i47.GSR = "ENABLED";
    FD1S3AX d5_i48 (.D(d5_71__N_706[48]), .CK(osc_clk), .Q(d5[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i48.GSR = "ENABLED";
    FD1S3AX d5_i49 (.D(d5_71__N_706[49]), .CK(osc_clk), .Q(d5[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i49.GSR = "ENABLED";
    FD1S3AX d5_i50 (.D(d5_71__N_706[50]), .CK(osc_clk), .Q(d5[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i50.GSR = "ENABLED";
    FD1S3AX d5_i51 (.D(d5_71__N_706[51]), .CK(osc_clk), .Q(d5[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i51.GSR = "ENABLED";
    FD1S3AX d5_i52 (.D(d5_71__N_706[52]), .CK(osc_clk), .Q(d5[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i52.GSR = "ENABLED";
    FD1S3AX d5_i53 (.D(d5_71__N_706[53]), .CK(osc_clk), .Q(d5[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i53.GSR = "ENABLED";
    FD1S3AX d5_i54 (.D(d5_71__N_706[54]), .CK(osc_clk), .Q(d5[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i54.GSR = "ENABLED";
    FD1S3AX d5_i55 (.D(d5_71__N_706[55]), .CK(osc_clk), .Q(d5[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i55.GSR = "ENABLED";
    FD1S3AX d5_i56 (.D(d5_71__N_706[56]), .CK(osc_clk), .Q(d5[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i56.GSR = "ENABLED";
    FD1S3AX d5_i57 (.D(d5_71__N_706[57]), .CK(osc_clk), .Q(d5[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i57.GSR = "ENABLED";
    FD1S3AX d5_i58 (.D(d5_71__N_706[58]), .CK(osc_clk), .Q(d5[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i58.GSR = "ENABLED";
    FD1S3AX d5_i59 (.D(d5_71__N_706[59]), .CK(osc_clk), .Q(d5[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i59.GSR = "ENABLED";
    FD1S3AX d5_i60 (.D(d5_71__N_706[60]), .CK(osc_clk), .Q(d5[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i60.GSR = "ENABLED";
    FD1S3AX d5_i61 (.D(d5_71__N_706[61]), .CK(osc_clk), .Q(d5[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i61.GSR = "ENABLED";
    FD1S3AX d5_i62 (.D(d5_71__N_706[62]), .CK(osc_clk), .Q(d5[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i62.GSR = "ENABLED";
    FD1S3AX d5_i63 (.D(d5_71__N_706[63]), .CK(osc_clk), .Q(d5[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i63.GSR = "ENABLED";
    FD1S3AX d5_i64 (.D(d5_71__N_706[64]), .CK(osc_clk), .Q(d5[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i64.GSR = "ENABLED";
    FD1S3AX d5_i65 (.D(d5_71__N_706[65]), .CK(osc_clk), .Q(d5[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i65.GSR = "ENABLED";
    FD1S3AX d5_i66 (.D(d5_71__N_706[66]), .CK(osc_clk), .Q(d5[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i66.GSR = "ENABLED";
    FD1S3AX d5_i67 (.D(d5_71__N_706[67]), .CK(osc_clk), .Q(d5[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i67.GSR = "ENABLED";
    FD1S3AX d5_i68 (.D(d5_71__N_706[68]), .CK(osc_clk), .Q(d5[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i68.GSR = "ENABLED";
    FD1S3AX d5_i69 (.D(d5_71__N_706[69]), .CK(osc_clk), .Q(d5[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i69.GSR = "ENABLED";
    FD1S3AX d5_i70 (.D(d5_71__N_706[70]), .CK(osc_clk), .Q(d5[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i70.GSR = "ENABLED";
    FD1S3AX d5_i71 (.D(d5_71__N_706[71]), .CK(osc_clk), .Q(d5[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i71.GSR = "ENABLED";
    FD1P3AX d6_i0_i1 (.D(d6_71__N_1459[1]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d6_i0_i2 (.D(d6_71__N_1459[2]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d6_i0_i3 (.D(d6_71__N_1459[3]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d6_i0_i4 (.D(d6_71__N_1459[4]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d6_i0_i5 (.D(d6_71__N_1459[5]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d6_i0_i6 (.D(d6_71__N_1459[6]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d6_i0_i7 (.D(d6_71__N_1459[7]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d6_i0_i8 (.D(d6_71__N_1459[8]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d6_i0_i9 (.D(d6_71__N_1459[9]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d6_i0_i10 (.D(d6_71__N_1459[10]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d6_i0_i11 (.D(d6_71__N_1459[11]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d6_i0_i12 (.D(d6_71__N_1459[12]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d6_i0_i13 (.D(d6_71__N_1459[13]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d6_i0_i14 (.D(d6_71__N_1459[14]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d6_i0_i15 (.D(d6_71__N_1459[15]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d6_i0_i16 (.D(d6_71__N_1459[16]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d6_i0_i17 (.D(d6_71__N_1459[17]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d6_i0_i18 (.D(d6_71__N_1459[18]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d6_i0_i19 (.D(d6_71__N_1459[19]), .SP(osc_clk_enable_160), .CK(osc_clk), 
            .Q(d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d6_i0_i20 (.D(d6_71__N_1459[20]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d6_i0_i21 (.D(d6_71__N_1459[21]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d6_i0_i22 (.D(d6_71__N_1459[22]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d6_i0_i23 (.D(d6_71__N_1459[23]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d6_i0_i24 (.D(d6_71__N_1459[24]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d6_i0_i25 (.D(d6_71__N_1459[25]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d6_i0_i26 (.D(d6_71__N_1459[26]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d6_i0_i27 (.D(d6_71__N_1459[27]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d6_i0_i28 (.D(d6_71__N_1459[28]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d6_i0_i29 (.D(d6_71__N_1459[29]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d6_i0_i30 (.D(d6_71__N_1459[30]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d6_i0_i31 (.D(d6_71__N_1459[31]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d6_i0_i32 (.D(d6_71__N_1459[32]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d6_i0_i33 (.D(d6_71__N_1459[33]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d6_i0_i34 (.D(d6_71__N_1459[34]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d6_i0_i35 (.D(d6_71__N_1459[35]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d6_i0_i36 (.D(d6_71__N_1459[36]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d6_i0_i37 (.D(d6_71__N_1459[37]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d6_i0_i38 (.D(d6_71__N_1459[38]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d6_i0_i39 (.D(d6_71__N_1459[39]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d6_i0_i40 (.D(d6_71__N_1459[40]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d6_i0_i41 (.D(d6_71__N_1459[41]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d6_i0_i42 (.D(d6_71__N_1459[42]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d6_i0_i43 (.D(d6_71__N_1459[43]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d6_i0_i44 (.D(d6_71__N_1459[44]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d6_i0_i45 (.D(d6_71__N_1459[45]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d6_i0_i46 (.D(d6_71__N_1459[46]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d6_i0_i47 (.D(d6_71__N_1459[47]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d6_i0_i48 (.D(d6_71__N_1459[48]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d6_i0_i49 (.D(d6_71__N_1459[49]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d6_i0_i50 (.D(d6_71__N_1459[50]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d6_i0_i51 (.D(d6_71__N_1459[51]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d6_i0_i52 (.D(d6_71__N_1459[52]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d6_i0_i53 (.D(d6_71__N_1459[53]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d6_i0_i54 (.D(d6_71__N_1459[54]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d6_i0_i55 (.D(d6_71__N_1459[55]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d6_i0_i56 (.D(d6_71__N_1459[56]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d6_i0_i57 (.D(d6_71__N_1459[57]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d6_i0_i58 (.D(d6_71__N_1459[58]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d6_i0_i59 (.D(d6_71__N_1459[59]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d6_i0_i60 (.D(d6_71__N_1459[60]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d6_i0_i61 (.D(d6_71__N_1459[61]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d6_i0_i62 (.D(d6_71__N_1459[62]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d6_i0_i63 (.D(d6_71__N_1459[63]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d6_i0_i64 (.D(d6_71__N_1459[64]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d6_i0_i65 (.D(d6_71__N_1459[65]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d6_i0_i66 (.D(d6_71__N_1459[66]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d6_i0_i67 (.D(d6_71__N_1459[67]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d6_i0_i68 (.D(d6_71__N_1459[68]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d6_i0_i69 (.D(d6_71__N_1459[69]), .SP(osc_clk_enable_210), .CK(osc_clk), 
            .Q(d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d6_i0_i70 (.D(d6_71__N_1459[70]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d6_i0_i71 (.D(d6_71__N_1459[71]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i1 (.D(d6[1]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i2 (.D(d6[2]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i3 (.D(d6[3]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i4 (.D(d6[4]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i5 (.D(d6[5]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i6 (.D(d6[6]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i7 (.D(d6[7]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i8 (.D(d6[8]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i9 (.D(d6[9]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i10 (.D(d6[10]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i11 (.D(d6[11]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i12 (.D(d6[12]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i13 (.D(d6[13]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i14 (.D(d6[14]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i15 (.D(d6[15]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i16 (.D(d6[16]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i17 (.D(d6[17]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i18 (.D(d6[18]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i19 (.D(d6[19]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i20 (.D(d6[20]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i21 (.D(d6[21]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i22 (.D(d6[22]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i23 (.D(d6[23]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i24 (.D(d6[24]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i25 (.D(d6[25]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i26 (.D(d6[26]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i27 (.D(d6[27]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i28 (.D(d6[28]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i29 (.D(d6[29]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i30 (.D(d6[30]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i31 (.D(d6[31]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i32 (.D(d6[32]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i33 (.D(d6[33]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i34 (.D(d6[34]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i35 (.D(d6[35]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i36 (.D(d6[36]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i37 (.D(d6[37]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i38 (.D(d6[38]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i39 (.D(d6[39]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i40 (.D(d6[40]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i41 (.D(d6[41]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i42 (.D(d6[42]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i43 (.D(d6[43]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i44 (.D(d6[44]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i45 (.D(d6[45]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i46 (.D(d6[46]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i47 (.D(d6[47]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i48 (.D(d6[48]), .SP(osc_clk_enable_260), .CK(osc_clk), 
            .Q(d_d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i49 (.D(d6[49]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d_d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i50 (.D(d6[50]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d_d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i51 (.D(d6[51]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d_d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i52 (.D(d6[52]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d_d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i53 (.D(d6[53]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d_d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i54 (.D(d6[54]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d_d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i55 (.D(d6[55]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d_d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i56 (.D(d6[56]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d_d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i57 (.D(d6[57]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d_d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i58 (.D(d6[58]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d_d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i59 (.D(d6[59]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d_d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i60 (.D(d6[60]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d_d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i61 (.D(d6[61]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d_d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i62 (.D(d6[62]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d_d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i63 (.D(d6[63]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d_d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i64 (.D(d6[64]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d_d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i65 (.D(d6[65]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d_d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i66 (.D(d6[66]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d_d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i67 (.D(d6[67]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d_d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i68 (.D(d6[68]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d_d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i69 (.D(d6[69]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d_d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i70 (.D(d6[70]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d_d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i71 (.D(d6[71]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d_d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d7_i0_i1 (.D(d7_71__N_1531[1]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d7_i0_i2 (.D(d7_71__N_1531[2]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d7_i0_i3 (.D(d7_71__N_1531[3]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d7_i0_i4 (.D(d7_71__N_1531[4]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d7_i0_i5 (.D(d7_71__N_1531[5]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d7_i0_i6 (.D(d7_71__N_1531[6]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d7_i0_i7 (.D(d7_71__N_1531[7]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d7_i0_i8 (.D(d7_71__N_1531[8]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d7_i0_i9 (.D(d7_71__N_1531[9]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d7_i0_i10 (.D(d7_71__N_1531[10]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d7_i0_i11 (.D(d7_71__N_1531[11]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d7_i0_i12 (.D(d7_71__N_1531[12]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d7_i0_i13 (.D(d7_71__N_1531[13]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d7_i0_i14 (.D(d7_71__N_1531[14]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d7_i0_i15 (.D(d7_71__N_1531[15]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d7_i0_i16 (.D(d7_71__N_1531[16]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d7_i0_i17 (.D(d7_71__N_1531[17]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d7_i0_i18 (.D(d7_71__N_1531[18]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d7_i0_i19 (.D(d7_71__N_1531[19]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d7_i0_i20 (.D(d7_71__N_1531[20]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d7_i0_i21 (.D(d7_71__N_1531[21]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d7_i0_i22 (.D(d7_71__N_1531[22]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d7_i0_i23 (.D(d7_71__N_1531[23]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d7_i0_i24 (.D(d7_71__N_1531[24]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d7_i0_i25 (.D(d7_71__N_1531[25]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d7_i0_i26 (.D(d7_71__N_1531[26]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d7_i0_i27 (.D(d7_71__N_1531[27]), .SP(osc_clk_enable_310), .CK(osc_clk), 
            .Q(d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d7_i0_i28 (.D(d7_71__N_1531[28]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d7_i0_i29 (.D(d7_71__N_1531[29]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d7_i0_i30 (.D(d7_71__N_1531[30]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d7_i0_i31 (.D(d7_71__N_1531[31]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d7_i0_i32 (.D(d7_71__N_1531[32]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d7_i0_i33 (.D(d7_71__N_1531[33]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d7_i0_i34 (.D(d7_71__N_1531[34]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d7_i0_i35 (.D(d7_71__N_1531[35]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d7_i0_i36 (.D(d7_71__N_1531[36]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d7_i0_i37 (.D(d7_71__N_1531[37]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d7_i0_i38 (.D(d7_71__N_1531[38]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d7_i0_i39 (.D(d7_71__N_1531[39]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d7_i0_i40 (.D(d7_71__N_1531[40]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d7_i0_i41 (.D(d7_71__N_1531[41]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d7_i0_i42 (.D(d7_71__N_1531[42]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d7_i0_i43 (.D(d7_71__N_1531[43]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d7_i0_i44 (.D(d7_71__N_1531[44]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d7_i0_i45 (.D(d7_71__N_1531[45]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d7_i0_i46 (.D(d7_71__N_1531[46]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d7_i0_i47 (.D(d7_71__N_1531[47]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d7_i0_i48 (.D(d7_71__N_1531[48]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d7_i0_i49 (.D(d7_71__N_1531[49]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d7_i0_i50 (.D(d7_71__N_1531[50]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d7_i0_i51 (.D(d7_71__N_1531[51]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d7_i0_i52 (.D(d7_71__N_1531[52]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d7_i0_i53 (.D(d7_71__N_1531[53]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d7_i0_i54 (.D(d7_71__N_1531[54]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d7_i0_i55 (.D(d7_71__N_1531[55]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d7_i0_i56 (.D(d7_71__N_1531[56]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d7_i0_i57 (.D(d7_71__N_1531[57]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d7_i0_i58 (.D(d7_71__N_1531[58]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d7_i0_i59 (.D(d7_71__N_1531[59]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d7_i0_i60 (.D(d7_71__N_1531[60]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d7_i0_i61 (.D(d7_71__N_1531[61]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d7_i0_i62 (.D(d7_71__N_1531[62]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d7_i0_i63 (.D(d7_71__N_1531[63]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d7_i0_i64 (.D(d7_71__N_1531[64]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d7_i0_i65 (.D(d7_71__N_1531[65]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d7_i0_i66 (.D(d7_71__N_1531[66]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d7_i0_i67 (.D(d7_71__N_1531[67]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d7_i0_i68 (.D(d7_71__N_1531[68]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d7_i0_i69 (.D(d7_71__N_1531[69]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d7_i0_i70 (.D(d7_71__N_1531[70]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d7_i0_i71 (.D(d7_71__N_1531[71]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i1 (.D(d7[1]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d_d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i2 (.D(d7[2]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d_d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i3 (.D(d7[3]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d_d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i4 (.D(d7[4]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d_d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i5 (.D(d7[5]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d_d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i6 (.D(d7[6]), .SP(osc_clk_enable_360), .CK(osc_clk), 
            .Q(d_d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i7 (.D(d7[7]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i8 (.D(d7[8]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i9 (.D(d7[9]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i10 (.D(d7[10]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i11 (.D(d7[11]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i12 (.D(d7[12]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i13 (.D(d7[13]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i14 (.D(d7[14]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i15 (.D(d7[15]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i16 (.D(d7[16]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i17 (.D(d7[17]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i18 (.D(d7[18]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i19 (.D(d7[19]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i20 (.D(d7[20]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i21 (.D(d7[21]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i22 (.D(d7[22]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i23 (.D(d7[23]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i24 (.D(d7[24]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i25 (.D(d7[25]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i26 (.D(d7[26]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i27 (.D(d7[27]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i28 (.D(d7[28]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i29 (.D(d7[29]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i30 (.D(d7[30]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i31 (.D(d7[31]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i32 (.D(d7[32]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i33 (.D(d7[33]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i34 (.D(d7[34]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i35 (.D(d7[35]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i36 (.D(d7[36]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i37 (.D(d7[37]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i38 (.D(d7[38]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i39 (.D(d7[39]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i40 (.D(d7[40]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i41 (.D(d7[41]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i42 (.D(d7[42]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i43 (.D(d7[43]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i44 (.D(d7[44]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i45 (.D(d7[45]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i46 (.D(d7[46]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i47 (.D(d7[47]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i48 (.D(d7[48]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i49 (.D(d7[49]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i50 (.D(d7[50]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i51 (.D(d7[51]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i52 (.D(d7[52]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i53 (.D(d7[53]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i54 (.D(d7[54]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i55 (.D(d7[55]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i56 (.D(d7[56]), .SP(osc_clk_enable_410), .CK(osc_clk), 
            .Q(d_d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i57 (.D(d7[57]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d_d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i58 (.D(d7[58]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d_d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i59 (.D(d7[59]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d_d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i60 (.D(d7[60]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d_d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i61 (.D(d7[61]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d_d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i62 (.D(d7[62]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d_d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i63 (.D(d7[63]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d_d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i64 (.D(d7[64]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d_d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i65 (.D(d7[65]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d_d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i66 (.D(d7[66]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d_d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i67 (.D(d7[67]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d_d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i68 (.D(d7[68]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d_d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i69 (.D(d7[69]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d_d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i70 (.D(d7[70]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d_d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i71 (.D(d7[71]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d_d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d8_i0_i1 (.D(d8_71__N_1603[1]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d8_i0_i2 (.D(d8_71__N_1603[2]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d8_i0_i3 (.D(d8_71__N_1603[3]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d8_i0_i4 (.D(d8_71__N_1603[4]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d8_i0_i5 (.D(d8_71__N_1603[5]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d8_i0_i6 (.D(d8_71__N_1603[6]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d8_i0_i7 (.D(d8_71__N_1603[7]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d8_i0_i8 (.D(d8_71__N_1603[8]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d8_i0_i9 (.D(d8_71__N_1603[9]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d8_i0_i10 (.D(d8_71__N_1603[10]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d8_i0_i11 (.D(d8_71__N_1603[11]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d8_i0_i12 (.D(d8_71__N_1603[12]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d8_i0_i13 (.D(d8_71__N_1603[13]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d8_i0_i14 (.D(d8_71__N_1603[14]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d8_i0_i15 (.D(d8_71__N_1603[15]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d8_i0_i16 (.D(d8_71__N_1603[16]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d8_i0_i17 (.D(d8_71__N_1603[17]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d8_i0_i18 (.D(d8_71__N_1603[18]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d8_i0_i19 (.D(d8_71__N_1603[19]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d8_i0_i20 (.D(d8_71__N_1603[20]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d8_i0_i21 (.D(d8_71__N_1603[21]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d8_i0_i22 (.D(d8_71__N_1603[22]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d8_i0_i23 (.D(d8_71__N_1603[23]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d8_i0_i24 (.D(d8_71__N_1603[24]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d8_i0_i25 (.D(d8_71__N_1603[25]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d8_i0_i26 (.D(d8_71__N_1603[26]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d8_i0_i27 (.D(d8_71__N_1603[27]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d8_i0_i28 (.D(d8_71__N_1603[28]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d8_i0_i29 (.D(d8_71__N_1603[29]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d8_i0_i30 (.D(d8_71__N_1603[30]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d8_i0_i31 (.D(d8_71__N_1603[31]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d8_i0_i32 (.D(d8_71__N_1603[32]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d8_i0_i33 (.D(d8_71__N_1603[33]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d8_i0_i34 (.D(d8_71__N_1603[34]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d8_i0_i35 (.D(d8_71__N_1603[35]), .SP(osc_clk_enable_460), .CK(osc_clk), 
            .Q(d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d8_i0_i36 (.D(d8_71__N_1603[36]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d8_i0_i37 (.D(d8_71__N_1603[37]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d8_i0_i38 (.D(d8_71__N_1603[38]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d8_i0_i39 (.D(d8_71__N_1603[39]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d8_i0_i40 (.D(d8_71__N_1603[40]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d8_i0_i41 (.D(d8_71__N_1603[41]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d8_i0_i42 (.D(d8_71__N_1603[42]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d8_i0_i43 (.D(d8_71__N_1603[43]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d8_i0_i44 (.D(d8_71__N_1603[44]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d8_i0_i45 (.D(d8_71__N_1603[45]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d8_i0_i46 (.D(d8_71__N_1603[46]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d8_i0_i47 (.D(d8_71__N_1603[47]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d8_i0_i48 (.D(d8_71__N_1603[48]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d8_i0_i49 (.D(d8_71__N_1603[49]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d8_i0_i50 (.D(d8_71__N_1603[50]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d8_i0_i51 (.D(d8_71__N_1603[51]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d8_i0_i52 (.D(d8_71__N_1603[52]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d8_i0_i53 (.D(d8_71__N_1603[53]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d8_i0_i54 (.D(d8_71__N_1603[54]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d8_i0_i55 (.D(d8_71__N_1603[55]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d8_i0_i56 (.D(d8_71__N_1603[56]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d8_i0_i57 (.D(d8_71__N_1603[57]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d8_i0_i58 (.D(d8_71__N_1603[58]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d8_i0_i59 (.D(d8_71__N_1603[59]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d8_i0_i60 (.D(d8_71__N_1603[60]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d8_i0_i61 (.D(d8_71__N_1603[61]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d8_i0_i62 (.D(d8_71__N_1603[62]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d8_i0_i63 (.D(d8_71__N_1603[63]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d8_i0_i64 (.D(d8_71__N_1603[64]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d8_i0_i65 (.D(d8_71__N_1603[65]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d8_i0_i66 (.D(d8_71__N_1603[66]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d8_i0_i67 (.D(d8_71__N_1603[67]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d8_i0_i68 (.D(d8_71__N_1603[68]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d8_i0_i69 (.D(d8_71__N_1603[69]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d8_i0_i70 (.D(d8_71__N_1603[70]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d8_i0_i71 (.D(d8_71__N_1603[71]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i1 (.D(d8[1]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d_d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i2 (.D(d8[2]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d_d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i3 (.D(d8[3]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d_d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i4 (.D(d8[4]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d_d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i5 (.D(d8[5]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d_d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i6 (.D(d8[6]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d_d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i7 (.D(d8[7]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d_d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i8 (.D(d8[8]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d_d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i9 (.D(d8[9]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d_d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i10 (.D(d8[10]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d_d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i11 (.D(d8[11]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d_d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i12 (.D(d8[12]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d_d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i13 (.D(d8[13]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d_d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i14 (.D(d8[14]), .SP(osc_clk_enable_510), .CK(osc_clk), 
            .Q(d_d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i15 (.D(d8[15]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i16 (.D(d8[16]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i17 (.D(d8[17]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i18 (.D(d8[18]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i19 (.D(d8[19]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i20 (.D(d8[20]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i21 (.D(d8[21]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i22 (.D(d8[22]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i23 (.D(d8[23]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i24 (.D(d8[24]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i25 (.D(d8[25]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i26 (.D(d8[26]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i27 (.D(d8[27]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i28 (.D(d8[28]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i29 (.D(d8[29]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i30 (.D(d8[30]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i31 (.D(d8[31]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i32 (.D(d8[32]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i33 (.D(d8[33]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i34 (.D(d8[34]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i35 (.D(d8[35]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i36 (.D(d8[36]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i37 (.D(d8[37]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i38 (.D(d8[38]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i39 (.D(d8[39]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i40 (.D(d8[40]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i41 (.D(d8[41]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i42 (.D(d8[42]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i43 (.D(d8[43]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i44 (.D(d8[44]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i45 (.D(d8[45]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i46 (.D(d8[46]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i47 (.D(d8[47]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i48 (.D(d8[48]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i49 (.D(d8[49]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i50 (.D(d8[50]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i51 (.D(d8[51]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i52 (.D(d8[52]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i53 (.D(d8[53]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i54 (.D(d8[54]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i55 (.D(d8[55]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i56 (.D(d8[56]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i57 (.D(d8[57]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i58 (.D(d8[58]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i59 (.D(d8[59]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i60 (.D(d8[60]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i61 (.D(d8[61]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i62 (.D(d8[62]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i63 (.D(d8[63]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i64 (.D(d8[64]), .SP(osc_clk_enable_560), .CK(osc_clk), 
            .Q(d_d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i65 (.D(d8[65]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d_d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i66 (.D(d8[66]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d_d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i67 (.D(d8[67]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d_d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i68 (.D(d8[68]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d_d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i69 (.D(d8[69]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d_d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i70 (.D(d8[70]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d_d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i71 (.D(d8[71]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d_d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d9_i0_i1 (.D(d9_71__N_1675[1]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d9_i0_i2 (.D(d9_71__N_1675[2]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d9_i0_i3 (.D(d9_71__N_1675[3]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d9_i0_i4 (.D(d9_71__N_1675[4]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d9_i0_i5 (.D(d9_71__N_1675[5]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d9_i0_i6 (.D(d9_71__N_1675[6]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d9_i0_i7 (.D(d9_71__N_1675[7]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d9_i0_i8 (.D(d9_71__N_1675[8]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d9_i0_i9 (.D(d9_71__N_1675[9]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d9_i0_i10 (.D(d9_71__N_1675[10]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d9_i0_i11 (.D(d9_71__N_1675[11]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d9_i0_i12 (.D(d9_71__N_1675[12]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d9_i0_i13 (.D(d9_71__N_1675[13]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d9_i0_i14 (.D(d9_71__N_1675[14]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d9_i0_i15 (.D(d9_71__N_1675[15]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d9_i0_i16 (.D(d9_71__N_1675[16]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d9_i0_i17 (.D(d9_71__N_1675[17]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d9_i0_i18 (.D(d9_71__N_1675[18]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d9_i0_i19 (.D(d9_71__N_1675[19]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d9_i0_i20 (.D(d9_71__N_1675[20]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d9_i0_i21 (.D(d9_71__N_1675[21]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d9_i0_i22 (.D(d9_71__N_1675[22]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d9_i0_i23 (.D(d9_71__N_1675[23]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d9_i0_i24 (.D(d9_71__N_1675[24]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d9_i0_i25 (.D(d9_71__N_1675[25]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d9_i0_i26 (.D(d9_71__N_1675[26]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d9_i0_i27 (.D(d9_71__N_1675[27]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d9_i0_i28 (.D(d9_71__N_1675[28]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d9_i0_i29 (.D(d9_71__N_1675[29]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d9_i0_i30 (.D(d9_71__N_1675[30]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d9_i0_i31 (.D(d9_71__N_1675[31]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d9_i0_i32 (.D(d9_71__N_1675[32]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d9_i0_i33 (.D(d9_71__N_1675[33]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d9_i0_i34 (.D(d9_71__N_1675[34]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d9_i0_i35 (.D(d9_71__N_1675[35]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d9_i0_i36 (.D(d9_71__N_1675[36]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d9_i0_i37 (.D(d9_71__N_1675[37]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d9_i0_i38 (.D(d9_71__N_1675[38]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d9_i0_i39 (.D(d9_71__N_1675[39]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d9_i0_i40 (.D(d9_71__N_1675[40]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d9_i0_i41 (.D(d9_71__N_1675[41]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d9_i0_i42 (.D(d9_71__N_1675[42]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d9_i0_i43 (.D(d9_71__N_1675[43]), .SP(osc_clk_enable_610), .CK(osc_clk), 
            .Q(d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d9_i0_i44 (.D(d9_71__N_1675[44]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d9_i0_i45 (.D(d9_71__N_1675[45]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d9_i0_i46 (.D(d9_71__N_1675[46]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d9_i0_i47 (.D(d9_71__N_1675[47]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d9_i0_i48 (.D(d9_71__N_1675[48]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d9_i0_i49 (.D(d9_71__N_1675[49]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d9_i0_i50 (.D(d9_71__N_1675[50]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d9_i0_i51 (.D(d9_71__N_1675[51]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d9_i0_i52 (.D(d9_71__N_1675[52]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d9_i0_i53 (.D(d9_71__N_1675[53]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d9_i0_i54 (.D(d9_71__N_1675[54]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d9_i0_i55 (.D(d9_71__N_1675[55]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d9_i0_i56 (.D(d9_71__N_1675[56]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d9_i0_i57 (.D(d9_71__N_1675[57]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d9_i0_i58 (.D(d9_71__N_1675[58]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d9_i0_i59 (.D(d9_71__N_1675[59]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d9_i0_i60 (.D(d9_71__N_1675[60]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d9_i0_i61 (.D(d9_71__N_1675[61]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d9_i0_i62 (.D(d9_71__N_1675[62]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d9_i0_i63 (.D(d9_71__N_1675[63]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d9_i0_i64 (.D(d9_71__N_1675[64]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d9_i0_i65 (.D(d9_71__N_1675[65]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d9_i0_i66 (.D(d9_71__N_1675[66]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d9_i0_i67 (.D(d9_71__N_1675[67]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d9_i0_i68 (.D(d9_71__N_1675[68]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d9_i0_i69 (.D(d9_71__N_1675[69]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d9_i0_i70 (.D(d9_71__N_1675[70]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d9_i0_i71 (.D(d9_71__N_1675[71]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i1 (.D(d9[1]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d_d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i2 (.D(d9[2]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d_d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i3 (.D(d9[3]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d_d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i4 (.D(d9[4]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d_d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i5 (.D(d9[5]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d_d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i6 (.D(d9[6]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d_d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i7 (.D(d9[7]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d_d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i8 (.D(d9[8]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d_d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i9 (.D(d9[9]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d_d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i10 (.D(d9[10]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d_d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i11 (.D(d9[11]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d_d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i12 (.D(d9[12]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d_d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i13 (.D(d9[13]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d_d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i14 (.D(d9[14]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d_d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i15 (.D(d9[15]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d_d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i16 (.D(d9[16]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d_d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i17 (.D(d9[17]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d_d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i18 (.D(d9[18]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d_d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i19 (.D(d9[19]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d_d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i20 (.D(d9[20]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d_d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i21 (.D(d9[21]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d_d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i22 (.D(d9[22]), .SP(osc_clk_enable_660), .CK(osc_clk), 
            .Q(d_d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i23 (.D(d9[23]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i24 (.D(d9[24]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i25 (.D(d9[25]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i26 (.D(d9[26]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i27 (.D(d9[27]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i28 (.D(d9[28]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i29 (.D(d9[29]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i30 (.D(d9[30]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i31 (.D(d9[31]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i32 (.D(d9[32]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i33 (.D(d9[33]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i34 (.D(d9[34]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i35 (.D(d9[35]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i36 (.D(d9[36]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i37 (.D(d9[37]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i38 (.D(d9[38]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i39 (.D(d9[39]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i40 (.D(d9[40]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i41 (.D(d9[41]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i42 (.D(d9[42]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i43 (.D(d9[43]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i44 (.D(d9[44]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i45 (.D(d9[45]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i46 (.D(d9[46]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i47 (.D(d9[47]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i48 (.D(d9[48]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i49 (.D(d9[49]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i50 (.D(d9[50]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i51 (.D(d9[51]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i52 (.D(d9[52]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i53 (.D(d9[53]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i54 (.D(d9[54]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i55 (.D(d9[55]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i56 (.D(d9[56]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i57 (.D(d9[57]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i58 (.D(d9[58]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i59 (.D(d9[59]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i60 (.D(d9[60]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i61 (.D(d9[61]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i62 (.D(d9[62]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i63 (.D(d9[63]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i64 (.D(d9[64]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i65 (.D(d9[65]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i66 (.D(d9[66]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i67 (.D(d9[67]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i68 (.D(d9[68]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i69 (.D(d9[69]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i70 (.D(d9[70]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i71 (.D(d9[71]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d_d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d10__i2 (.D(d10_71__N_1747[57]), .SP(osc_clk_enable_710), .CK(osc_clk), 
            .Q(d10[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i2.GSR = "ENABLED";
    FD1P3AX d10__i3 (.D(d10_71__N_1747[58]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i3.GSR = "ENABLED";
    FD1P3AX d10__i4 (.D(d10_71__N_1747[59]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i4.GSR = "ENABLED";
    FD1P3AX d10__i5 (.D(d10_71__N_1747[60]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i5.GSR = "ENABLED";
    FD1P3AX d10__i6 (.D(d10_71__N_1747[61]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i6.GSR = "ENABLED";
    FD1P3AX d10__i7 (.D(d10_71__N_1747[62]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i7.GSR = "ENABLED";
    FD1P3AX d10__i8 (.D(d10_71__N_1747[63]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i8.GSR = "ENABLED";
    FD1P3AX d10__i9 (.D(d10_71__N_1747[64]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i9.GSR = "ENABLED";
    FD1P3AX d10__i10 (.D(d10_71__N_1747[65]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i10.GSR = "ENABLED";
    FD1P3AX d10__i11 (.D(d10_71__N_1747[66]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i11.GSR = "ENABLED";
    FD1P3AX d10__i12 (.D(d10_71__N_1747[67]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i12.GSR = "ENABLED";
    FD1P3AX d10__i13 (.D(d10_71__N_1747[68]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i13.GSR = "ENABLED";
    FD1P3AX d10__i14 (.D(d10_71__N_1747[69]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i14.GSR = "ENABLED";
    FD1P3AX d10__i15 (.D(d10_71__N_1747[70]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i15.GSR = "ENABLED";
    FD1P3AX d10__i16 (.D(d10_71__N_1747[71]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i16.GSR = "ENABLED";
    FD1P3AX d_out_i0_i1 (.D(d_out_11__N_1819[1]), .SP(v_comb), .CK(osc_clk), 
            .Q(\CIC1_outSin[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i1.GSR = "ENABLED";
    FD1P3AX d_out_i0_i2 (.D(d_out_11__N_1819[2]), .SP(v_comb), .CK(osc_clk), 
            .Q(\CIC1_outSin[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i2.GSR = "ENABLED";
    FD1P3AX d_out_i0_i3 (.D(d_out_11__N_1819[3]), .SP(v_comb), .CK(osc_clk), 
            .Q(\CIC1_outSin[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i3.GSR = "ENABLED";
    FD1P3AX d_out_i0_i4 (.D(d_out_11__N_1819[4]), .SP(v_comb), .CK(osc_clk), 
            .Q(\CIC1_outSin[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i4.GSR = "ENABLED";
    FD1P3AX d_out_i0_i5 (.D(d_out_11__N_1819[5]), .SP(v_comb), .CK(osc_clk), 
            .Q(\CIC1_outSin[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i5.GSR = "ENABLED";
    FD1P3AX d_out_i0_i6 (.D(d_out_11__N_1819[6]), .SP(v_comb), .CK(osc_clk), 
            .Q(MYLED_c_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i6.GSR = "ENABLED";
    FD1P3AX d_out_i0_i7 (.D(d_out_11__N_1819[7]), .SP(v_comb), .CK(osc_clk), 
            .Q(MYLED_c_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i7.GSR = "ENABLED";
    FD1P3AX d_out_i0_i8 (.D(d_out_11__N_1819[8]), .SP(v_comb), .CK(osc_clk), 
            .Q(MYLED_c_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i8.GSR = "ENABLED";
    FD1P3AX d_out_i0_i9 (.D(d_out_11__N_1819[9]), .SP(v_comb), .CK(osc_clk), 
            .Q(MYLED_c_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i9.GSR = "ENABLED";
    FD1P3AX d_out_i0_i10 (.D(d_out_11__N_1819[10]), .SP(v_comb), .CK(osc_clk), 
            .Q(MYLED_c_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i10.GSR = "ENABLED";
    FD1P3AX d_out_i0_i11 (.D(d_out_11__N_1819[11]), .SP(v_comb), .CK(osc_clk), 
            .Q(MYLED_c_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i11.GSR = "ENABLED";
    FD1S3AX d1_i1 (.D(d1_71__N_418[1]), .CK(osc_clk), .Q(d1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i1.GSR = "ENABLED";
    FD1S3AX d1_i2 (.D(d1_71__N_418[2]), .CK(osc_clk), .Q(d1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i2.GSR = "ENABLED";
    FD1S3AX d1_i3 (.D(d1_71__N_418[3]), .CK(osc_clk), .Q(d1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i3.GSR = "ENABLED";
    FD1S3AX d1_i4 (.D(d1_71__N_418[4]), .CK(osc_clk), .Q(d1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i4.GSR = "ENABLED";
    FD1S3AX d1_i5 (.D(d1_71__N_418[5]), .CK(osc_clk), .Q(d1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i5.GSR = "ENABLED";
    FD1S3AX d1_i6 (.D(d1_71__N_418[6]), .CK(osc_clk), .Q(d1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i6.GSR = "ENABLED";
    FD1S3AX d1_i7 (.D(d1_71__N_418[7]), .CK(osc_clk), .Q(d1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i7.GSR = "ENABLED";
    FD1S3AX d1_i8 (.D(d1_71__N_418[8]), .CK(osc_clk), .Q(d1[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i8.GSR = "ENABLED";
    FD1S3AX d1_i9 (.D(d1_71__N_418[9]), .CK(osc_clk), .Q(d1[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i9.GSR = "ENABLED";
    FD1S3AX d1_i10 (.D(d1_71__N_418[10]), .CK(osc_clk), .Q(d1[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i10.GSR = "ENABLED";
    FD1S3AX d1_i11 (.D(d1_71__N_418[11]), .CK(osc_clk), .Q(d1[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i11.GSR = "ENABLED";
    FD1S3AX d1_i12 (.D(d1_71__N_418[12]), .CK(osc_clk), .Q(d1[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i12.GSR = "ENABLED";
    FD1S3AX d1_i13 (.D(d1_71__N_418[13]), .CK(osc_clk), .Q(d1[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i13.GSR = "ENABLED";
    FD1S3AX d1_i14 (.D(d1_71__N_418[14]), .CK(osc_clk), .Q(d1[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i14.GSR = "ENABLED";
    FD1S3AX d1_i15 (.D(d1_71__N_418[15]), .CK(osc_clk), .Q(d1[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i15.GSR = "ENABLED";
    FD1S3AX d1_i16 (.D(d1_71__N_418[16]), .CK(osc_clk), .Q(d1[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i16.GSR = "ENABLED";
    FD1S3AX d1_i17 (.D(d1_71__N_418[17]), .CK(osc_clk), .Q(d1[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i17.GSR = "ENABLED";
    FD1S3AX d1_i18 (.D(d1_71__N_418[18]), .CK(osc_clk), .Q(d1[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i18.GSR = "ENABLED";
    FD1S3AX d1_i19 (.D(d1_71__N_418[19]), .CK(osc_clk), .Q(d1[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i19.GSR = "ENABLED";
    FD1S3AX d1_i20 (.D(d1_71__N_418[20]), .CK(osc_clk), .Q(d1[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i20.GSR = "ENABLED";
    FD1S3AX d1_i21 (.D(d1_71__N_418[21]), .CK(osc_clk), .Q(d1[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i21.GSR = "ENABLED";
    FD1S3AX d1_i22 (.D(d1_71__N_418[22]), .CK(osc_clk), .Q(d1[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i22.GSR = "ENABLED";
    FD1S3AX d1_i23 (.D(d1_71__N_418[23]), .CK(osc_clk), .Q(d1[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i23.GSR = "ENABLED";
    FD1S3AX d1_i24 (.D(d1_71__N_418[24]), .CK(osc_clk), .Q(d1[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i24.GSR = "ENABLED";
    FD1S3AX d1_i25 (.D(d1_71__N_418[25]), .CK(osc_clk), .Q(d1[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i25.GSR = "ENABLED";
    FD1S3AX d1_i26 (.D(d1_71__N_418[26]), .CK(osc_clk), .Q(d1[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i26.GSR = "ENABLED";
    FD1S3AX d1_i27 (.D(d1_71__N_418[27]), .CK(osc_clk), .Q(d1[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i27.GSR = "ENABLED";
    FD1S3AX d1_i28 (.D(d1_71__N_418[28]), .CK(osc_clk), .Q(d1[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i28.GSR = "ENABLED";
    FD1S3AX d1_i29 (.D(d1_71__N_418[29]), .CK(osc_clk), .Q(d1[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i29.GSR = "ENABLED";
    FD1S3AX d1_i30 (.D(d1_71__N_418[30]), .CK(osc_clk), .Q(d1[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i30.GSR = "ENABLED";
    FD1S3AX d1_i31 (.D(d1_71__N_418[31]), .CK(osc_clk), .Q(d1[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i31.GSR = "ENABLED";
    FD1S3AX d1_i32 (.D(d1_71__N_418[32]), .CK(osc_clk), .Q(d1[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i32.GSR = "ENABLED";
    FD1S3AX d1_i33 (.D(d1_71__N_418[33]), .CK(osc_clk), .Q(d1[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i33.GSR = "ENABLED";
    FD1S3AX d1_i34 (.D(d1_71__N_418[34]), .CK(osc_clk), .Q(d1[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i34.GSR = "ENABLED";
    FD1S3AX d1_i35 (.D(d1_71__N_418[35]), .CK(osc_clk), .Q(d1[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i35.GSR = "ENABLED";
    FD1S3AX d1_i36 (.D(d1_71__N_418[36]), .CK(osc_clk), .Q(d1[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i36.GSR = "ENABLED";
    FD1S3AX d1_i37 (.D(d1_71__N_418[37]), .CK(osc_clk), .Q(d1[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i37.GSR = "ENABLED";
    FD1S3AX d1_i38 (.D(d1_71__N_418[38]), .CK(osc_clk), .Q(d1[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i38.GSR = "ENABLED";
    FD1S3AX d1_i39 (.D(d1_71__N_418[39]), .CK(osc_clk), .Q(d1[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i39.GSR = "ENABLED";
    FD1S3AX d1_i40 (.D(d1_71__N_418[40]), .CK(osc_clk), .Q(d1[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i40.GSR = "ENABLED";
    FD1S3AX d1_i41 (.D(d1_71__N_418[41]), .CK(osc_clk), .Q(d1[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i41.GSR = "ENABLED";
    FD1S3AX d1_i42 (.D(d1_71__N_418[42]), .CK(osc_clk), .Q(d1[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i42.GSR = "ENABLED";
    FD1S3AX d1_i43 (.D(d1_71__N_418[43]), .CK(osc_clk), .Q(d1[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i43.GSR = "ENABLED";
    FD1S3AX d1_i44 (.D(d1_71__N_418[44]), .CK(osc_clk), .Q(d1[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i44.GSR = "ENABLED";
    FD1S3AX d1_i45 (.D(d1_71__N_418[45]), .CK(osc_clk), .Q(d1[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i45.GSR = "ENABLED";
    FD1S3AX d1_i46 (.D(d1_71__N_418[46]), .CK(osc_clk), .Q(d1[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i46.GSR = "ENABLED";
    FD1S3AX d1_i47 (.D(d1_71__N_418[47]), .CK(osc_clk), .Q(d1[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i47.GSR = "ENABLED";
    FD1S3AX d1_i48 (.D(d1_71__N_418[48]), .CK(osc_clk), .Q(d1[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i48.GSR = "ENABLED";
    FD1S3AX d1_i49 (.D(d1_71__N_418[49]), .CK(osc_clk), .Q(d1[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i49.GSR = "ENABLED";
    FD1S3AX d1_i50 (.D(d1_71__N_418[50]), .CK(osc_clk), .Q(d1[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i50.GSR = "ENABLED";
    FD1S3AX d1_i51 (.D(d1_71__N_418[51]), .CK(osc_clk), .Q(d1[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i51.GSR = "ENABLED";
    FD1S3AX d1_i52 (.D(d1_71__N_418[52]), .CK(osc_clk), .Q(d1[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i52.GSR = "ENABLED";
    FD1S3AX d1_i53 (.D(d1_71__N_418[53]), .CK(osc_clk), .Q(d1[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i53.GSR = "ENABLED";
    FD1S3AX d1_i54 (.D(d1_71__N_418[54]), .CK(osc_clk), .Q(d1[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i54.GSR = "ENABLED";
    FD1S3AX d1_i55 (.D(d1_71__N_418[55]), .CK(osc_clk), .Q(d1[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i55.GSR = "ENABLED";
    FD1S3AX d1_i56 (.D(d1_71__N_418[56]), .CK(osc_clk), .Q(d1[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i56.GSR = "ENABLED";
    FD1S3AX d1_i57 (.D(d1_71__N_418[57]), .CK(osc_clk), .Q(d1[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i57.GSR = "ENABLED";
    FD1S3AX d1_i58 (.D(d1_71__N_418[58]), .CK(osc_clk), .Q(d1[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i58.GSR = "ENABLED";
    FD1S3AX d1_i59 (.D(d1_71__N_418[59]), .CK(osc_clk), .Q(d1[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i59.GSR = "ENABLED";
    FD1S3AX d1_i60 (.D(d1_71__N_418[60]), .CK(osc_clk), .Q(d1[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i60.GSR = "ENABLED";
    FD1S3AX d1_i61 (.D(d1_71__N_418[61]), .CK(osc_clk), .Q(d1[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i61.GSR = "ENABLED";
    FD1S3AX d1_i62 (.D(d1_71__N_418[62]), .CK(osc_clk), .Q(d1[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i62.GSR = "ENABLED";
    FD1S3AX d1_i63 (.D(d1_71__N_418[63]), .CK(osc_clk), .Q(d1[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i63.GSR = "ENABLED";
    FD1S3AX d1_i64 (.D(d1_71__N_418[64]), .CK(osc_clk), .Q(d1[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i64.GSR = "ENABLED";
    FD1S3AX d1_i65 (.D(d1_71__N_418[65]), .CK(osc_clk), .Q(d1[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i65.GSR = "ENABLED";
    FD1S3AX d1_i66 (.D(d1_71__N_418[66]), .CK(osc_clk), .Q(d1[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i66.GSR = "ENABLED";
    FD1S3AX d1_i67 (.D(d1_71__N_418[67]), .CK(osc_clk), .Q(d1[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i67.GSR = "ENABLED";
    FD1S3AX d1_i68 (.D(d1_71__N_418[68]), .CK(osc_clk), .Q(d1[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i68.GSR = "ENABLED";
    FD1S3AX d1_i69 (.D(d1_71__N_418[69]), .CK(osc_clk), .Q(d1[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i69.GSR = "ENABLED";
    FD1S3AX d1_i70 (.D(d1_71__N_418[70]), .CK(osc_clk), .Q(d1[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i70.GSR = "ENABLED";
    FD1S3AX d1_i71 (.D(d1_71__N_418[71]), .CK(osc_clk), .Q(d1[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i71.GSR = "ENABLED";
    CCU2D add_1057_37 (.A0(d2[70]), .B0(n4451), .C0(n4452[34]), .D0(d1[70]), 
          .A1(d2[71]), .B1(n4451), .C1(n4452[35]), .D1(d1[71]), .CIN(n11936), 
          .S0(d2_71__N_490[70]), .S1(d2_71__N_490[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1057_37.INIT0 = 16'h74b8;
    defparam add_1057_37.INIT1 = 16'h74b8;
    defparam add_1057_37.INJECT1_0 = "NO";
    defparam add_1057_37.INJECT1_1 = "NO";
    CCU2D add_1057_35 (.A0(d2[68]), .B0(n4451), .C0(n4452[32]), .D0(d1[68]), 
          .A1(d2[69]), .B1(n4451), .C1(n4452[33]), .D1(d1[69]), .CIN(n11935), 
          .COUT(n11936), .S0(d2_71__N_490[68]), .S1(d2_71__N_490[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1057_35.INIT0 = 16'h74b8;
    defparam add_1057_35.INIT1 = 16'h74b8;
    defparam add_1057_35.INJECT1_0 = "NO";
    defparam add_1057_35.INJECT1_1 = "NO";
    CCU2D add_1057_33 (.A0(d2[66]), .B0(n4451), .C0(n4452[30]), .D0(d1[66]), 
          .A1(d2[67]), .B1(n4451), .C1(n4452[31]), .D1(d1[67]), .CIN(n11934), 
          .COUT(n11935), .S0(d2_71__N_490[66]), .S1(d2_71__N_490[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1057_33.INIT0 = 16'h74b8;
    defparam add_1057_33.INIT1 = 16'h74b8;
    defparam add_1057_33.INJECT1_0 = "NO";
    defparam add_1057_33.INJECT1_1 = "NO";
    CCU2D add_1057_31 (.A0(d2[64]), .B0(n4451), .C0(n4452[28]), .D0(d1[64]), 
          .A1(d2[65]), .B1(n4451), .C1(n4452[29]), .D1(d1[65]), .CIN(n11933), 
          .COUT(n11934), .S0(d2_71__N_490[64]), .S1(d2_71__N_490[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1057_31.INIT0 = 16'h74b8;
    defparam add_1057_31.INIT1 = 16'h74b8;
    defparam add_1057_31.INJECT1_0 = "NO";
    defparam add_1057_31.INJECT1_1 = "NO";
    CCU2D add_1057_29 (.A0(d2[62]), .B0(n4451), .C0(n4452[26]), .D0(d1[62]), 
          .A1(d2[63]), .B1(n4451), .C1(n4452[27]), .D1(d1[63]), .CIN(n11932), 
          .COUT(n11933), .S0(d2_71__N_490[62]), .S1(d2_71__N_490[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1057_29.INIT0 = 16'h74b8;
    defparam add_1057_29.INIT1 = 16'h74b8;
    defparam add_1057_29.INJECT1_0 = "NO";
    defparam add_1057_29.INJECT1_1 = "NO";
    CCU2D add_1057_27 (.A0(d2[60]), .B0(n4451), .C0(n4452[24]), .D0(d1[60]), 
          .A1(d2[61]), .B1(n4451), .C1(n4452[25]), .D1(d1[61]), .CIN(n11931), 
          .COUT(n11932), .S0(d2_71__N_490[60]), .S1(d2_71__N_490[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1057_27.INIT0 = 16'h74b8;
    defparam add_1057_27.INIT1 = 16'h74b8;
    defparam add_1057_27.INJECT1_0 = "NO";
    defparam add_1057_27.INJECT1_1 = "NO";
    CCU2D add_1057_25 (.A0(d2[58]), .B0(n4451), .C0(n4452[22]), .D0(d1[58]), 
          .A1(d2[59]), .B1(n4451), .C1(n4452[23]), .D1(d1[59]), .CIN(n11930), 
          .COUT(n11931), .S0(d2_71__N_490[58]), .S1(d2_71__N_490[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1057_25.INIT0 = 16'h74b8;
    defparam add_1057_25.INIT1 = 16'h74b8;
    defparam add_1057_25.INJECT1_0 = "NO";
    defparam add_1057_25.INJECT1_1 = "NO";
    CCU2D add_1057_23 (.A0(d2[56]), .B0(n4451), .C0(n4452[20]), .D0(d1[56]), 
          .A1(d2[57]), .B1(n4451), .C1(n4452[21]), .D1(d1[57]), .CIN(n11929), 
          .COUT(n11930), .S0(d2_71__N_490[56]), .S1(d2_71__N_490[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1057_23.INIT0 = 16'h74b8;
    defparam add_1057_23.INIT1 = 16'h74b8;
    defparam add_1057_23.INJECT1_0 = "NO";
    defparam add_1057_23.INJECT1_1 = "NO";
    CCU2D add_1057_21 (.A0(d2[54]), .B0(n4451), .C0(n4452[18]), .D0(d1[54]), 
          .A1(d2[55]), .B1(n4451), .C1(n4452[19]), .D1(d1[55]), .CIN(n11928), 
          .COUT(n11929), .S0(d2_71__N_490[54]), .S1(d2_71__N_490[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1057_21.INIT0 = 16'h74b8;
    defparam add_1057_21.INIT1 = 16'h74b8;
    defparam add_1057_21.INJECT1_0 = "NO";
    defparam add_1057_21.INJECT1_1 = "NO";
    CCU2D add_1057_19 (.A0(d2[52]), .B0(n4451), .C0(n4452[16]), .D0(d1[52]), 
          .A1(d2[53]), .B1(n4451), .C1(n4452[17]), .D1(d1[53]), .CIN(n11927), 
          .COUT(n11928), .S0(d2_71__N_490[52]), .S1(d2_71__N_490[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1057_19.INIT0 = 16'h74b8;
    defparam add_1057_19.INIT1 = 16'h74b8;
    defparam add_1057_19.INJECT1_0 = "NO";
    defparam add_1057_19.INJECT1_1 = "NO";
    CCU2D add_1057_17 (.A0(d2[50]), .B0(n4451), .C0(n4452[14]), .D0(d1[50]), 
          .A1(d2[51]), .B1(n4451), .C1(n4452[15]), .D1(d1[51]), .CIN(n11926), 
          .COUT(n11927), .S0(d2_71__N_490[50]), .S1(d2_71__N_490[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1057_17.INIT0 = 16'h74b8;
    defparam add_1057_17.INIT1 = 16'h74b8;
    defparam add_1057_17.INJECT1_0 = "NO";
    defparam add_1057_17.INJECT1_1 = "NO";
    CCU2D add_1057_15 (.A0(d2[48]), .B0(n4451), .C0(n4452[12]), .D0(d1[48]), 
          .A1(d2[49]), .B1(n4451), .C1(n4452[13]), .D1(d1[49]), .CIN(n11925), 
          .COUT(n11926), .S0(d2_71__N_490[48]), .S1(d2_71__N_490[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1057_15.INIT0 = 16'h74b8;
    defparam add_1057_15.INIT1 = 16'h74b8;
    defparam add_1057_15.INJECT1_0 = "NO";
    defparam add_1057_15.INJECT1_1 = "NO";
    CCU2D add_1057_13 (.A0(d2[46]), .B0(n4451), .C0(n4452[10]), .D0(d1[46]), 
          .A1(d2[47]), .B1(n4451), .C1(n4452[11]), .D1(d1[47]), .CIN(n11924), 
          .COUT(n11925), .S0(d2_71__N_490[46]), .S1(d2_71__N_490[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1057_13.INIT0 = 16'h74b8;
    defparam add_1057_13.INIT1 = 16'h74b8;
    defparam add_1057_13.INJECT1_0 = "NO";
    defparam add_1057_13.INJECT1_1 = "NO";
    CCU2D add_1057_11 (.A0(d2[44]), .B0(n4451), .C0(n4452[8]), .D0(d1[44]), 
          .A1(d2[45]), .B1(n4451), .C1(n4452[9]), .D1(d1[45]), .CIN(n11923), 
          .COUT(n11924), .S0(d2_71__N_490[44]), .S1(d2_71__N_490[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1057_11.INIT0 = 16'h74b8;
    defparam add_1057_11.INIT1 = 16'h74b8;
    defparam add_1057_11.INJECT1_0 = "NO";
    defparam add_1057_11.INJECT1_1 = "NO";
    FD1S3IX count__i2 (.D(n375[2]), .CK(osc_clk), .CD(n8425), .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n375[3]), .CK(osc_clk), .CD(n8425), .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n375[4]), .CK(osc_clk), .CD(n8425), .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n375[5]), .CK(osc_clk), .CD(n8425), .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n375[6]), .CK(osc_clk), .CD(n8425), .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n375[7]), .CK(osc_clk), .CD(n8425), .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n375[8]), .CK(osc_clk), .CD(n8425), .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n375[9]), .CK(osc_clk), .CD(n8425), .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n375[10]), .CK(osc_clk), .CD(n8425), .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_15__N_1442[11]), .CK(osc_clk), .CD(d_clk_tmp_N_1831), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(n375[12]), .CK(osc_clk), .CD(n8425), .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(n375[13]), .CK(osc_clk), .CD(n8425), .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(n375[14]), .CK(osc_clk), .CD(n8425), .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(n375[15]), .CK(osc_clk), .CD(n8425), .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i15.GSR = "ENABLED";
    CCU2D add_1057_9 (.A0(d2[42]), .B0(n4451), .C0(n4452[6]), .D0(d1[42]), 
          .A1(d2[43]), .B1(n4451), .C1(n4452[7]), .D1(d1[43]), .CIN(n11922), 
          .COUT(n11923), .S0(d2_71__N_490[42]), .S1(d2_71__N_490[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1057_9.INIT0 = 16'h74b8;
    defparam add_1057_9.INIT1 = 16'h74b8;
    defparam add_1057_9.INJECT1_0 = "NO";
    defparam add_1057_9.INJECT1_1 = "NO";
    LUT4 i7_2_lut_3_lut (.A(count[13]), .B(count[15]), .C(count[3]), .Z(n21_adj_2495)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i7_2_lut_3_lut.init = 16'h1010;
    CCU2D add_1106_15 (.A0(d9[49]), .B0(d_d9[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[50]), .B1(d_d9[50]), .C1(GND_net), .D1(GND_net), .CIN(n11536), 
          .COUT(n11537));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1106_15.INIT0 = 16'h5999;
    defparam add_1106_15.INIT1 = 16'h5999;
    defparam add_1106_15.INJECT1_0 = "NO";
    defparam add_1106_15.INJECT1_1 = "NO";
    CCU2D add_1057_7 (.A0(d2[40]), .B0(n4451), .C0(n4452[4]), .D0(d1[40]), 
          .A1(d2[41]), .B1(n4451), .C1(n4452[5]), .D1(d1[41]), .CIN(n11921), 
          .COUT(n11922), .S0(d2_71__N_490[40]), .S1(d2_71__N_490[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1057_7.INIT0 = 16'h74b8;
    defparam add_1057_7.INIT1 = 16'h74b8;
    defparam add_1057_7.INJECT1_0 = "NO";
    defparam add_1057_7.INJECT1_1 = "NO";
    CCU2D add_1057_5 (.A0(d2[38]), .B0(n4451), .C0(n4452[2]), .D0(d1[38]), 
          .A1(d2[39]), .B1(n4451), .C1(n4452[3]), .D1(d1[39]), .CIN(n11920), 
          .COUT(n11921), .S0(d2_71__N_490[38]), .S1(d2_71__N_490[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1057_5.INIT0 = 16'h74b8;
    defparam add_1057_5.INIT1 = 16'h74b8;
    defparam add_1057_5.INJECT1_0 = "NO";
    defparam add_1057_5.INJECT1_1 = "NO";
    CCU2D add_1057_3 (.A0(d2[36]), .B0(n4451), .C0(n4452[0]), .D0(d1[36]), 
          .A1(d2[37]), .B1(n4451), .C1(n4452[1]), .D1(d1[37]), .CIN(n11919), 
          .COUT(n11920), .S0(d2_71__N_490[36]), .S1(d2_71__N_490[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1057_3.INIT0 = 16'h74b8;
    defparam add_1057_3.INIT1 = 16'h74b8;
    defparam add_1057_3.INJECT1_0 = "NO";
    defparam add_1057_3.INJECT1_1 = "NO";
    CCU2D add_1057_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n4451), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11919));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1057_1.INIT0 = 16'hF000;
    defparam add_1057_1.INIT1 = 16'h0555;
    defparam add_1057_1.INJECT1_0 = "NO";
    defparam add_1057_1.INJECT1_1 = "NO";
    CCU2D add_1061_36 (.A0(d2[70]), .B0(d3[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[71]), .B1(d3[71]), .C1(GND_net), .D1(GND_net), .CIN(n11914), 
          .S0(n4604[34]), .S1(n4604[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1061_36.INIT0 = 16'h5666;
    defparam add_1061_36.INIT1 = 16'h5666;
    defparam add_1061_36.INJECT1_0 = "NO";
    defparam add_1061_36.INJECT1_1 = "NO";
    CCU2D add_1061_34 (.A0(d2[68]), .B0(d3[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[69]), .B1(d3[69]), .C1(GND_net), .D1(GND_net), .CIN(n11913), 
          .COUT(n11914), .S0(n4604[32]), .S1(n4604[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1061_34.INIT0 = 16'h5666;
    defparam add_1061_34.INIT1 = 16'h5666;
    defparam add_1061_34.INJECT1_0 = "NO";
    defparam add_1061_34.INJECT1_1 = "NO";
    CCU2D add_1061_32 (.A0(d2[66]), .B0(d3[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[67]), .B1(d3[67]), .C1(GND_net), .D1(GND_net), .CIN(n11912), 
          .COUT(n11913), .S0(n4604[30]), .S1(n4604[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1061_32.INIT0 = 16'h5666;
    defparam add_1061_32.INIT1 = 16'h5666;
    defparam add_1061_32.INJECT1_0 = "NO";
    defparam add_1061_32.INJECT1_1 = "NO";
    CCU2D add_1061_30 (.A0(d2[64]), .B0(d3[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[65]), .B1(d3[65]), .C1(GND_net), .D1(GND_net), .CIN(n11911), 
          .COUT(n11912), .S0(n4604[28]), .S1(n4604[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1061_30.INIT0 = 16'h5666;
    defparam add_1061_30.INIT1 = 16'h5666;
    defparam add_1061_30.INJECT1_0 = "NO";
    defparam add_1061_30.INJECT1_1 = "NO";
    LUT4 i75_2_lut_rep_96 (.A(count[12]), .B(count[14]), .Z(n13070)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i75_2_lut_rep_96.init = 16'heeee;
    CCU2D add_1106_13 (.A0(d9[47]), .B0(d_d9[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[48]), .B1(d_d9[48]), .C1(GND_net), .D1(GND_net), .CIN(n11535), 
          .COUT(n11536));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1106_13.INIT0 = 16'h5999;
    defparam add_1106_13.INIT1 = 16'h5999;
    defparam add_1106_13.INJECT1_0 = "NO";
    defparam add_1106_13.INJECT1_1 = "NO";
    CCU2D add_1061_28 (.A0(d2[62]), .B0(d3[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[63]), .B1(d3[63]), .C1(GND_net), .D1(GND_net), .CIN(n11910), 
          .COUT(n11911), .S0(n4604[26]), .S1(n4604[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1061_28.INIT0 = 16'h5666;
    defparam add_1061_28.INIT1 = 16'h5666;
    defparam add_1061_28.INJECT1_0 = "NO";
    defparam add_1061_28.INJECT1_1 = "NO";
    CCU2D add_1106_11 (.A0(d9[45]), .B0(d_d9[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[46]), .B1(d_d9[46]), .C1(GND_net), .D1(GND_net), .CIN(n11534), 
          .COUT(n11535));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1106_11.INIT0 = 16'h5999;
    defparam add_1106_11.INIT1 = 16'h5999;
    defparam add_1106_11.INJECT1_0 = "NO";
    defparam add_1106_11.INJECT1_1 = "NO";
    CCU2D add_1061_26 (.A0(d2[60]), .B0(d3[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[61]), .B1(d3[61]), .C1(GND_net), .D1(GND_net), .CIN(n11909), 
          .COUT(n11910), .S0(n4604[24]), .S1(n4604[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1061_26.INIT0 = 16'h5666;
    defparam add_1061_26.INIT1 = 16'h5666;
    defparam add_1061_26.INJECT1_0 = "NO";
    defparam add_1061_26.INJECT1_1 = "NO";
    CCU2D add_1061_24 (.A0(d2[58]), .B0(d3[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[59]), .B1(d3[59]), .C1(GND_net), .D1(GND_net), .CIN(n11908), 
          .COUT(n11909), .S0(n4604[22]), .S1(n4604[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1061_24.INIT0 = 16'h5666;
    defparam add_1061_24.INIT1 = 16'h5666;
    defparam add_1061_24.INJECT1_0 = "NO";
    defparam add_1061_24.INJECT1_1 = "NO";
    LUT4 i4646_2_lut (.A(d4[36]), .B(d5[36]), .Z(n4908[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4646_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_3_lut (.A(count[12]), .B(count[14]), .C(count[2]), .Z(n15)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h1010;
    CCU2D add_1136_37 (.A0(d7[71]), .B0(d_d7[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11134), 
          .S0(n6884[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1136_37.INIT0 = 16'h5999;
    defparam add_1136_37.INIT1 = 16'h0000;
    defparam add_1136_37.INJECT1_0 = "NO";
    defparam add_1136_37.INJECT1_1 = "NO";
    CCU2D add_1136_35 (.A0(d7[69]), .B0(d_d7[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[70]), .B1(d_d7[70]), .C1(GND_net), .D1(GND_net), .CIN(n11133), 
          .COUT(n11134), .S0(n6884[33]), .S1(n6884[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1136_35.INIT0 = 16'h5999;
    defparam add_1136_35.INIT1 = 16'h5999;
    defparam add_1136_35.INJECT1_0 = "NO";
    defparam add_1136_35.INJECT1_1 = "NO";
    CCU2D add_1136_33 (.A0(d7[67]), .B0(d_d7[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[68]), .B1(d_d7[68]), .C1(GND_net), .D1(GND_net), .CIN(n11132), 
          .COUT(n11133), .S0(n6884[31]), .S1(n6884[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1136_33.INIT0 = 16'h5999;
    defparam add_1136_33.INIT1 = 16'h5999;
    defparam add_1136_33.INJECT1_0 = "NO";
    defparam add_1136_33.INJECT1_1 = "NO";
    CCU2D add_1136_31 (.A0(d7[65]), .B0(d_d7[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[66]), .B1(d_d7[66]), .C1(GND_net), .D1(GND_net), .CIN(n11131), 
          .COUT(n11132), .S0(n6884[29]), .S1(n6884[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1136_31.INIT0 = 16'h5999;
    defparam add_1136_31.INIT1 = 16'h5999;
    defparam add_1136_31.INJECT1_0 = "NO";
    defparam add_1136_31.INJECT1_1 = "NO";
    CCU2D add_1136_29 (.A0(d7[63]), .B0(d_d7[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[64]), .B1(d_d7[64]), .C1(GND_net), .D1(GND_net), .CIN(n11130), 
          .COUT(n11131), .S0(n6884[27]), .S1(n6884[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1136_29.INIT0 = 16'h5999;
    defparam add_1136_29.INIT1 = 16'h5999;
    defparam add_1136_29.INJECT1_0 = "NO";
    defparam add_1136_29.INJECT1_1 = "NO";
    CCU2D add_1136_27 (.A0(d7[61]), .B0(d_d7[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[62]), .B1(d_d7[62]), .C1(GND_net), .D1(GND_net), .CIN(n11129), 
          .COUT(n11130), .S0(n6884[25]), .S1(n6884[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1136_27.INIT0 = 16'h5999;
    defparam add_1136_27.INIT1 = 16'h5999;
    defparam add_1136_27.INJECT1_0 = "NO";
    defparam add_1136_27.INJECT1_1 = "NO";
    CCU2D add_1136_25 (.A0(d7[59]), .B0(d_d7[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[60]), .B1(d_d7[60]), .C1(GND_net), .D1(GND_net), .CIN(n11128), 
          .COUT(n11129), .S0(n6884[23]), .S1(n6884[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1136_25.INIT0 = 16'h5999;
    defparam add_1136_25.INIT1 = 16'h5999;
    defparam add_1136_25.INJECT1_0 = "NO";
    defparam add_1136_25.INJECT1_1 = "NO";
    CCU2D add_1136_23 (.A0(d7[57]), .B0(d_d7[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[58]), .B1(d_d7[58]), .C1(GND_net), .D1(GND_net), .CIN(n11127), 
          .COUT(n11128), .S0(n6884[21]), .S1(n6884[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1136_23.INIT0 = 16'h5999;
    defparam add_1136_23.INIT1 = 16'h5999;
    defparam add_1136_23.INJECT1_0 = "NO";
    defparam add_1136_23.INJECT1_1 = "NO";
    CCU2D add_1136_21 (.A0(d7[55]), .B0(d_d7[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[56]), .B1(d_d7[56]), .C1(GND_net), .D1(GND_net), .CIN(n11126), 
          .COUT(n11127), .S0(n6884[19]), .S1(n6884[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1136_21.INIT0 = 16'h5999;
    defparam add_1136_21.INIT1 = 16'h5999;
    defparam add_1136_21.INJECT1_0 = "NO";
    defparam add_1136_21.INJECT1_1 = "NO";
    CCU2D add_1136_19 (.A0(d7[53]), .B0(d_d7[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[54]), .B1(d_d7[54]), .C1(GND_net), .D1(GND_net), .CIN(n11125), 
          .COUT(n11126), .S0(n6884[17]), .S1(n6884[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1136_19.INIT0 = 16'h5999;
    defparam add_1136_19.INIT1 = 16'h5999;
    defparam add_1136_19.INJECT1_0 = "NO";
    defparam add_1136_19.INJECT1_1 = "NO";
    CCU2D add_1136_17 (.A0(d7[51]), .B0(d_d7[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[52]), .B1(d_d7[52]), .C1(GND_net), .D1(GND_net), .CIN(n11124), 
          .COUT(n11125), .S0(n6884[15]), .S1(n6884[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1136_17.INIT0 = 16'h5999;
    defparam add_1136_17.INIT1 = 16'h5999;
    defparam add_1136_17.INJECT1_0 = "NO";
    defparam add_1136_17.INJECT1_1 = "NO";
    CCU2D add_1136_15 (.A0(d7[49]), .B0(d_d7[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[50]), .B1(d_d7[50]), .C1(GND_net), .D1(GND_net), .CIN(n11123), 
          .COUT(n11124), .S0(n6884[13]), .S1(n6884[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1136_15.INIT0 = 16'h5999;
    defparam add_1136_15.INIT1 = 16'h5999;
    defparam add_1136_15.INJECT1_0 = "NO";
    defparam add_1136_15.INJECT1_1 = "NO";
    CCU2D add_1136_13 (.A0(d7[47]), .B0(d_d7[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[48]), .B1(d_d7[48]), .C1(GND_net), .D1(GND_net), .CIN(n11122), 
          .COUT(n11123), .S0(n6884[11]), .S1(n6884[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1136_13.INIT0 = 16'h5999;
    defparam add_1136_13.INIT1 = 16'h5999;
    defparam add_1136_13.INJECT1_0 = "NO";
    defparam add_1136_13.INJECT1_1 = "NO";
    CCU2D add_1136_11 (.A0(d7[45]), .B0(d_d7[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[46]), .B1(d_d7[46]), .C1(GND_net), .D1(GND_net), .CIN(n11121), 
          .COUT(n11122), .S0(n6884[9]), .S1(n6884[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1136_11.INIT0 = 16'h5999;
    defparam add_1136_11.INIT1 = 16'h5999;
    defparam add_1136_11.INJECT1_0 = "NO";
    defparam add_1136_11.INJECT1_1 = "NO";
    CCU2D add_1136_9 (.A0(d7[43]), .B0(d_d7[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[44]), .B1(d_d7[44]), .C1(GND_net), .D1(GND_net), .CIN(n11120), 
          .COUT(n11121), .S0(n6884[7]), .S1(n6884[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1136_9.INIT0 = 16'h5999;
    defparam add_1136_9.INIT1 = 16'h5999;
    defparam add_1136_9.INJECT1_0 = "NO";
    defparam add_1136_9.INJECT1_1 = "NO";
    CCU2D add_1136_7 (.A0(d7[41]), .B0(d_d7[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[42]), .B1(d_d7[42]), .C1(GND_net), .D1(GND_net), .CIN(n11119), 
          .COUT(n11120), .S0(n6884[5]), .S1(n6884[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1136_7.INIT0 = 16'h5999;
    defparam add_1136_7.INIT1 = 16'h5999;
    defparam add_1136_7.INJECT1_0 = "NO";
    defparam add_1136_7.INJECT1_1 = "NO";
    CCU2D add_1136_5 (.A0(d7[39]), .B0(d_d7[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[40]), .B1(d_d7[40]), .C1(GND_net), .D1(GND_net), .CIN(n11118), 
          .COUT(n11119), .S0(n6884[3]), .S1(n6884[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1136_5.INIT0 = 16'h5999;
    defparam add_1136_5.INIT1 = 16'h5999;
    defparam add_1136_5.INJECT1_0 = "NO";
    defparam add_1136_5.INJECT1_1 = "NO";
    CCU2D add_1136_3 (.A0(d7[37]), .B0(d_d7[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[38]), .B1(d_d7[38]), .C1(GND_net), .D1(GND_net), .CIN(n11117), 
          .COUT(n11118), .S0(n6884[1]), .S1(n6884[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1136_3.INIT0 = 16'h5999;
    defparam add_1136_3.INIT1 = 16'h5999;
    defparam add_1136_3.INJECT1_0 = "NO";
    defparam add_1136_3.INJECT1_1 = "NO";
    CCU2D add_1136_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d7[36]), .B1(d_d7[36]), .C1(GND_net), .D1(GND_net), .COUT(n11117), 
          .S1(n6884[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1136_1.INIT0 = 16'hF000;
    defparam add_1136_1.INIT1 = 16'h5999;
    defparam add_1136_1.INJECT1_0 = "NO";
    defparam add_1136_1.INJECT1_1 = "NO";
    CCU2D add_1137_37 (.A0(d_d7[70]), .B0(n6883), .C0(n6884[34]), .D0(d7[70]), 
          .A1(d_d7[71]), .B1(n6883), .C1(n6884[35]), .D1(d7[71]), .CIN(n11115), 
          .S0(d8_71__N_1603[70]), .S1(d8_71__N_1603[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1137_37.INIT0 = 16'hb874;
    defparam add_1137_37.INIT1 = 16'hb874;
    defparam add_1137_37.INJECT1_0 = "NO";
    defparam add_1137_37.INJECT1_1 = "NO";
    CCU2D add_1137_35 (.A0(d_d7[68]), .B0(n6883), .C0(n6884[32]), .D0(d7[68]), 
          .A1(d_d7[69]), .B1(n6883), .C1(n6884[33]), .D1(d7[69]), .CIN(n11114), 
          .COUT(n11115), .S0(d8_71__N_1603[68]), .S1(d8_71__N_1603[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1137_35.INIT0 = 16'hb874;
    defparam add_1137_35.INIT1 = 16'hb874;
    defparam add_1137_35.INJECT1_0 = "NO";
    defparam add_1137_35.INJECT1_1 = "NO";
    CCU2D add_1137_33 (.A0(d_d7[66]), .B0(n6883), .C0(n6884[30]), .D0(d7[66]), 
          .A1(d_d7[67]), .B1(n6883), .C1(n6884[31]), .D1(d7[67]), .CIN(n11113), 
          .COUT(n11114), .S0(d8_71__N_1603[66]), .S1(d8_71__N_1603[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1137_33.INIT0 = 16'hb874;
    defparam add_1137_33.INIT1 = 16'hb874;
    defparam add_1137_33.INJECT1_0 = "NO";
    defparam add_1137_33.INJECT1_1 = "NO";
    CCU2D add_1137_31 (.A0(d_d7[64]), .B0(n6883), .C0(n6884[28]), .D0(d7[64]), 
          .A1(d_d7[65]), .B1(n6883), .C1(n6884[29]), .D1(d7[65]), .CIN(n11112), 
          .COUT(n11113), .S0(d8_71__N_1603[64]), .S1(d8_71__N_1603[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1137_31.INIT0 = 16'hb874;
    defparam add_1137_31.INIT1 = 16'hb874;
    defparam add_1137_31.INJECT1_0 = "NO";
    defparam add_1137_31.INJECT1_1 = "NO";
    CCU2D add_1137_29 (.A0(d_d7[62]), .B0(n6883), .C0(n6884[26]), .D0(d7[62]), 
          .A1(d_d7[63]), .B1(n6883), .C1(n6884[27]), .D1(d7[63]), .CIN(n11111), 
          .COUT(n11112), .S0(d8_71__N_1603[62]), .S1(d8_71__N_1603[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1137_29.INIT0 = 16'hb874;
    defparam add_1137_29.INIT1 = 16'hb874;
    defparam add_1137_29.INJECT1_0 = "NO";
    defparam add_1137_29.INJECT1_1 = "NO";
    CCU2D add_1137_27 (.A0(d_d7[60]), .B0(n6883), .C0(n6884[24]), .D0(d7[60]), 
          .A1(d_d7[61]), .B1(n6883), .C1(n6884[25]), .D1(d7[61]), .CIN(n11110), 
          .COUT(n11111), .S0(d8_71__N_1603[60]), .S1(d8_71__N_1603[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1137_27.INIT0 = 16'hb874;
    defparam add_1137_27.INIT1 = 16'hb874;
    defparam add_1137_27.INJECT1_0 = "NO";
    defparam add_1137_27.INJECT1_1 = "NO";
    CCU2D add_1137_25 (.A0(d_d7[58]), .B0(n6883), .C0(n6884[22]), .D0(d7[58]), 
          .A1(d_d7[59]), .B1(n6883), .C1(n6884[23]), .D1(d7[59]), .CIN(n11109), 
          .COUT(n11110), .S0(d8_71__N_1603[58]), .S1(d8_71__N_1603[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1137_25.INIT0 = 16'hb874;
    defparam add_1137_25.INIT1 = 16'hb874;
    defparam add_1137_25.INJECT1_0 = "NO";
    defparam add_1137_25.INJECT1_1 = "NO";
    CCU2D add_1137_23 (.A0(d_d7[56]), .B0(n6883), .C0(n6884[20]), .D0(d7[56]), 
          .A1(d_d7[57]), .B1(n6883), .C1(n6884[21]), .D1(d7[57]), .CIN(n11108), 
          .COUT(n11109), .S0(d8_71__N_1603[56]), .S1(d8_71__N_1603[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1137_23.INIT0 = 16'hb874;
    defparam add_1137_23.INIT1 = 16'hb874;
    defparam add_1137_23.INJECT1_0 = "NO";
    defparam add_1137_23.INJECT1_1 = "NO";
    CCU2D add_1137_21 (.A0(d_d7[54]), .B0(n6883), .C0(n6884[18]), .D0(d7[54]), 
          .A1(d_d7[55]), .B1(n6883), .C1(n6884[19]), .D1(d7[55]), .CIN(n11107), 
          .COUT(n11108), .S0(d8_71__N_1603[54]), .S1(d8_71__N_1603[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1137_21.INIT0 = 16'hb874;
    defparam add_1137_21.INIT1 = 16'hb874;
    defparam add_1137_21.INJECT1_0 = "NO";
    defparam add_1137_21.INJECT1_1 = "NO";
    CCU2D add_1137_19 (.A0(d_d7[52]), .B0(n6883), .C0(n6884[16]), .D0(d7[52]), 
          .A1(d_d7[53]), .B1(n6883), .C1(n6884[17]), .D1(d7[53]), .CIN(n11106), 
          .COUT(n11107), .S0(d8_71__N_1603[52]), .S1(d8_71__N_1603[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1137_19.INIT0 = 16'hb874;
    defparam add_1137_19.INIT1 = 16'hb874;
    defparam add_1137_19.INJECT1_0 = "NO";
    defparam add_1137_19.INJECT1_1 = "NO";
    CCU2D add_1137_17 (.A0(d_d7[50]), .B0(n6883), .C0(n6884[14]), .D0(d7[50]), 
          .A1(d_d7[51]), .B1(n6883), .C1(n6884[15]), .D1(d7[51]), .CIN(n11105), 
          .COUT(n11106), .S0(d8_71__N_1603[50]), .S1(d8_71__N_1603[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1137_17.INIT0 = 16'hb874;
    defparam add_1137_17.INIT1 = 16'hb874;
    defparam add_1137_17.INJECT1_0 = "NO";
    defparam add_1137_17.INJECT1_1 = "NO";
    CCU2D add_1137_15 (.A0(d_d7[48]), .B0(n6883), .C0(n6884[12]), .D0(d7[48]), 
          .A1(d_d7[49]), .B1(n6883), .C1(n6884[13]), .D1(d7[49]), .CIN(n11104), 
          .COUT(n11105), .S0(d8_71__N_1603[48]), .S1(d8_71__N_1603[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1137_15.INIT0 = 16'hb874;
    defparam add_1137_15.INIT1 = 16'hb874;
    defparam add_1137_15.INJECT1_0 = "NO";
    defparam add_1137_15.INJECT1_1 = "NO";
    CCU2D add_1137_13 (.A0(d_d7[46]), .B0(n6883), .C0(n6884[10]), .D0(d7[46]), 
          .A1(d_d7[47]), .B1(n6883), .C1(n6884[11]), .D1(d7[47]), .CIN(n11103), 
          .COUT(n11104), .S0(d8_71__N_1603[46]), .S1(d8_71__N_1603[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1137_13.INIT0 = 16'hb874;
    defparam add_1137_13.INIT1 = 16'hb874;
    defparam add_1137_13.INJECT1_0 = "NO";
    defparam add_1137_13.INJECT1_1 = "NO";
    CCU2D add_1137_11 (.A0(d_d7[44]), .B0(n6883), .C0(n6884[8]), .D0(d7[44]), 
          .A1(d_d7[45]), .B1(n6883), .C1(n6884[9]), .D1(d7[45]), .CIN(n11102), 
          .COUT(n11103), .S0(d8_71__N_1603[44]), .S1(d8_71__N_1603[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1137_11.INIT0 = 16'hb874;
    defparam add_1137_11.INIT1 = 16'hb874;
    defparam add_1137_11.INJECT1_0 = "NO";
    defparam add_1137_11.INJECT1_1 = "NO";
    CCU2D add_1137_9 (.A0(d_d7[42]), .B0(n6883), .C0(n6884[6]), .D0(d7[42]), 
          .A1(d_d7[43]), .B1(n6883), .C1(n6884[7]), .D1(d7[43]), .CIN(n11101), 
          .COUT(n11102), .S0(d8_71__N_1603[42]), .S1(d8_71__N_1603[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1137_9.INIT0 = 16'hb874;
    defparam add_1137_9.INIT1 = 16'hb874;
    defparam add_1137_9.INJECT1_0 = "NO";
    defparam add_1137_9.INJECT1_1 = "NO";
    CCU2D add_1137_7 (.A0(d_d7[40]), .B0(n6883), .C0(n6884[4]), .D0(d7[40]), 
          .A1(d_d7[41]), .B1(n6883), .C1(n6884[5]), .D1(d7[41]), .CIN(n11100), 
          .COUT(n11101), .S0(d8_71__N_1603[40]), .S1(d8_71__N_1603[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1137_7.INIT0 = 16'hb874;
    defparam add_1137_7.INIT1 = 16'hb874;
    defparam add_1137_7.INJECT1_0 = "NO";
    defparam add_1137_7.INJECT1_1 = "NO";
    CCU2D add_1137_5 (.A0(d_d7[38]), .B0(n6883), .C0(n6884[2]), .D0(d7[38]), 
          .A1(d_d7[39]), .B1(n6883), .C1(n6884[3]), .D1(d7[39]), .CIN(n11099), 
          .COUT(n11100), .S0(d8_71__N_1603[38]), .S1(d8_71__N_1603[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1137_5.INIT0 = 16'hb874;
    defparam add_1137_5.INIT1 = 16'hb874;
    defparam add_1137_5.INJECT1_0 = "NO";
    defparam add_1137_5.INJECT1_1 = "NO";
    CCU2D add_1137_3 (.A0(d_d7[36]), .B0(n6883), .C0(n6884[0]), .D0(d7[36]), 
          .A1(d_d7[37]), .B1(n6883), .C1(n6884[1]), .D1(d7[37]), .CIN(n11098), 
          .COUT(n11099), .S0(d8_71__N_1603[36]), .S1(d8_71__N_1603[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1137_3.INIT0 = 16'hb874;
    defparam add_1137_3.INIT1 = 16'hb874;
    defparam add_1137_3.INJECT1_0 = "NO";
    defparam add_1137_3.INJECT1_1 = "NO";
    CCU2D add_1137_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n6883), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11098));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1137_1.INIT0 = 16'hF000;
    defparam add_1137_1.INIT1 = 16'h0555;
    defparam add_1137_1.INJECT1_0 = "NO";
    defparam add_1137_1.INJECT1_1 = "NO";
    CCU2D add_1141_37 (.A0(d6[71]), .B0(d_d6[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11094), 
          .S0(n7036[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1141_37.INIT0 = 16'h5999;
    defparam add_1141_37.INIT1 = 16'h0000;
    defparam add_1141_37.INJECT1_0 = "NO";
    defparam add_1141_37.INJECT1_1 = "NO";
    CCU2D add_1141_35 (.A0(d6[69]), .B0(d_d6[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[70]), .B1(d_d6[70]), .C1(GND_net), .D1(GND_net), .CIN(n11093), 
          .COUT(n11094), .S0(n7036[33]), .S1(n7036[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1141_35.INIT0 = 16'h5999;
    defparam add_1141_35.INIT1 = 16'h5999;
    defparam add_1141_35.INJECT1_0 = "NO";
    defparam add_1141_35.INJECT1_1 = "NO";
    CCU2D add_1141_33 (.A0(d6[67]), .B0(d_d6[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[68]), .B1(d_d6[68]), .C1(GND_net), .D1(GND_net), .CIN(n11092), 
          .COUT(n11093), .S0(n7036[31]), .S1(n7036[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1141_33.INIT0 = 16'h5999;
    defparam add_1141_33.INIT1 = 16'h5999;
    defparam add_1141_33.INJECT1_0 = "NO";
    defparam add_1141_33.INJECT1_1 = "NO";
    CCU2D add_1141_31 (.A0(d6[65]), .B0(d_d6[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[66]), .B1(d_d6[66]), .C1(GND_net), .D1(GND_net), .CIN(n11091), 
          .COUT(n11092), .S0(n7036[29]), .S1(n7036[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1141_31.INIT0 = 16'h5999;
    defparam add_1141_31.INIT1 = 16'h5999;
    defparam add_1141_31.INJECT1_0 = "NO";
    defparam add_1141_31.INJECT1_1 = "NO";
    CCU2D add_1141_29 (.A0(d6[63]), .B0(d_d6[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[64]), .B1(d_d6[64]), .C1(GND_net), .D1(GND_net), .CIN(n11090), 
          .COUT(n11091), .S0(n7036[27]), .S1(n7036[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1141_29.INIT0 = 16'h5999;
    defparam add_1141_29.INIT1 = 16'h5999;
    defparam add_1141_29.INJECT1_0 = "NO";
    defparam add_1141_29.INJECT1_1 = "NO";
    CCU2D add_1141_27 (.A0(d6[61]), .B0(d_d6[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[62]), .B1(d_d6[62]), .C1(GND_net), .D1(GND_net), .CIN(n11089), 
          .COUT(n11090), .S0(n7036[25]), .S1(n7036[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1141_27.INIT0 = 16'h5999;
    defparam add_1141_27.INIT1 = 16'h5999;
    defparam add_1141_27.INJECT1_0 = "NO";
    defparam add_1141_27.INJECT1_1 = "NO";
    CCU2D add_1141_25 (.A0(d6[59]), .B0(d_d6[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[60]), .B1(d_d6[60]), .C1(GND_net), .D1(GND_net), .CIN(n11088), 
          .COUT(n11089), .S0(n7036[23]), .S1(n7036[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1141_25.INIT0 = 16'h5999;
    defparam add_1141_25.INIT1 = 16'h5999;
    defparam add_1141_25.INJECT1_0 = "NO";
    defparam add_1141_25.INJECT1_1 = "NO";
    CCU2D add_1141_23 (.A0(d6[57]), .B0(d_d6[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[58]), .B1(d_d6[58]), .C1(GND_net), .D1(GND_net), .CIN(n11087), 
          .COUT(n11088), .S0(n7036[21]), .S1(n7036[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1141_23.INIT0 = 16'h5999;
    defparam add_1141_23.INIT1 = 16'h5999;
    defparam add_1141_23.INJECT1_0 = "NO";
    defparam add_1141_23.INJECT1_1 = "NO";
    CCU2D add_1141_21 (.A0(d6[55]), .B0(d_d6[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[56]), .B1(d_d6[56]), .C1(GND_net), .D1(GND_net), .CIN(n11086), 
          .COUT(n11087), .S0(n7036[19]), .S1(n7036[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1141_21.INIT0 = 16'h5999;
    defparam add_1141_21.INIT1 = 16'h5999;
    defparam add_1141_21.INJECT1_0 = "NO";
    defparam add_1141_21.INJECT1_1 = "NO";
    CCU2D add_1141_19 (.A0(d6[53]), .B0(d_d6[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[54]), .B1(d_d6[54]), .C1(GND_net), .D1(GND_net), .CIN(n11085), 
          .COUT(n11086), .S0(n7036[17]), .S1(n7036[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1141_19.INIT0 = 16'h5999;
    defparam add_1141_19.INIT1 = 16'h5999;
    defparam add_1141_19.INJECT1_0 = "NO";
    defparam add_1141_19.INJECT1_1 = "NO";
    CCU2D add_1141_17 (.A0(d6[51]), .B0(d_d6[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[52]), .B1(d_d6[52]), .C1(GND_net), .D1(GND_net), .CIN(n11084), 
          .COUT(n11085), .S0(n7036[15]), .S1(n7036[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1141_17.INIT0 = 16'h5999;
    defparam add_1141_17.INIT1 = 16'h5999;
    defparam add_1141_17.INJECT1_0 = "NO";
    defparam add_1141_17.INJECT1_1 = "NO";
    CCU2D add_1141_15 (.A0(d6[49]), .B0(d_d6[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[50]), .B1(d_d6[50]), .C1(GND_net), .D1(GND_net), .CIN(n11083), 
          .COUT(n11084), .S0(n7036[13]), .S1(n7036[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1141_15.INIT0 = 16'h5999;
    defparam add_1141_15.INIT1 = 16'h5999;
    defparam add_1141_15.INJECT1_0 = "NO";
    defparam add_1141_15.INJECT1_1 = "NO";
    CCU2D add_1141_13 (.A0(d6[47]), .B0(d_d6[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[48]), .B1(d_d6[48]), .C1(GND_net), .D1(GND_net), .CIN(n11082), 
          .COUT(n11083), .S0(n7036[11]), .S1(n7036[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1141_13.INIT0 = 16'h5999;
    defparam add_1141_13.INIT1 = 16'h5999;
    defparam add_1141_13.INJECT1_0 = "NO";
    defparam add_1141_13.INJECT1_1 = "NO";
    CCU2D add_1141_11 (.A0(d6[45]), .B0(d_d6[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[46]), .B1(d_d6[46]), .C1(GND_net), .D1(GND_net), .CIN(n11081), 
          .COUT(n11082), .S0(n7036[9]), .S1(n7036[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1141_11.INIT0 = 16'h5999;
    defparam add_1141_11.INIT1 = 16'h5999;
    defparam add_1141_11.INJECT1_0 = "NO";
    defparam add_1141_11.INJECT1_1 = "NO";
    CCU2D add_1141_9 (.A0(d6[43]), .B0(d_d6[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[44]), .B1(d_d6[44]), .C1(GND_net), .D1(GND_net), .CIN(n11080), 
          .COUT(n11081), .S0(n7036[7]), .S1(n7036[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1141_9.INIT0 = 16'h5999;
    defparam add_1141_9.INIT1 = 16'h5999;
    defparam add_1141_9.INJECT1_0 = "NO";
    defparam add_1141_9.INJECT1_1 = "NO";
    CCU2D add_1141_7 (.A0(d6[41]), .B0(d_d6[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[42]), .B1(d_d6[42]), .C1(GND_net), .D1(GND_net), .CIN(n11079), 
          .COUT(n11080), .S0(n7036[5]), .S1(n7036[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1141_7.INIT0 = 16'h5999;
    defparam add_1141_7.INIT1 = 16'h5999;
    defparam add_1141_7.INJECT1_0 = "NO";
    defparam add_1141_7.INJECT1_1 = "NO";
    CCU2D add_1141_5 (.A0(d6[39]), .B0(d_d6[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[40]), .B1(d_d6[40]), .C1(GND_net), .D1(GND_net), .CIN(n11078), 
          .COUT(n11079), .S0(n7036[3]), .S1(n7036[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1141_5.INIT0 = 16'h5999;
    defparam add_1141_5.INIT1 = 16'h5999;
    defparam add_1141_5.INJECT1_0 = "NO";
    defparam add_1141_5.INJECT1_1 = "NO";
    CCU2D add_1141_3 (.A0(d6[37]), .B0(d_d6[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[38]), .B1(d_d6[38]), .C1(GND_net), .D1(GND_net), .CIN(n11077), 
          .COUT(n11078), .S0(n7036[1]), .S1(n7036[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1141_3.INIT0 = 16'h5999;
    defparam add_1141_3.INIT1 = 16'h5999;
    defparam add_1141_3.INJECT1_0 = "NO";
    defparam add_1141_3.INJECT1_1 = "NO";
    CCU2D add_1141_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d6[36]), .B1(d_d6[36]), .C1(GND_net), .D1(GND_net), .COUT(n11077), 
          .S1(n7036[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1141_1.INIT0 = 16'hF000;
    defparam add_1141_1.INIT1 = 16'h5999;
    defparam add_1141_1.INJECT1_0 = "NO";
    defparam add_1141_1.INJECT1_1 = "NO";
    CCU2D add_1142_37 (.A0(d_d6[70]), .B0(n7035), .C0(n7036[34]), .D0(d6[70]), 
          .A1(d_d6[71]), .B1(n7035), .C1(n7036[35]), .D1(d6[71]), .CIN(n11075), 
          .S0(d7_71__N_1531[70]), .S1(d7_71__N_1531[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1142_37.INIT0 = 16'hb874;
    defparam add_1142_37.INIT1 = 16'hb874;
    defparam add_1142_37.INJECT1_0 = "NO";
    defparam add_1142_37.INJECT1_1 = "NO";
    CCU2D add_1142_35 (.A0(d_d6[68]), .B0(n7035), .C0(n7036[32]), .D0(d6[68]), 
          .A1(d_d6[69]), .B1(n7035), .C1(n7036[33]), .D1(d6[69]), .CIN(n11074), 
          .COUT(n11075), .S0(d7_71__N_1531[68]), .S1(d7_71__N_1531[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1142_35.INIT0 = 16'hb874;
    defparam add_1142_35.INIT1 = 16'hb874;
    defparam add_1142_35.INJECT1_0 = "NO";
    defparam add_1142_35.INJECT1_1 = "NO";
    CCU2D add_1142_33 (.A0(d_d6[66]), .B0(n7035), .C0(n7036[30]), .D0(d6[66]), 
          .A1(d_d6[67]), .B1(n7035), .C1(n7036[31]), .D1(d6[67]), .CIN(n11073), 
          .COUT(n11074), .S0(d7_71__N_1531[66]), .S1(d7_71__N_1531[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1142_33.INIT0 = 16'hb874;
    defparam add_1142_33.INIT1 = 16'hb874;
    defparam add_1142_33.INJECT1_0 = "NO";
    defparam add_1142_33.INJECT1_1 = "NO";
    CCU2D add_1142_31 (.A0(d_d6[64]), .B0(n7035), .C0(n7036[28]), .D0(d6[64]), 
          .A1(d_d6[65]), .B1(n7035), .C1(n7036[29]), .D1(d6[65]), .CIN(n11072), 
          .COUT(n11073), .S0(d7_71__N_1531[64]), .S1(d7_71__N_1531[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1142_31.INIT0 = 16'hb874;
    defparam add_1142_31.INIT1 = 16'hb874;
    defparam add_1142_31.INJECT1_0 = "NO";
    defparam add_1142_31.INJECT1_1 = "NO";
    CCU2D add_1142_29 (.A0(d_d6[62]), .B0(n7035), .C0(n7036[26]), .D0(d6[62]), 
          .A1(d_d6[63]), .B1(n7035), .C1(n7036[27]), .D1(d6[63]), .CIN(n11071), 
          .COUT(n11072), .S0(d7_71__N_1531[62]), .S1(d7_71__N_1531[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1142_29.INIT0 = 16'hb874;
    defparam add_1142_29.INIT1 = 16'hb874;
    defparam add_1142_29.INJECT1_0 = "NO";
    defparam add_1142_29.INJECT1_1 = "NO";
    CCU2D add_1142_27 (.A0(d_d6[60]), .B0(n7035), .C0(n7036[24]), .D0(d6[60]), 
          .A1(d_d6[61]), .B1(n7035), .C1(n7036[25]), .D1(d6[61]), .CIN(n11070), 
          .COUT(n11071), .S0(d7_71__N_1531[60]), .S1(d7_71__N_1531[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1142_27.INIT0 = 16'hb874;
    defparam add_1142_27.INIT1 = 16'hb874;
    defparam add_1142_27.INJECT1_0 = "NO";
    defparam add_1142_27.INJECT1_1 = "NO";
    CCU2D add_1142_25 (.A0(d_d6[58]), .B0(n7035), .C0(n7036[22]), .D0(d6[58]), 
          .A1(d_d6[59]), .B1(n7035), .C1(n7036[23]), .D1(d6[59]), .CIN(n11069), 
          .COUT(n11070), .S0(d7_71__N_1531[58]), .S1(d7_71__N_1531[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1142_25.INIT0 = 16'hb874;
    defparam add_1142_25.INIT1 = 16'hb874;
    defparam add_1142_25.INJECT1_0 = "NO";
    defparam add_1142_25.INJECT1_1 = "NO";
    CCU2D add_1142_23 (.A0(d_d6[56]), .B0(n7035), .C0(n7036[20]), .D0(d6[56]), 
          .A1(d_d6[57]), .B1(n7035), .C1(n7036[21]), .D1(d6[57]), .CIN(n11068), 
          .COUT(n11069), .S0(d7_71__N_1531[56]), .S1(d7_71__N_1531[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1142_23.INIT0 = 16'hb874;
    defparam add_1142_23.INIT1 = 16'hb874;
    defparam add_1142_23.INJECT1_0 = "NO";
    defparam add_1142_23.INJECT1_1 = "NO";
    CCU2D add_1142_21 (.A0(d_d6[54]), .B0(n7035), .C0(n7036[18]), .D0(d6[54]), 
          .A1(d_d6[55]), .B1(n7035), .C1(n7036[19]), .D1(d6[55]), .CIN(n11067), 
          .COUT(n11068), .S0(d7_71__N_1531[54]), .S1(d7_71__N_1531[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1142_21.INIT0 = 16'hb874;
    defparam add_1142_21.INIT1 = 16'hb874;
    defparam add_1142_21.INJECT1_0 = "NO";
    defparam add_1142_21.INJECT1_1 = "NO";
    CCU2D add_1142_19 (.A0(d_d6[52]), .B0(n7035), .C0(n7036[16]), .D0(d6[52]), 
          .A1(d_d6[53]), .B1(n7035), .C1(n7036[17]), .D1(d6[53]), .CIN(n11066), 
          .COUT(n11067), .S0(d7_71__N_1531[52]), .S1(d7_71__N_1531[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1142_19.INIT0 = 16'hb874;
    defparam add_1142_19.INIT1 = 16'hb874;
    defparam add_1142_19.INJECT1_0 = "NO";
    defparam add_1142_19.INJECT1_1 = "NO";
    CCU2D add_1142_17 (.A0(d_d6[50]), .B0(n7035), .C0(n7036[14]), .D0(d6[50]), 
          .A1(d_d6[51]), .B1(n7035), .C1(n7036[15]), .D1(d6[51]), .CIN(n11065), 
          .COUT(n11066), .S0(d7_71__N_1531[50]), .S1(d7_71__N_1531[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1142_17.INIT0 = 16'hb874;
    defparam add_1142_17.INIT1 = 16'hb874;
    defparam add_1142_17.INJECT1_0 = "NO";
    defparam add_1142_17.INJECT1_1 = "NO";
    CCU2D add_1142_15 (.A0(d_d6[48]), .B0(n7035), .C0(n7036[12]), .D0(d6[48]), 
          .A1(d_d6[49]), .B1(n7035), .C1(n7036[13]), .D1(d6[49]), .CIN(n11064), 
          .COUT(n11065), .S0(d7_71__N_1531[48]), .S1(d7_71__N_1531[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1142_15.INIT0 = 16'hb874;
    defparam add_1142_15.INIT1 = 16'hb874;
    defparam add_1142_15.INJECT1_0 = "NO";
    defparam add_1142_15.INJECT1_1 = "NO";
    CCU2D add_1142_13 (.A0(d_d6[46]), .B0(n7035), .C0(n7036[10]), .D0(d6[46]), 
          .A1(d_d6[47]), .B1(n7035), .C1(n7036[11]), .D1(d6[47]), .CIN(n11063), 
          .COUT(n11064), .S0(d7_71__N_1531[46]), .S1(d7_71__N_1531[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1142_13.INIT0 = 16'hb874;
    defparam add_1142_13.INIT1 = 16'hb874;
    defparam add_1142_13.INJECT1_0 = "NO";
    defparam add_1142_13.INJECT1_1 = "NO";
    CCU2D add_1142_11 (.A0(d_d6[44]), .B0(n7035), .C0(n7036[8]), .D0(d6[44]), 
          .A1(d_d6[45]), .B1(n7035), .C1(n7036[9]), .D1(d6[45]), .CIN(n11062), 
          .COUT(n11063), .S0(d7_71__N_1531[44]), .S1(d7_71__N_1531[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1142_11.INIT0 = 16'hb874;
    defparam add_1142_11.INIT1 = 16'hb874;
    defparam add_1142_11.INJECT1_0 = "NO";
    defparam add_1142_11.INJECT1_1 = "NO";
    CCU2D add_1142_9 (.A0(d_d6[42]), .B0(n7035), .C0(n7036[6]), .D0(d6[42]), 
          .A1(d_d6[43]), .B1(n7035), .C1(n7036[7]), .D1(d6[43]), .CIN(n11061), 
          .COUT(n11062), .S0(d7_71__N_1531[42]), .S1(d7_71__N_1531[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1142_9.INIT0 = 16'hb874;
    defparam add_1142_9.INIT1 = 16'hb874;
    defparam add_1142_9.INJECT1_0 = "NO";
    defparam add_1142_9.INJECT1_1 = "NO";
    CCU2D add_1142_7 (.A0(d_d6[40]), .B0(n7035), .C0(n7036[4]), .D0(d6[40]), 
          .A1(d_d6[41]), .B1(n7035), .C1(n7036[5]), .D1(d6[41]), .CIN(n11060), 
          .COUT(n11061), .S0(d7_71__N_1531[40]), .S1(d7_71__N_1531[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1142_7.INIT0 = 16'hb874;
    defparam add_1142_7.INIT1 = 16'hb874;
    defparam add_1142_7.INJECT1_0 = "NO";
    defparam add_1142_7.INJECT1_1 = "NO";
    CCU2D add_1142_5 (.A0(d_d6[38]), .B0(n7035), .C0(n7036[2]), .D0(d6[38]), 
          .A1(d_d6[39]), .B1(n7035), .C1(n7036[3]), .D1(d6[39]), .CIN(n11059), 
          .COUT(n11060), .S0(d7_71__N_1531[38]), .S1(d7_71__N_1531[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1142_5.INIT0 = 16'hb874;
    defparam add_1142_5.INIT1 = 16'hb874;
    defparam add_1142_5.INJECT1_0 = "NO";
    defparam add_1142_5.INJECT1_1 = "NO";
    CCU2D add_1142_3 (.A0(d_d6[36]), .B0(n7035), .C0(n7036[0]), .D0(d6[36]), 
          .A1(d_d6[37]), .B1(n7035), .C1(n7036[1]), .D1(d6[37]), .CIN(n11058), 
          .COUT(n11059), .S0(d7_71__N_1531[36]), .S1(d7_71__N_1531[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1142_3.INIT0 = 16'hb874;
    defparam add_1142_3.INIT1 = 16'hb874;
    defparam add_1142_3.INJECT1_0 = "NO";
    defparam add_1142_3.INJECT1_1 = "NO";
    CCU2D add_1142_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n7035), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11058));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1142_1.INIT0 = 16'hF000;
    defparam add_1142_1.INIT1 = 16'h0555;
    defparam add_1142_1.INJECT1_0 = "NO";
    defparam add_1142_1.INJECT1_1 = "NO";
    CCU2D add_1045_37 (.A0(d_tmp[35]), .B0(d_d_tmp[35]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n10969), .S0(d6_71__N_1459[35]), .S1(n4147));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1045_37.INIT0 = 16'h5999;
    defparam add_1045_37.INIT1 = 16'h0000;
    defparam add_1045_37.INJECT1_0 = "NO";
    defparam add_1045_37.INJECT1_1 = "NO";
    CCU2D add_1045_35 (.A0(d_tmp[33]), .B0(d_d_tmp[33]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[34]), .B1(d_d_tmp[34]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10968), .COUT(n10969), .S0(d6_71__N_1459[33]), 
          .S1(d6_71__N_1459[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1045_35.INIT0 = 16'h5999;
    defparam add_1045_35.INIT1 = 16'h5999;
    defparam add_1045_35.INJECT1_0 = "NO";
    defparam add_1045_35.INJECT1_1 = "NO";
    CCU2D add_1045_33 (.A0(d_tmp[31]), .B0(d_d_tmp[31]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[32]), .B1(d_d_tmp[32]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10967), .COUT(n10968), .S0(d6_71__N_1459[31]), 
          .S1(d6_71__N_1459[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1045_33.INIT0 = 16'h5999;
    defparam add_1045_33.INIT1 = 16'h5999;
    defparam add_1045_33.INJECT1_0 = "NO";
    defparam add_1045_33.INJECT1_1 = "NO";
    CCU2D add_1045_31 (.A0(d_tmp[29]), .B0(d_d_tmp[29]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[30]), .B1(d_d_tmp[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10966), .COUT(n10967), .S0(d6_71__N_1459[29]), 
          .S1(d6_71__N_1459[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1045_31.INIT0 = 16'h5999;
    defparam add_1045_31.INIT1 = 16'h5999;
    defparam add_1045_31.INJECT1_0 = "NO";
    defparam add_1045_31.INJECT1_1 = "NO";
    CCU2D add_1045_29 (.A0(d_tmp[27]), .B0(d_d_tmp[27]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[28]), .B1(d_d_tmp[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10965), .COUT(n10966), .S0(d6_71__N_1459[27]), 
          .S1(d6_71__N_1459[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1045_29.INIT0 = 16'h5999;
    defparam add_1045_29.INIT1 = 16'h5999;
    defparam add_1045_29.INJECT1_0 = "NO";
    defparam add_1045_29.INJECT1_1 = "NO";
    CCU2D add_1045_27 (.A0(d_tmp[25]), .B0(d_d_tmp[25]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[26]), .B1(d_d_tmp[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10964), .COUT(n10965), .S0(d6_71__N_1459[25]), 
          .S1(d6_71__N_1459[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1045_27.INIT0 = 16'h5999;
    defparam add_1045_27.INIT1 = 16'h5999;
    defparam add_1045_27.INJECT1_0 = "NO";
    defparam add_1045_27.INJECT1_1 = "NO";
    CCU2D add_1045_25 (.A0(d_tmp[23]), .B0(d_d_tmp[23]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[24]), .B1(d_d_tmp[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10963), .COUT(n10964), .S0(d6_71__N_1459[23]), 
          .S1(d6_71__N_1459[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1045_25.INIT0 = 16'h5999;
    defparam add_1045_25.INIT1 = 16'h5999;
    defparam add_1045_25.INJECT1_0 = "NO";
    defparam add_1045_25.INJECT1_1 = "NO";
    CCU2D add_1045_23 (.A0(d_tmp[21]), .B0(d_d_tmp[21]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[22]), .B1(d_d_tmp[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10962), .COUT(n10963), .S0(d6_71__N_1459[21]), 
          .S1(d6_71__N_1459[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1045_23.INIT0 = 16'h5999;
    defparam add_1045_23.INIT1 = 16'h5999;
    defparam add_1045_23.INJECT1_0 = "NO";
    defparam add_1045_23.INJECT1_1 = "NO";
    CCU2D add_1045_21 (.A0(d_tmp[19]), .B0(d_d_tmp[19]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[20]), .B1(d_d_tmp[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10961), .COUT(n10962), .S0(d6_71__N_1459[19]), 
          .S1(d6_71__N_1459[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1045_21.INIT0 = 16'h5999;
    defparam add_1045_21.INIT1 = 16'h5999;
    defparam add_1045_21.INJECT1_0 = "NO";
    defparam add_1045_21.INJECT1_1 = "NO";
    CCU2D add_1045_19 (.A0(d_tmp[17]), .B0(d_d_tmp[17]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[18]), .B1(d_d_tmp[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10960), .COUT(n10961), .S0(d6_71__N_1459[17]), 
          .S1(d6_71__N_1459[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1045_19.INIT0 = 16'h5999;
    defparam add_1045_19.INIT1 = 16'h5999;
    defparam add_1045_19.INJECT1_0 = "NO";
    defparam add_1045_19.INJECT1_1 = "NO";
    CCU2D add_1045_17 (.A0(d_tmp[15]), .B0(d_d_tmp[15]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[16]), .B1(d_d_tmp[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10959), .COUT(n10960), .S0(d6_71__N_1459[15]), 
          .S1(d6_71__N_1459[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1045_17.INIT0 = 16'h5999;
    defparam add_1045_17.INIT1 = 16'h5999;
    defparam add_1045_17.INJECT1_0 = "NO";
    defparam add_1045_17.INJECT1_1 = "NO";
    CCU2D add_1045_15 (.A0(d_tmp[13]), .B0(d_d_tmp[13]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[14]), .B1(d_d_tmp[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10958), .COUT(n10959), .S0(d6_71__N_1459[13]), 
          .S1(d6_71__N_1459[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1045_15.INIT0 = 16'h5999;
    defparam add_1045_15.INIT1 = 16'h5999;
    defparam add_1045_15.INJECT1_0 = "NO";
    defparam add_1045_15.INJECT1_1 = "NO";
    CCU2D add_1045_13 (.A0(d_tmp[11]), .B0(d_d_tmp[11]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[12]), .B1(d_d_tmp[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10957), .COUT(n10958), .S0(d6_71__N_1459[11]), 
          .S1(d6_71__N_1459[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1045_13.INIT0 = 16'h5999;
    defparam add_1045_13.INIT1 = 16'h5999;
    defparam add_1045_13.INJECT1_0 = "NO";
    defparam add_1045_13.INJECT1_1 = "NO";
    CCU2D add_1045_11 (.A0(d_tmp[9]), .B0(d_d_tmp[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[10]), .B1(d_d_tmp[10]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10956), .COUT(n10957), .S0(d6_71__N_1459[9]), .S1(d6_71__N_1459[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1045_11.INIT0 = 16'h5999;
    defparam add_1045_11.INIT1 = 16'h5999;
    defparam add_1045_11.INJECT1_0 = "NO";
    defparam add_1045_11.INJECT1_1 = "NO";
    CCU2D add_1045_9 (.A0(d_tmp[7]), .B0(d_d_tmp[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[8]), .B1(d_d_tmp[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10955), .COUT(n10956), .S0(d6_71__N_1459[7]), .S1(d6_71__N_1459[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1045_9.INIT0 = 16'h5999;
    defparam add_1045_9.INIT1 = 16'h5999;
    defparam add_1045_9.INJECT1_0 = "NO";
    defparam add_1045_9.INJECT1_1 = "NO";
    CCU2D add_1045_7 (.A0(d_tmp[5]), .B0(d_d_tmp[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[6]), .B1(d_d_tmp[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10954), .COUT(n10955), .S0(d6_71__N_1459[5]), .S1(d6_71__N_1459[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1045_7.INIT0 = 16'h5999;
    defparam add_1045_7.INIT1 = 16'h5999;
    defparam add_1045_7.INJECT1_0 = "NO";
    defparam add_1045_7.INJECT1_1 = "NO";
    CCU2D add_1045_5 (.A0(d_tmp[3]), .B0(d_d_tmp[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[4]), .B1(d_d_tmp[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10953), .COUT(n10954), .S0(d6_71__N_1459[3]), .S1(d6_71__N_1459[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1045_5.INIT0 = 16'h5999;
    defparam add_1045_5.INIT1 = 16'h5999;
    defparam add_1045_5.INJECT1_0 = "NO";
    defparam add_1045_5.INJECT1_1 = "NO";
    CCU2D add_1045_3 (.A0(d_tmp[1]), .B0(d_d_tmp[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[2]), .B1(d_d_tmp[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10952), .COUT(n10953), .S0(d6_71__N_1459[1]), .S1(d6_71__N_1459[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1045_3.INIT0 = 16'h5999;
    defparam add_1045_3.INIT1 = 16'h5999;
    defparam add_1045_3.INJECT1_0 = "NO";
    defparam add_1045_3.INJECT1_1 = "NO";
    CCU2D add_1045_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[0]), .B1(d_d_tmp[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n10952), .S1(d6_71__N_1459[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1045_1.INIT0 = 16'h0000;
    defparam add_1045_1.INIT1 = 16'h5999;
    defparam add_1045_1.INJECT1_0 = "NO";
    defparam add_1045_1.INJECT1_1 = "NO";
    CCU2D add_1100_37 (.A0(d8[35]), .B0(d_d8[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10930), 
          .S0(d9_71__N_1675[35]), .S1(n5819));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1100_37.INIT0 = 16'h5999;
    defparam add_1100_37.INIT1 = 16'h0000;
    defparam add_1100_37.INJECT1_0 = "NO";
    defparam add_1100_37.INJECT1_1 = "NO";
    CCU2D add_1100_35 (.A0(d8[33]), .B0(d_d8[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[34]), .B1(d_d8[34]), .C1(GND_net), .D1(GND_net), .CIN(n10929), 
          .COUT(n10930), .S0(d9_71__N_1675[33]), .S1(d9_71__N_1675[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1100_35.INIT0 = 16'h5999;
    defparam add_1100_35.INIT1 = 16'h5999;
    defparam add_1100_35.INJECT1_0 = "NO";
    defparam add_1100_35.INJECT1_1 = "NO";
    CCU2D add_1100_33 (.A0(d8[31]), .B0(d_d8[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[32]), .B1(d_d8[32]), .C1(GND_net), .D1(GND_net), .CIN(n10928), 
          .COUT(n10929), .S0(d9_71__N_1675[31]), .S1(d9_71__N_1675[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1100_33.INIT0 = 16'h5999;
    defparam add_1100_33.INIT1 = 16'h5999;
    defparam add_1100_33.INJECT1_0 = "NO";
    defparam add_1100_33.INJECT1_1 = "NO";
    CCU2D add_1100_31 (.A0(d8[29]), .B0(d_d8[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[30]), .B1(d_d8[30]), .C1(GND_net), .D1(GND_net), .CIN(n10927), 
          .COUT(n10928), .S0(d9_71__N_1675[29]), .S1(d9_71__N_1675[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1100_31.INIT0 = 16'h5999;
    defparam add_1100_31.INIT1 = 16'h5999;
    defparam add_1100_31.INJECT1_0 = "NO";
    defparam add_1100_31.INJECT1_1 = "NO";
    CCU2D add_1100_29 (.A0(d8[27]), .B0(d_d8[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[28]), .B1(d_d8[28]), .C1(GND_net), .D1(GND_net), .CIN(n10926), 
          .COUT(n10927), .S0(d9_71__N_1675[27]), .S1(d9_71__N_1675[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1100_29.INIT0 = 16'h5999;
    defparam add_1100_29.INIT1 = 16'h5999;
    defparam add_1100_29.INJECT1_0 = "NO";
    defparam add_1100_29.INJECT1_1 = "NO";
    CCU2D add_1100_27 (.A0(d8[25]), .B0(d_d8[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[26]), .B1(d_d8[26]), .C1(GND_net), .D1(GND_net), .CIN(n10925), 
          .COUT(n10926), .S0(d9_71__N_1675[25]), .S1(d9_71__N_1675[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1100_27.INIT0 = 16'h5999;
    defparam add_1100_27.INIT1 = 16'h5999;
    defparam add_1100_27.INJECT1_0 = "NO";
    defparam add_1100_27.INJECT1_1 = "NO";
    CCU2D add_1100_25 (.A0(d8[23]), .B0(d_d8[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[24]), .B1(d_d8[24]), .C1(GND_net), .D1(GND_net), .CIN(n10924), 
          .COUT(n10925), .S0(d9_71__N_1675[23]), .S1(d9_71__N_1675[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1100_25.INIT0 = 16'h5999;
    defparam add_1100_25.INIT1 = 16'h5999;
    defparam add_1100_25.INJECT1_0 = "NO";
    defparam add_1100_25.INJECT1_1 = "NO";
    CCU2D add_1100_23 (.A0(d8[21]), .B0(d_d8[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[22]), .B1(d_d8[22]), .C1(GND_net), .D1(GND_net), .CIN(n10923), 
          .COUT(n10924), .S0(d9_71__N_1675[21]), .S1(d9_71__N_1675[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1100_23.INIT0 = 16'h5999;
    defparam add_1100_23.INIT1 = 16'h5999;
    defparam add_1100_23.INJECT1_0 = "NO";
    defparam add_1100_23.INJECT1_1 = "NO";
    CCU2D add_1100_21 (.A0(d8[19]), .B0(d_d8[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[20]), .B1(d_d8[20]), .C1(GND_net), .D1(GND_net), .CIN(n10922), 
          .COUT(n10923), .S0(d9_71__N_1675[19]), .S1(d9_71__N_1675[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1100_21.INIT0 = 16'h5999;
    defparam add_1100_21.INIT1 = 16'h5999;
    defparam add_1100_21.INJECT1_0 = "NO";
    defparam add_1100_21.INJECT1_1 = "NO";
    CCU2D add_1100_19 (.A0(d8[17]), .B0(d_d8[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[18]), .B1(d_d8[18]), .C1(GND_net), .D1(GND_net), .CIN(n10921), 
          .COUT(n10922), .S0(d9_71__N_1675[17]), .S1(d9_71__N_1675[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1100_19.INIT0 = 16'h5999;
    defparam add_1100_19.INIT1 = 16'h5999;
    defparam add_1100_19.INJECT1_0 = "NO";
    defparam add_1100_19.INJECT1_1 = "NO";
    CCU2D add_1100_17 (.A0(d8[15]), .B0(d_d8[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[16]), .B1(d_d8[16]), .C1(GND_net), .D1(GND_net), .CIN(n10920), 
          .COUT(n10921), .S0(d9_71__N_1675[15]), .S1(d9_71__N_1675[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1100_17.INIT0 = 16'h5999;
    defparam add_1100_17.INIT1 = 16'h5999;
    defparam add_1100_17.INJECT1_0 = "NO";
    defparam add_1100_17.INJECT1_1 = "NO";
    CCU2D add_1100_15 (.A0(d8[13]), .B0(d_d8[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[14]), .B1(d_d8[14]), .C1(GND_net), .D1(GND_net), .CIN(n10919), 
          .COUT(n10920), .S0(d9_71__N_1675[13]), .S1(d9_71__N_1675[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1100_15.INIT0 = 16'h5999;
    defparam add_1100_15.INIT1 = 16'h5999;
    defparam add_1100_15.INJECT1_0 = "NO";
    defparam add_1100_15.INJECT1_1 = "NO";
    CCU2D add_1100_13 (.A0(d8[11]), .B0(d_d8[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[12]), .B1(d_d8[12]), .C1(GND_net), .D1(GND_net), .CIN(n10918), 
          .COUT(n10919), .S0(d9_71__N_1675[11]), .S1(d9_71__N_1675[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1100_13.INIT0 = 16'h5999;
    defparam add_1100_13.INIT1 = 16'h5999;
    defparam add_1100_13.INJECT1_0 = "NO";
    defparam add_1100_13.INJECT1_1 = "NO";
    CCU2D add_1100_11 (.A0(d8[9]), .B0(d_d8[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[10]), .B1(d_d8[10]), .C1(GND_net), .D1(GND_net), .CIN(n10917), 
          .COUT(n10918), .S0(d9_71__N_1675[9]), .S1(d9_71__N_1675[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1100_11.INIT0 = 16'h5999;
    defparam add_1100_11.INIT1 = 16'h5999;
    defparam add_1100_11.INJECT1_0 = "NO";
    defparam add_1100_11.INJECT1_1 = "NO";
    CCU2D add_1100_9 (.A0(d8[7]), .B0(d_d8[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[8]), .B1(d_d8[8]), .C1(GND_net), .D1(GND_net), .CIN(n10916), 
          .COUT(n10917), .S0(d9_71__N_1675[7]), .S1(d9_71__N_1675[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1100_9.INIT0 = 16'h5999;
    defparam add_1100_9.INIT1 = 16'h5999;
    defparam add_1100_9.INJECT1_0 = "NO";
    defparam add_1100_9.INJECT1_1 = "NO";
    CCU2D add_1100_7 (.A0(d8[5]), .B0(d_d8[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[6]), .B1(d_d8[6]), .C1(GND_net), .D1(GND_net), .CIN(n10915), 
          .COUT(n10916), .S0(d9_71__N_1675[5]), .S1(d9_71__N_1675[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1100_7.INIT0 = 16'h5999;
    defparam add_1100_7.INIT1 = 16'h5999;
    defparam add_1100_7.INJECT1_0 = "NO";
    defparam add_1100_7.INJECT1_1 = "NO";
    CCU2D add_1100_5 (.A0(d8[3]), .B0(d_d8[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[4]), .B1(d_d8[4]), .C1(GND_net), .D1(GND_net), .CIN(n10914), 
          .COUT(n10915), .S0(d9_71__N_1675[3]), .S1(d9_71__N_1675[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1100_5.INIT0 = 16'h5999;
    defparam add_1100_5.INIT1 = 16'h5999;
    defparam add_1100_5.INJECT1_0 = "NO";
    defparam add_1100_5.INJECT1_1 = "NO";
    CCU2D add_1100_3 (.A0(d8[1]), .B0(d_d8[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[2]), .B1(d_d8[2]), .C1(GND_net), .D1(GND_net), .CIN(n10913), 
          .COUT(n10914), .S0(d9_71__N_1675[1]), .S1(d9_71__N_1675[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1100_3.INIT0 = 16'h5999;
    defparam add_1100_3.INIT1 = 16'h5999;
    defparam add_1100_3.INJECT1_0 = "NO";
    defparam add_1100_3.INJECT1_1 = "NO";
    CCU2D add_1100_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d8[0]), .B1(d_d8[0]), .C1(GND_net), .D1(GND_net), .COUT(n10913), 
          .S1(d9_71__N_1675[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1100_1.INIT0 = 16'h0000;
    defparam add_1100_1.INIT1 = 16'h5999;
    defparam add_1100_1.INJECT1_0 = "NO";
    defparam add_1100_1.INJECT1_1 = "NO";
    CCU2D add_10_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10806), 
          .S0(n375[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_17.INIT0 = 16'h5aaa;
    defparam add_10_17.INIT1 = 16'h0000;
    defparam add_10_17.INJECT1_0 = "NO";
    defparam add_10_17.INJECT1_1 = "NO";
    CCU2D add_10_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n10805), .COUT(n10806), .S0(n375[13]), .S1(n375[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_15.INIT0 = 16'h5aaa;
    defparam add_10_15.INIT1 = 16'h5aaa;
    defparam add_10_15.INJECT1_0 = "NO";
    defparam add_10_15.INJECT1_1 = "NO";
    CCU2D add_10_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n10804), .COUT(n10805), .S0(n375[11]), .S1(n375[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_13.INIT0 = 16'h5aaa;
    defparam add_10_13.INIT1 = 16'h5aaa;
    defparam add_10_13.INJECT1_0 = "NO";
    defparam add_10_13.INJECT1_1 = "NO";
    CCU2D add_10_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n10803), .COUT(n10804), .S0(n375[9]), .S1(n375[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_11.INIT0 = 16'h5aaa;
    defparam add_10_11.INIT1 = 16'h5aaa;
    defparam add_10_11.INJECT1_0 = "NO";
    defparam add_10_11.INJECT1_1 = "NO";
    CCU2D add_10_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10802), 
          .COUT(n10803), .S0(n375[7]), .S1(n375[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_9.INIT0 = 16'h5aaa;
    defparam add_10_9.INIT1 = 16'h5aaa;
    defparam add_10_9.INJECT1_0 = "NO";
    defparam add_10_9.INJECT1_1 = "NO";
    CCU2D add_10_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10801), 
          .COUT(n10802), .S0(n375[5]), .S1(n375[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_7.INIT0 = 16'h5aaa;
    defparam add_10_7.INIT1 = 16'h5aaa;
    defparam add_10_7.INJECT1_0 = "NO";
    defparam add_10_7.INJECT1_1 = "NO";
    CCU2D add_10_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10800), 
          .COUT(n10801), .S0(n375[3]), .S1(n375[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_5.INIT0 = 16'h5aaa;
    defparam add_10_5.INIT1 = 16'h5aaa;
    defparam add_10_5.INJECT1_0 = "NO";
    defparam add_10_5.INJECT1_1 = "NO";
    CCU2D add_10_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10799), 
          .COUT(n10800), .S0(n375[1]), .S1(n375[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_3.INIT0 = 16'h5aaa;
    defparam add_10_3.INIT1 = 16'h5aaa;
    defparam add_10_3.INJECT1_0 = "NO";
    defparam add_10_3.INJECT1_1 = "NO";
    CCU2D add_10_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n10799), 
          .S1(n375[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_1.INIT0 = 16'hF000;
    defparam add_10_1.INIT1 = 16'h5555;
    defparam add_10_1.INJECT1_0 = "NO";
    defparam add_10_1.INJECT1_1 = "NO";
    CCU2D add_1070_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10779), 
          .S0(n4907));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1070_cout.INIT0 = 16'h0000;
    defparam add_1070_cout.INIT1 = 16'h0000;
    defparam add_1070_cout.INJECT1_0 = "NO";
    defparam add_1070_cout.INJECT1_1 = "NO";
    CCU2D add_1070_36 (.A0(d4[34]), .B0(d5[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[35]), .B1(d5[35]), .C1(GND_net), .D1(GND_net), .CIN(n10778), 
          .COUT(n10779), .S0(d5_71__N_706[34]), .S1(d5_71__N_706[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1070_36.INIT0 = 16'h5666;
    defparam add_1070_36.INIT1 = 16'h5666;
    defparam add_1070_36.INJECT1_0 = "NO";
    defparam add_1070_36.INJECT1_1 = "NO";
    CCU2D add_1070_34 (.A0(d4[32]), .B0(d5[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[33]), .B1(d5[33]), .C1(GND_net), .D1(GND_net), .CIN(n10777), 
          .COUT(n10778), .S0(d5_71__N_706[32]), .S1(d5_71__N_706[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1070_34.INIT0 = 16'h5666;
    defparam add_1070_34.INIT1 = 16'h5666;
    defparam add_1070_34.INJECT1_0 = "NO";
    defparam add_1070_34.INJECT1_1 = "NO";
    CCU2D add_1070_32 (.A0(d4[30]), .B0(d5[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[31]), .B1(d5[31]), .C1(GND_net), .D1(GND_net), .CIN(n10776), 
          .COUT(n10777), .S0(d5_71__N_706[30]), .S1(d5_71__N_706[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1070_32.INIT0 = 16'h5666;
    defparam add_1070_32.INIT1 = 16'h5666;
    defparam add_1070_32.INJECT1_0 = "NO";
    defparam add_1070_32.INJECT1_1 = "NO";
    CCU2D add_1070_30 (.A0(d4[28]), .B0(d5[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[29]), .B1(d5[29]), .C1(GND_net), .D1(GND_net), .CIN(n10775), 
          .COUT(n10776), .S0(d5_71__N_706[28]), .S1(d5_71__N_706[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1070_30.INIT0 = 16'h5666;
    defparam add_1070_30.INIT1 = 16'h5666;
    defparam add_1070_30.INJECT1_0 = "NO";
    defparam add_1070_30.INJECT1_1 = "NO";
    CCU2D add_1070_28 (.A0(d4[26]), .B0(d5[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[27]), .B1(d5[27]), .C1(GND_net), .D1(GND_net), .CIN(n10774), 
          .COUT(n10775), .S0(d5_71__N_706[26]), .S1(d5_71__N_706[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1070_28.INIT0 = 16'h5666;
    defparam add_1070_28.INIT1 = 16'h5666;
    defparam add_1070_28.INJECT1_0 = "NO";
    defparam add_1070_28.INJECT1_1 = "NO";
    CCU2D add_1070_26 (.A0(d4[24]), .B0(d5[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[25]), .B1(d5[25]), .C1(GND_net), .D1(GND_net), .CIN(n10773), 
          .COUT(n10774), .S0(d5_71__N_706[24]), .S1(d5_71__N_706[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1070_26.INIT0 = 16'h5666;
    defparam add_1070_26.INIT1 = 16'h5666;
    defparam add_1070_26.INJECT1_0 = "NO";
    defparam add_1070_26.INJECT1_1 = "NO";
    CCU2D add_1070_24 (.A0(d4[22]), .B0(d5[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[23]), .B1(d5[23]), .C1(GND_net), .D1(GND_net), .CIN(n10772), 
          .COUT(n10773), .S0(d5_71__N_706[22]), .S1(d5_71__N_706[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1070_24.INIT0 = 16'h5666;
    defparam add_1070_24.INIT1 = 16'h5666;
    defparam add_1070_24.INJECT1_0 = "NO";
    defparam add_1070_24.INJECT1_1 = "NO";
    CCU2D add_1070_22 (.A0(d4[20]), .B0(d5[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[21]), .B1(d5[21]), .C1(GND_net), .D1(GND_net), .CIN(n10771), 
          .COUT(n10772), .S0(d5_71__N_706[20]), .S1(d5_71__N_706[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1070_22.INIT0 = 16'h5666;
    defparam add_1070_22.INIT1 = 16'h5666;
    defparam add_1070_22.INJECT1_0 = "NO";
    defparam add_1070_22.INJECT1_1 = "NO";
    CCU2D add_1070_20 (.A0(d4[18]), .B0(d5[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[19]), .B1(d5[19]), .C1(GND_net), .D1(GND_net), .CIN(n10770), 
          .COUT(n10771), .S0(d5_71__N_706[18]), .S1(d5_71__N_706[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1070_20.INIT0 = 16'h5666;
    defparam add_1070_20.INIT1 = 16'h5666;
    defparam add_1070_20.INJECT1_0 = "NO";
    defparam add_1070_20.INJECT1_1 = "NO";
    CCU2D add_1070_18 (.A0(d4[16]), .B0(d5[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[17]), .B1(d5[17]), .C1(GND_net), .D1(GND_net), .CIN(n10769), 
          .COUT(n10770), .S0(d5_71__N_706[16]), .S1(d5_71__N_706[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1070_18.INIT0 = 16'h5666;
    defparam add_1070_18.INIT1 = 16'h5666;
    defparam add_1070_18.INJECT1_0 = "NO";
    defparam add_1070_18.INJECT1_1 = "NO";
    CCU2D add_1070_16 (.A0(d4[14]), .B0(d5[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[15]), .B1(d5[15]), .C1(GND_net), .D1(GND_net), .CIN(n10768), 
          .COUT(n10769), .S0(d5_71__N_706[14]), .S1(d5_71__N_706[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1070_16.INIT0 = 16'h5666;
    defparam add_1070_16.INIT1 = 16'h5666;
    defparam add_1070_16.INJECT1_0 = "NO";
    defparam add_1070_16.INJECT1_1 = "NO";
    CCU2D add_1070_14 (.A0(d4[12]), .B0(d5[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[13]), .B1(d5[13]), .C1(GND_net), .D1(GND_net), .CIN(n10767), 
          .COUT(n10768), .S0(d5_71__N_706[12]), .S1(d5_71__N_706[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1070_14.INIT0 = 16'h5666;
    defparam add_1070_14.INIT1 = 16'h5666;
    defparam add_1070_14.INJECT1_0 = "NO";
    defparam add_1070_14.INJECT1_1 = "NO";
    CCU2D add_1070_12 (.A0(d4[10]), .B0(d5[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[11]), .B1(d5[11]), .C1(GND_net), .D1(GND_net), .CIN(n10766), 
          .COUT(n10767), .S0(d5_71__N_706[10]), .S1(d5_71__N_706[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1070_12.INIT0 = 16'h5666;
    defparam add_1070_12.INIT1 = 16'h5666;
    defparam add_1070_12.INJECT1_0 = "NO";
    defparam add_1070_12.INJECT1_1 = "NO";
    CCU2D add_1070_10 (.A0(d4[8]), .B0(d5[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[9]), .B1(d5[9]), .C1(GND_net), .D1(GND_net), .CIN(n10765), 
          .COUT(n10766), .S0(d5_71__N_706[8]), .S1(d5_71__N_706[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1070_10.INIT0 = 16'h5666;
    defparam add_1070_10.INIT1 = 16'h5666;
    defparam add_1070_10.INJECT1_0 = "NO";
    defparam add_1070_10.INJECT1_1 = "NO";
    CCU2D add_1070_8 (.A0(d4[6]), .B0(d5[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[7]), .B1(d5[7]), .C1(GND_net), .D1(GND_net), .CIN(n10764), 
          .COUT(n10765), .S0(d5_71__N_706[6]), .S1(d5_71__N_706[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1070_8.INIT0 = 16'h5666;
    defparam add_1070_8.INIT1 = 16'h5666;
    defparam add_1070_8.INJECT1_0 = "NO";
    defparam add_1070_8.INJECT1_1 = "NO";
    CCU2D add_1070_6 (.A0(d4[4]), .B0(d5[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[5]), .B1(d5[5]), .C1(GND_net), .D1(GND_net), .CIN(n10763), 
          .COUT(n10764), .S0(d5_71__N_706[4]), .S1(d5_71__N_706[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1070_6.INIT0 = 16'h5666;
    defparam add_1070_6.INIT1 = 16'h5666;
    defparam add_1070_6.INJECT1_0 = "NO";
    defparam add_1070_6.INJECT1_1 = "NO";
    CCU2D add_1070_4 (.A0(d4[2]), .B0(d5[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[3]), .B1(d5[3]), .C1(GND_net), .D1(GND_net), .CIN(n10762), 
          .COUT(n10763), .S0(d5_71__N_706[2]), .S1(d5_71__N_706[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1070_4.INIT0 = 16'h5666;
    defparam add_1070_4.INIT1 = 16'h5666;
    defparam add_1070_4.INJECT1_0 = "NO";
    defparam add_1070_4.INJECT1_1 = "NO";
    CCU2D add_1070_2 (.A0(d4[0]), .B0(d5[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[1]), .B1(d5[1]), .C1(GND_net), .D1(GND_net), .COUT(n10762), 
          .S1(d5_71__N_706[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1070_2.INIT0 = 16'h7000;
    defparam add_1070_2.INIT1 = 16'h5666;
    defparam add_1070_2.INJECT1_0 = "NO";
    defparam add_1070_2.INJECT1_1 = "NO";
    CCU2D add_1065_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10760), 
          .S0(n4755));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1065_cout.INIT0 = 16'h0000;
    defparam add_1065_cout.INIT1 = 16'h0000;
    defparam add_1065_cout.INJECT1_0 = "NO";
    defparam add_1065_cout.INJECT1_1 = "NO";
    CCU2D add_1065_36 (.A0(d3[34]), .B0(d4[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[35]), .B1(d4[35]), .C1(GND_net), .D1(GND_net), .CIN(n10759), 
          .COUT(n10760), .S0(d4_71__N_634[34]), .S1(d4_71__N_634[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1065_36.INIT0 = 16'h5666;
    defparam add_1065_36.INIT1 = 16'h5666;
    defparam add_1065_36.INJECT1_0 = "NO";
    defparam add_1065_36.INJECT1_1 = "NO";
    CCU2D add_1065_34 (.A0(d3[32]), .B0(d4[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[33]), .B1(d4[33]), .C1(GND_net), .D1(GND_net), .CIN(n10758), 
          .COUT(n10759), .S0(d4_71__N_634[32]), .S1(d4_71__N_634[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1065_34.INIT0 = 16'h5666;
    defparam add_1065_34.INIT1 = 16'h5666;
    defparam add_1065_34.INJECT1_0 = "NO";
    defparam add_1065_34.INJECT1_1 = "NO";
    CCU2D add_1065_32 (.A0(d3[30]), .B0(d4[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[31]), .B1(d4[31]), .C1(GND_net), .D1(GND_net), .CIN(n10757), 
          .COUT(n10758), .S0(d4_71__N_634[30]), .S1(d4_71__N_634[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1065_32.INIT0 = 16'h5666;
    defparam add_1065_32.INIT1 = 16'h5666;
    defparam add_1065_32.INJECT1_0 = "NO";
    defparam add_1065_32.INJECT1_1 = "NO";
    CCU2D add_1065_30 (.A0(d3[28]), .B0(d4[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[29]), .B1(d4[29]), .C1(GND_net), .D1(GND_net), .CIN(n10756), 
          .COUT(n10757), .S0(d4_71__N_634[28]), .S1(d4_71__N_634[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1065_30.INIT0 = 16'h5666;
    defparam add_1065_30.INIT1 = 16'h5666;
    defparam add_1065_30.INJECT1_0 = "NO";
    defparam add_1065_30.INJECT1_1 = "NO";
    CCU2D add_1065_28 (.A0(d3[26]), .B0(d4[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[27]), .B1(d4[27]), .C1(GND_net), .D1(GND_net), .CIN(n10755), 
          .COUT(n10756), .S0(d4_71__N_634[26]), .S1(d4_71__N_634[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1065_28.INIT0 = 16'h5666;
    defparam add_1065_28.INIT1 = 16'h5666;
    defparam add_1065_28.INJECT1_0 = "NO";
    defparam add_1065_28.INJECT1_1 = "NO";
    CCU2D add_1065_26 (.A0(d3[24]), .B0(d4[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[25]), .B1(d4[25]), .C1(GND_net), .D1(GND_net), .CIN(n10754), 
          .COUT(n10755), .S0(d4_71__N_634[24]), .S1(d4_71__N_634[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1065_26.INIT0 = 16'h5666;
    defparam add_1065_26.INIT1 = 16'h5666;
    defparam add_1065_26.INJECT1_0 = "NO";
    defparam add_1065_26.INJECT1_1 = "NO";
    CCU2D add_1065_24 (.A0(d3[22]), .B0(d4[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[23]), .B1(d4[23]), .C1(GND_net), .D1(GND_net), .CIN(n10753), 
          .COUT(n10754), .S0(d4_71__N_634[22]), .S1(d4_71__N_634[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1065_24.INIT0 = 16'h5666;
    defparam add_1065_24.INIT1 = 16'h5666;
    defparam add_1065_24.INJECT1_0 = "NO";
    defparam add_1065_24.INJECT1_1 = "NO";
    CCU2D add_1065_22 (.A0(d3[20]), .B0(d4[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[21]), .B1(d4[21]), .C1(GND_net), .D1(GND_net), .CIN(n10752), 
          .COUT(n10753), .S0(d4_71__N_634[20]), .S1(d4_71__N_634[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1065_22.INIT0 = 16'h5666;
    defparam add_1065_22.INIT1 = 16'h5666;
    defparam add_1065_22.INJECT1_0 = "NO";
    defparam add_1065_22.INJECT1_1 = "NO";
    CCU2D add_1065_20 (.A0(d3[18]), .B0(d4[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[19]), .B1(d4[19]), .C1(GND_net), .D1(GND_net), .CIN(n10751), 
          .COUT(n10752), .S0(d4_71__N_634[18]), .S1(d4_71__N_634[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1065_20.INIT0 = 16'h5666;
    defparam add_1065_20.INIT1 = 16'h5666;
    defparam add_1065_20.INJECT1_0 = "NO";
    defparam add_1065_20.INJECT1_1 = "NO";
    CCU2D add_1065_18 (.A0(d3[16]), .B0(d4[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[17]), .B1(d4[17]), .C1(GND_net), .D1(GND_net), .CIN(n10750), 
          .COUT(n10751), .S0(d4_71__N_634[16]), .S1(d4_71__N_634[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1065_18.INIT0 = 16'h5666;
    defparam add_1065_18.INIT1 = 16'h5666;
    defparam add_1065_18.INJECT1_0 = "NO";
    defparam add_1065_18.INJECT1_1 = "NO";
    CCU2D add_1065_16 (.A0(d3[14]), .B0(d4[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[15]), .B1(d4[15]), .C1(GND_net), .D1(GND_net), .CIN(n10749), 
          .COUT(n10750), .S0(d4_71__N_634[14]), .S1(d4_71__N_634[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1065_16.INIT0 = 16'h5666;
    defparam add_1065_16.INIT1 = 16'h5666;
    defparam add_1065_16.INJECT1_0 = "NO";
    defparam add_1065_16.INJECT1_1 = "NO";
    CCU2D add_1065_14 (.A0(d3[12]), .B0(d4[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[13]), .B1(d4[13]), .C1(GND_net), .D1(GND_net), .CIN(n10748), 
          .COUT(n10749), .S0(d4_71__N_634[12]), .S1(d4_71__N_634[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1065_14.INIT0 = 16'h5666;
    defparam add_1065_14.INIT1 = 16'h5666;
    defparam add_1065_14.INJECT1_0 = "NO";
    defparam add_1065_14.INJECT1_1 = "NO";
    CCU2D add_1065_12 (.A0(d3[10]), .B0(d4[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[11]), .B1(d4[11]), .C1(GND_net), .D1(GND_net), .CIN(n10747), 
          .COUT(n10748), .S0(d4_71__N_634[10]), .S1(d4_71__N_634[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1065_12.INIT0 = 16'h5666;
    defparam add_1065_12.INIT1 = 16'h5666;
    defparam add_1065_12.INJECT1_0 = "NO";
    defparam add_1065_12.INJECT1_1 = "NO";
    CCU2D add_1065_10 (.A0(d3[8]), .B0(d4[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[9]), .B1(d4[9]), .C1(GND_net), .D1(GND_net), .CIN(n10746), 
          .COUT(n10747), .S0(d4_71__N_634[8]), .S1(d4_71__N_634[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1065_10.INIT0 = 16'h5666;
    defparam add_1065_10.INIT1 = 16'h5666;
    defparam add_1065_10.INJECT1_0 = "NO";
    defparam add_1065_10.INJECT1_1 = "NO";
    CCU2D add_1065_8 (.A0(d3[6]), .B0(d4[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[7]), .B1(d4[7]), .C1(GND_net), .D1(GND_net), .CIN(n10745), 
          .COUT(n10746), .S0(d4_71__N_634[6]), .S1(d4_71__N_634[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1065_8.INIT0 = 16'h5666;
    defparam add_1065_8.INIT1 = 16'h5666;
    defparam add_1065_8.INJECT1_0 = "NO";
    defparam add_1065_8.INJECT1_1 = "NO";
    CCU2D add_1065_6 (.A0(d3[4]), .B0(d4[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[5]), .B1(d4[5]), .C1(GND_net), .D1(GND_net), .CIN(n10744), 
          .COUT(n10745), .S0(d4_71__N_634[4]), .S1(d4_71__N_634[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1065_6.INIT0 = 16'h5666;
    defparam add_1065_6.INIT1 = 16'h5666;
    defparam add_1065_6.INJECT1_0 = "NO";
    defparam add_1065_6.INJECT1_1 = "NO";
    CCU2D add_1065_4 (.A0(d3[2]), .B0(d4[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[3]), .B1(d4[3]), .C1(GND_net), .D1(GND_net), .CIN(n10743), 
          .COUT(n10744), .S0(d4_71__N_634[2]), .S1(d4_71__N_634[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1065_4.INIT0 = 16'h5666;
    defparam add_1065_4.INIT1 = 16'h5666;
    defparam add_1065_4.INJECT1_0 = "NO";
    defparam add_1065_4.INJECT1_1 = "NO";
    CCU2D add_1065_2 (.A0(d3[0]), .B0(d4[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[1]), .B1(d4[1]), .C1(GND_net), .D1(GND_net), .COUT(n10743), 
          .S1(d4_71__N_634[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1065_2.INIT0 = 16'h7000;
    defparam add_1065_2.INIT1 = 16'h5666;
    defparam add_1065_2.INJECT1_0 = "NO";
    defparam add_1065_2.INJECT1_1 = "NO";
    CCU2D add_1060_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10741), 
          .S0(n4603));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1060_cout.INIT0 = 16'h0000;
    defparam add_1060_cout.INIT1 = 16'h0000;
    defparam add_1060_cout.INJECT1_0 = "NO";
    defparam add_1060_cout.INJECT1_1 = "NO";
    CCU2D add_1060_36 (.A0(d2[34]), .B0(d3[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[35]), .B1(d3[35]), .C1(GND_net), .D1(GND_net), .CIN(n10740), 
          .COUT(n10741), .S0(d3_71__N_562[34]), .S1(d3_71__N_562[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1060_36.INIT0 = 16'h5666;
    defparam add_1060_36.INIT1 = 16'h5666;
    defparam add_1060_36.INJECT1_0 = "NO";
    defparam add_1060_36.INJECT1_1 = "NO";
    CCU2D add_1060_34 (.A0(d2[32]), .B0(d3[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[33]), .B1(d3[33]), .C1(GND_net), .D1(GND_net), .CIN(n10739), 
          .COUT(n10740), .S0(d3_71__N_562[32]), .S1(d3_71__N_562[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1060_34.INIT0 = 16'h5666;
    defparam add_1060_34.INIT1 = 16'h5666;
    defparam add_1060_34.INJECT1_0 = "NO";
    defparam add_1060_34.INJECT1_1 = "NO";
    CCU2D add_1060_32 (.A0(d2[30]), .B0(d3[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[31]), .B1(d3[31]), .C1(GND_net), .D1(GND_net), .CIN(n10738), 
          .COUT(n10739), .S0(d3_71__N_562[30]), .S1(d3_71__N_562[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1060_32.INIT0 = 16'h5666;
    defparam add_1060_32.INIT1 = 16'h5666;
    defparam add_1060_32.INJECT1_0 = "NO";
    defparam add_1060_32.INJECT1_1 = "NO";
    CCU2D add_1060_30 (.A0(d2[28]), .B0(d3[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[29]), .B1(d3[29]), .C1(GND_net), .D1(GND_net), .CIN(n10737), 
          .COUT(n10738), .S0(d3_71__N_562[28]), .S1(d3_71__N_562[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1060_30.INIT0 = 16'h5666;
    defparam add_1060_30.INIT1 = 16'h5666;
    defparam add_1060_30.INJECT1_0 = "NO";
    defparam add_1060_30.INJECT1_1 = "NO";
    CCU2D add_1060_28 (.A0(d2[26]), .B0(d3[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[27]), .B1(d3[27]), .C1(GND_net), .D1(GND_net), .CIN(n10736), 
          .COUT(n10737), .S0(d3_71__N_562[26]), .S1(d3_71__N_562[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1060_28.INIT0 = 16'h5666;
    defparam add_1060_28.INIT1 = 16'h5666;
    defparam add_1060_28.INJECT1_0 = "NO";
    defparam add_1060_28.INJECT1_1 = "NO";
    CCU2D add_1060_26 (.A0(d2[24]), .B0(d3[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[25]), .B1(d3[25]), .C1(GND_net), .D1(GND_net), .CIN(n10735), 
          .COUT(n10736), .S0(d3_71__N_562[24]), .S1(d3_71__N_562[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1060_26.INIT0 = 16'h5666;
    defparam add_1060_26.INIT1 = 16'h5666;
    defparam add_1060_26.INJECT1_0 = "NO";
    defparam add_1060_26.INJECT1_1 = "NO";
    CCU2D add_1060_24 (.A0(d2[22]), .B0(d3[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[23]), .B1(d3[23]), .C1(GND_net), .D1(GND_net), .CIN(n10734), 
          .COUT(n10735), .S0(d3_71__N_562[22]), .S1(d3_71__N_562[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1060_24.INIT0 = 16'h5666;
    defparam add_1060_24.INIT1 = 16'h5666;
    defparam add_1060_24.INJECT1_0 = "NO";
    defparam add_1060_24.INJECT1_1 = "NO";
    CCU2D add_1060_22 (.A0(d2[20]), .B0(d3[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[21]), .B1(d3[21]), .C1(GND_net), .D1(GND_net), .CIN(n10733), 
          .COUT(n10734), .S0(d3_71__N_562[20]), .S1(d3_71__N_562[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1060_22.INIT0 = 16'h5666;
    defparam add_1060_22.INIT1 = 16'h5666;
    defparam add_1060_22.INJECT1_0 = "NO";
    defparam add_1060_22.INJECT1_1 = "NO";
    CCU2D add_1060_20 (.A0(d2[18]), .B0(d3[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[19]), .B1(d3[19]), .C1(GND_net), .D1(GND_net), .CIN(n10732), 
          .COUT(n10733), .S0(d3_71__N_562[18]), .S1(d3_71__N_562[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1060_20.INIT0 = 16'h5666;
    defparam add_1060_20.INIT1 = 16'h5666;
    defparam add_1060_20.INJECT1_0 = "NO";
    defparam add_1060_20.INJECT1_1 = "NO";
    CCU2D add_1060_18 (.A0(d2[16]), .B0(d3[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[17]), .B1(d3[17]), .C1(GND_net), .D1(GND_net), .CIN(n10731), 
          .COUT(n10732), .S0(d3_71__N_562[16]), .S1(d3_71__N_562[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1060_18.INIT0 = 16'h5666;
    defparam add_1060_18.INIT1 = 16'h5666;
    defparam add_1060_18.INJECT1_0 = "NO";
    defparam add_1060_18.INJECT1_1 = "NO";
    CCU2D add_1060_16 (.A0(d2[14]), .B0(d3[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[15]), .B1(d3[15]), .C1(GND_net), .D1(GND_net), .CIN(n10730), 
          .COUT(n10731), .S0(d3_71__N_562[14]), .S1(d3_71__N_562[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1060_16.INIT0 = 16'h5666;
    defparam add_1060_16.INIT1 = 16'h5666;
    defparam add_1060_16.INJECT1_0 = "NO";
    defparam add_1060_16.INJECT1_1 = "NO";
    CCU2D add_1060_14 (.A0(d2[12]), .B0(d3[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[13]), .B1(d3[13]), .C1(GND_net), .D1(GND_net), .CIN(n10729), 
          .COUT(n10730), .S0(d3_71__N_562[12]), .S1(d3_71__N_562[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1060_14.INIT0 = 16'h5666;
    defparam add_1060_14.INIT1 = 16'h5666;
    defparam add_1060_14.INJECT1_0 = "NO";
    defparam add_1060_14.INJECT1_1 = "NO";
    CCU2D add_1060_12 (.A0(d2[10]), .B0(d3[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[11]), .B1(d3[11]), .C1(GND_net), .D1(GND_net), .CIN(n10728), 
          .COUT(n10729), .S0(d3_71__N_562[10]), .S1(d3_71__N_562[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1060_12.INIT0 = 16'h5666;
    defparam add_1060_12.INIT1 = 16'h5666;
    defparam add_1060_12.INJECT1_0 = "NO";
    defparam add_1060_12.INJECT1_1 = "NO";
    CCU2D add_1060_10 (.A0(d2[8]), .B0(d3[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[9]), .B1(d3[9]), .C1(GND_net), .D1(GND_net), .CIN(n10727), 
          .COUT(n10728), .S0(d3_71__N_562[8]), .S1(d3_71__N_562[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1060_10.INIT0 = 16'h5666;
    defparam add_1060_10.INIT1 = 16'h5666;
    defparam add_1060_10.INJECT1_0 = "NO";
    defparam add_1060_10.INJECT1_1 = "NO";
    CCU2D add_1060_8 (.A0(d2[6]), .B0(d3[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[7]), .B1(d3[7]), .C1(GND_net), .D1(GND_net), .CIN(n10726), 
          .COUT(n10727), .S0(d3_71__N_562[6]), .S1(d3_71__N_562[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1060_8.INIT0 = 16'h5666;
    defparam add_1060_8.INIT1 = 16'h5666;
    defparam add_1060_8.INJECT1_0 = "NO";
    defparam add_1060_8.INJECT1_1 = "NO";
    CCU2D add_1060_6 (.A0(d2[4]), .B0(d3[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[5]), .B1(d3[5]), .C1(GND_net), .D1(GND_net), .CIN(n10725), 
          .COUT(n10726), .S0(d3_71__N_562[4]), .S1(d3_71__N_562[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1060_6.INIT0 = 16'h5666;
    defparam add_1060_6.INIT1 = 16'h5666;
    defparam add_1060_6.INJECT1_0 = "NO";
    defparam add_1060_6.INJECT1_1 = "NO";
    CCU2D add_1060_4 (.A0(d2[2]), .B0(d3[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[3]), .B1(d3[3]), .C1(GND_net), .D1(GND_net), .CIN(n10724), 
          .COUT(n10725), .S0(d3_71__N_562[2]), .S1(d3_71__N_562[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1060_4.INIT0 = 16'h5666;
    defparam add_1060_4.INIT1 = 16'h5666;
    defparam add_1060_4.INJECT1_0 = "NO";
    defparam add_1060_4.INJECT1_1 = "NO";
    CCU2D add_1060_2 (.A0(d2[0]), .B0(d3[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[1]), .B1(d3[1]), .C1(GND_net), .D1(GND_net), .COUT(n10724), 
          .S1(d3_71__N_562[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1060_2.INIT0 = 16'h7000;
    defparam add_1060_2.INIT1 = 16'h5666;
    defparam add_1060_2.INJECT1_0 = "NO";
    defparam add_1060_2.INJECT1_1 = "NO";
    CCU2D add_1055_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10722), 
          .S0(n4451));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1055_cout.INIT0 = 16'h0000;
    defparam add_1055_cout.INIT1 = 16'h0000;
    defparam add_1055_cout.INJECT1_0 = "NO";
    defparam add_1055_cout.INJECT1_1 = "NO";
    CCU2D add_1055_36 (.A0(d1[34]), .B0(d2[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[35]), .B1(d2[35]), .C1(GND_net), .D1(GND_net), .CIN(n10721), 
          .COUT(n10722), .S0(d2_71__N_490[34]), .S1(d2_71__N_490[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1055_36.INIT0 = 16'h5666;
    defparam add_1055_36.INIT1 = 16'h5666;
    defparam add_1055_36.INJECT1_0 = "NO";
    defparam add_1055_36.INJECT1_1 = "NO";
    CCU2D add_1055_34 (.A0(d1[32]), .B0(d2[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[33]), .B1(d2[33]), .C1(GND_net), .D1(GND_net), .CIN(n10720), 
          .COUT(n10721), .S0(d2_71__N_490[32]), .S1(d2_71__N_490[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1055_34.INIT0 = 16'h5666;
    defparam add_1055_34.INIT1 = 16'h5666;
    defparam add_1055_34.INJECT1_0 = "NO";
    defparam add_1055_34.INJECT1_1 = "NO";
    CCU2D add_1055_32 (.A0(d1[30]), .B0(d2[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[31]), .B1(d2[31]), .C1(GND_net), .D1(GND_net), .CIN(n10719), 
          .COUT(n10720), .S0(d2_71__N_490[30]), .S1(d2_71__N_490[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1055_32.INIT0 = 16'h5666;
    defparam add_1055_32.INIT1 = 16'h5666;
    defparam add_1055_32.INJECT1_0 = "NO";
    defparam add_1055_32.INJECT1_1 = "NO";
    CCU2D add_1055_30 (.A0(d1[28]), .B0(d2[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[29]), .B1(d2[29]), .C1(GND_net), .D1(GND_net), .CIN(n10718), 
          .COUT(n10719), .S0(d2_71__N_490[28]), .S1(d2_71__N_490[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1055_30.INIT0 = 16'h5666;
    defparam add_1055_30.INIT1 = 16'h5666;
    defparam add_1055_30.INJECT1_0 = "NO";
    defparam add_1055_30.INJECT1_1 = "NO";
    CCU2D add_1055_28 (.A0(d1[26]), .B0(d2[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[27]), .B1(d2[27]), .C1(GND_net), .D1(GND_net), .CIN(n10717), 
          .COUT(n10718), .S0(d2_71__N_490[26]), .S1(d2_71__N_490[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1055_28.INIT0 = 16'h5666;
    defparam add_1055_28.INIT1 = 16'h5666;
    defparam add_1055_28.INJECT1_0 = "NO";
    defparam add_1055_28.INJECT1_1 = "NO";
    CCU2D add_1055_26 (.A0(d1[24]), .B0(d2[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[25]), .B1(d2[25]), .C1(GND_net), .D1(GND_net), .CIN(n10716), 
          .COUT(n10717), .S0(d2_71__N_490[24]), .S1(d2_71__N_490[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1055_26.INIT0 = 16'h5666;
    defparam add_1055_26.INIT1 = 16'h5666;
    defparam add_1055_26.INJECT1_0 = "NO";
    defparam add_1055_26.INJECT1_1 = "NO";
    CCU2D add_1055_24 (.A0(d1[22]), .B0(d2[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[23]), .B1(d2[23]), .C1(GND_net), .D1(GND_net), .CIN(n10715), 
          .COUT(n10716), .S0(d2_71__N_490[22]), .S1(d2_71__N_490[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1055_24.INIT0 = 16'h5666;
    defparam add_1055_24.INIT1 = 16'h5666;
    defparam add_1055_24.INJECT1_0 = "NO";
    defparam add_1055_24.INJECT1_1 = "NO";
    CCU2D add_1055_22 (.A0(d1[20]), .B0(d2[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[21]), .B1(d2[21]), .C1(GND_net), .D1(GND_net), .CIN(n10714), 
          .COUT(n10715), .S0(d2_71__N_490[20]), .S1(d2_71__N_490[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1055_22.INIT0 = 16'h5666;
    defparam add_1055_22.INIT1 = 16'h5666;
    defparam add_1055_22.INJECT1_0 = "NO";
    defparam add_1055_22.INJECT1_1 = "NO";
    CCU2D add_1055_20 (.A0(d1[18]), .B0(d2[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[19]), .B1(d2[19]), .C1(GND_net), .D1(GND_net), .CIN(n10713), 
          .COUT(n10714), .S0(d2_71__N_490[18]), .S1(d2_71__N_490[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1055_20.INIT0 = 16'h5666;
    defparam add_1055_20.INIT1 = 16'h5666;
    defparam add_1055_20.INJECT1_0 = "NO";
    defparam add_1055_20.INJECT1_1 = "NO";
    CCU2D add_1055_18 (.A0(d1[16]), .B0(d2[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[17]), .B1(d2[17]), .C1(GND_net), .D1(GND_net), .CIN(n10712), 
          .COUT(n10713), .S0(d2_71__N_490[16]), .S1(d2_71__N_490[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1055_18.INIT0 = 16'h5666;
    defparam add_1055_18.INIT1 = 16'h5666;
    defparam add_1055_18.INJECT1_0 = "NO";
    defparam add_1055_18.INJECT1_1 = "NO";
    CCU2D add_1055_16 (.A0(d1[14]), .B0(d2[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[15]), .B1(d2[15]), .C1(GND_net), .D1(GND_net), .CIN(n10711), 
          .COUT(n10712), .S0(d2_71__N_490[14]), .S1(d2_71__N_490[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1055_16.INIT0 = 16'h5666;
    defparam add_1055_16.INIT1 = 16'h5666;
    defparam add_1055_16.INJECT1_0 = "NO";
    defparam add_1055_16.INJECT1_1 = "NO";
    CCU2D add_1055_14 (.A0(d1[12]), .B0(d2[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[13]), .B1(d2[13]), .C1(GND_net), .D1(GND_net), .CIN(n10710), 
          .COUT(n10711), .S0(d2_71__N_490[12]), .S1(d2_71__N_490[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1055_14.INIT0 = 16'h5666;
    defparam add_1055_14.INIT1 = 16'h5666;
    defparam add_1055_14.INJECT1_0 = "NO";
    defparam add_1055_14.INJECT1_1 = "NO";
    CCU2D add_1055_12 (.A0(d1[10]), .B0(d2[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[11]), .B1(d2[11]), .C1(GND_net), .D1(GND_net), .CIN(n10709), 
          .COUT(n10710), .S0(d2_71__N_490[10]), .S1(d2_71__N_490[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1055_12.INIT0 = 16'h5666;
    defparam add_1055_12.INIT1 = 16'h5666;
    defparam add_1055_12.INJECT1_0 = "NO";
    defparam add_1055_12.INJECT1_1 = "NO";
    CCU2D add_1055_10 (.A0(d1[8]), .B0(d2[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[9]), .B1(d2[9]), .C1(GND_net), .D1(GND_net), .CIN(n10708), 
          .COUT(n10709), .S0(d2_71__N_490[8]), .S1(d2_71__N_490[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1055_10.INIT0 = 16'h5666;
    defparam add_1055_10.INIT1 = 16'h5666;
    defparam add_1055_10.INJECT1_0 = "NO";
    defparam add_1055_10.INJECT1_1 = "NO";
    CCU2D add_1055_8 (.A0(d1[6]), .B0(d2[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[7]), .B1(d2[7]), .C1(GND_net), .D1(GND_net), .CIN(n10707), 
          .COUT(n10708), .S0(d2_71__N_490[6]), .S1(d2_71__N_490[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1055_8.INIT0 = 16'h5666;
    defparam add_1055_8.INIT1 = 16'h5666;
    defparam add_1055_8.INJECT1_0 = "NO";
    defparam add_1055_8.INJECT1_1 = "NO";
    CCU2D add_1055_6 (.A0(d1[4]), .B0(d2[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[5]), .B1(d2[5]), .C1(GND_net), .D1(GND_net), .CIN(n10706), 
          .COUT(n10707), .S0(d2_71__N_490[4]), .S1(d2_71__N_490[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1055_6.INIT0 = 16'h5666;
    defparam add_1055_6.INIT1 = 16'h5666;
    defparam add_1055_6.INJECT1_0 = "NO";
    defparam add_1055_6.INJECT1_1 = "NO";
    CCU2D add_1055_4 (.A0(d1[2]), .B0(d2[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[3]), .B1(d2[3]), .C1(GND_net), .D1(GND_net), .CIN(n10705), 
          .COUT(n10706), .S0(d2_71__N_490[2]), .S1(d2_71__N_490[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1055_4.INIT0 = 16'h5666;
    defparam add_1055_4.INIT1 = 16'h5666;
    defparam add_1055_4.INJECT1_0 = "NO";
    defparam add_1055_4.INJECT1_1 = "NO";
    CCU2D add_1055_2 (.A0(d1[0]), .B0(d2[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[1]), .B1(d2[1]), .C1(GND_net), .D1(GND_net), .COUT(n10705), 
          .S1(d2_71__N_490[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1055_2.INIT0 = 16'h7000;
    defparam add_1055_2.INIT1 = 16'h5666;
    defparam add_1055_2.INJECT1_0 = "NO";
    defparam add_1055_2.INJECT1_1 = "NO";
    CCU2D add_1050_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10660), 
          .S0(n4299));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1050_cout.INIT0 = 16'h0000;
    defparam add_1050_cout.INIT1 = 16'h0000;
    defparam add_1050_cout.INJECT1_0 = "NO";
    defparam add_1050_cout.INJECT1_1 = "NO";
    CCU2D add_1050_36 (.A0(MixerOutSin[11]), .B0(d1[34]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[35]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10659), .COUT(n10660), .S0(d1_71__N_418[34]), 
          .S1(d1_71__N_418[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1050_36.INIT0 = 16'h5666;
    defparam add_1050_36.INIT1 = 16'h5666;
    defparam add_1050_36.INJECT1_0 = "NO";
    defparam add_1050_36.INJECT1_1 = "NO";
    CCU2D add_1050_34 (.A0(MixerOutSin[11]), .B0(d1[32]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[33]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10658), .COUT(n10659), .S0(d1_71__N_418[32]), 
          .S1(d1_71__N_418[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1050_34.INIT0 = 16'h5666;
    defparam add_1050_34.INIT1 = 16'h5666;
    defparam add_1050_34.INJECT1_0 = "NO";
    defparam add_1050_34.INJECT1_1 = "NO";
    CCU2D add_1050_32 (.A0(MixerOutSin[11]), .B0(d1[30]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10657), .COUT(n10658), .S0(d1_71__N_418[30]), 
          .S1(d1_71__N_418[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1050_32.INIT0 = 16'h5666;
    defparam add_1050_32.INIT1 = 16'h5666;
    defparam add_1050_32.INJECT1_0 = "NO";
    defparam add_1050_32.INJECT1_1 = "NO";
    CCU2D add_1050_30 (.A0(MixerOutSin[11]), .B0(d1[28]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10656), .COUT(n10657), .S0(d1_71__N_418[28]), 
          .S1(d1_71__N_418[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1050_30.INIT0 = 16'h5666;
    defparam add_1050_30.INIT1 = 16'h5666;
    defparam add_1050_30.INJECT1_0 = "NO";
    defparam add_1050_30.INJECT1_1 = "NO";
    CCU2D add_1050_28 (.A0(MixerOutSin[11]), .B0(d1[26]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10655), .COUT(n10656), .S0(d1_71__N_418[26]), 
          .S1(d1_71__N_418[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1050_28.INIT0 = 16'h5666;
    defparam add_1050_28.INIT1 = 16'h5666;
    defparam add_1050_28.INJECT1_0 = "NO";
    defparam add_1050_28.INJECT1_1 = "NO";
    CCU2D add_1050_26 (.A0(MixerOutSin[11]), .B0(d1[24]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10654), .COUT(n10655), .S0(d1_71__N_418[24]), 
          .S1(d1_71__N_418[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1050_26.INIT0 = 16'h5666;
    defparam add_1050_26.INIT1 = 16'h5666;
    defparam add_1050_26.INJECT1_0 = "NO";
    defparam add_1050_26.INJECT1_1 = "NO";
    CCU2D add_1050_24 (.A0(MixerOutSin[11]), .B0(d1[22]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10653), .COUT(n10654), .S0(d1_71__N_418[22]), 
          .S1(d1_71__N_418[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1050_24.INIT0 = 16'h5666;
    defparam add_1050_24.INIT1 = 16'h5666;
    defparam add_1050_24.INJECT1_0 = "NO";
    defparam add_1050_24.INJECT1_1 = "NO";
    CCU2D add_1050_22 (.A0(MixerOutSin[11]), .B0(d1[20]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10652), .COUT(n10653), .S0(d1_71__N_418[20]), 
          .S1(d1_71__N_418[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1050_22.INIT0 = 16'h5666;
    defparam add_1050_22.INIT1 = 16'h5666;
    defparam add_1050_22.INJECT1_0 = "NO";
    defparam add_1050_22.INJECT1_1 = "NO";
    CCU2D add_1050_20 (.A0(MixerOutSin[11]), .B0(d1[18]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10651), .COUT(n10652), .S0(d1_71__N_418[18]), 
          .S1(d1_71__N_418[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1050_20.INIT0 = 16'h5666;
    defparam add_1050_20.INIT1 = 16'h5666;
    defparam add_1050_20.INJECT1_0 = "NO";
    defparam add_1050_20.INJECT1_1 = "NO";
    CCU2D add_1050_18 (.A0(MixerOutSin[11]), .B0(d1[16]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10650), .COUT(n10651), .S0(d1_71__N_418[16]), 
          .S1(d1_71__N_418[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1050_18.INIT0 = 16'h5666;
    defparam add_1050_18.INIT1 = 16'h5666;
    defparam add_1050_18.INJECT1_0 = "NO";
    defparam add_1050_18.INJECT1_1 = "NO";
    CCU2D add_1050_16 (.A0(MixerOutSin[11]), .B0(d1[14]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10649), .COUT(n10650), .S0(d1_71__N_418[14]), 
          .S1(d1_71__N_418[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1050_16.INIT0 = 16'h5666;
    defparam add_1050_16.INIT1 = 16'h5666;
    defparam add_1050_16.INJECT1_0 = "NO";
    defparam add_1050_16.INJECT1_1 = "NO";
    CCU2D add_1050_14 (.A0(MixerOutSin[11]), .B0(d1[12]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10648), .COUT(n10649), .S0(d1_71__N_418[12]), 
          .S1(d1_71__N_418[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1050_14.INIT0 = 16'h5666;
    defparam add_1050_14.INIT1 = 16'h5666;
    defparam add_1050_14.INJECT1_0 = "NO";
    defparam add_1050_14.INJECT1_1 = "NO";
    CCU2D add_1050_12 (.A0(MixerOutSin[10]), .B0(d1[10]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10647), .COUT(n10648), .S0(d1_71__N_418[10]), 
          .S1(d1_71__N_418[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1050_12.INIT0 = 16'h5666;
    defparam add_1050_12.INIT1 = 16'h5666;
    defparam add_1050_12.INJECT1_0 = "NO";
    defparam add_1050_12.INJECT1_1 = "NO";
    CCU2D add_1050_10 (.A0(MixerOutSin[8]), .B0(d1[8]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[9]), .B1(d1[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10646), .COUT(n10647), .S0(d1_71__N_418[8]), 
          .S1(d1_71__N_418[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1050_10.INIT0 = 16'h5666;
    defparam add_1050_10.INIT1 = 16'h5666;
    defparam add_1050_10.INJECT1_0 = "NO";
    defparam add_1050_10.INJECT1_1 = "NO";
    CCU2D add_1050_8 (.A0(MixerOutSin[6]), .B0(d1[6]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutSin[7]), .B1(d1[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10645), .COUT(n10646), .S0(d1_71__N_418[6]), .S1(d1_71__N_418[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1050_8.INIT0 = 16'h5666;
    defparam add_1050_8.INIT1 = 16'h5666;
    defparam add_1050_8.INJECT1_0 = "NO";
    defparam add_1050_8.INJECT1_1 = "NO";
    CCU2D add_1050_6 (.A0(MixerOutSin[4]), .B0(d1[4]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutSin[5]), .B1(d1[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10644), .COUT(n10645), .S0(d1_71__N_418[4]), .S1(d1_71__N_418[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1050_6.INIT0 = 16'h5666;
    defparam add_1050_6.INIT1 = 16'h5666;
    defparam add_1050_6.INJECT1_0 = "NO";
    defparam add_1050_6.INJECT1_1 = "NO";
    CCU2D add_1050_4 (.A0(MixerOutSin[2]), .B0(d1[2]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutSin[3]), .B1(d1[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10643), .COUT(n10644), .S0(d1_71__N_418[2]), .S1(d1_71__N_418[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1050_4.INIT0 = 16'h5666;
    defparam add_1050_4.INIT1 = 16'h5666;
    defparam add_1050_4.INJECT1_0 = "NO";
    defparam add_1050_4.INJECT1_1 = "NO";
    CCU2D add_1050_2 (.A0(MixerOutSin[0]), .B0(d1[0]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutSin[1]), .B1(d1[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n10643), .S1(d1_71__N_418[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1050_2.INIT0 = 16'h7000;
    defparam add_1050_2.INIT1 = 16'h5666;
    defparam add_1050_2.INJECT1_0 = "NO";
    defparam add_1050_2.INJECT1_1 = "NO";
    CCU2D add_1140_37 (.A0(d6[35]), .B0(d_d6[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n12131), 
          .S0(d7_71__N_1531[35]), .S1(n7035));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1140_37.INIT0 = 16'h5999;
    defparam add_1140_37.INIT1 = 16'h0000;
    defparam add_1140_37.INJECT1_0 = "NO";
    defparam add_1140_37.INJECT1_1 = "NO";
    CCU2D add_1140_35 (.A0(d6[33]), .B0(d_d6[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[34]), .B1(d_d6[34]), .C1(GND_net), .D1(GND_net), .CIN(n12130), 
          .COUT(n12131), .S0(d7_71__N_1531[33]), .S1(d7_71__N_1531[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1140_35.INIT0 = 16'h5999;
    defparam add_1140_35.INIT1 = 16'h5999;
    defparam add_1140_35.INJECT1_0 = "NO";
    defparam add_1140_35.INJECT1_1 = "NO";
    CCU2D add_1140_33 (.A0(d6[31]), .B0(d_d6[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[32]), .B1(d_d6[32]), .C1(GND_net), .D1(GND_net), .CIN(n12129), 
          .COUT(n12130), .S0(d7_71__N_1531[31]), .S1(d7_71__N_1531[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1140_33.INIT0 = 16'h5999;
    defparam add_1140_33.INIT1 = 16'h5999;
    defparam add_1140_33.INJECT1_0 = "NO";
    defparam add_1140_33.INJECT1_1 = "NO";
    CCU2D add_1140_31 (.A0(d6[29]), .B0(d_d6[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[30]), .B1(d_d6[30]), .C1(GND_net), .D1(GND_net), .CIN(n12128), 
          .COUT(n12129), .S0(d7_71__N_1531[29]), .S1(d7_71__N_1531[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1140_31.INIT0 = 16'h5999;
    defparam add_1140_31.INIT1 = 16'h5999;
    defparam add_1140_31.INJECT1_0 = "NO";
    defparam add_1140_31.INJECT1_1 = "NO";
    CCU2D add_1140_29 (.A0(d6[27]), .B0(d_d6[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[28]), .B1(d_d6[28]), .C1(GND_net), .D1(GND_net), .CIN(n12127), 
          .COUT(n12128), .S0(d7_71__N_1531[27]), .S1(d7_71__N_1531[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1140_29.INIT0 = 16'h5999;
    defparam add_1140_29.INIT1 = 16'h5999;
    defparam add_1140_29.INJECT1_0 = "NO";
    defparam add_1140_29.INJECT1_1 = "NO";
    CCU2D add_1140_27 (.A0(d6[25]), .B0(d_d6[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[26]), .B1(d_d6[26]), .C1(GND_net), .D1(GND_net), .CIN(n12126), 
          .COUT(n12127), .S0(d7_71__N_1531[25]), .S1(d7_71__N_1531[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1140_27.INIT0 = 16'h5999;
    defparam add_1140_27.INIT1 = 16'h5999;
    defparam add_1140_27.INJECT1_0 = "NO";
    defparam add_1140_27.INJECT1_1 = "NO";
    CCU2D add_1140_25 (.A0(d6[23]), .B0(d_d6[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[24]), .B1(d_d6[24]), .C1(GND_net), .D1(GND_net), .CIN(n12125), 
          .COUT(n12126), .S0(d7_71__N_1531[23]), .S1(d7_71__N_1531[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1140_25.INIT0 = 16'h5999;
    defparam add_1140_25.INIT1 = 16'h5999;
    defparam add_1140_25.INJECT1_0 = "NO";
    defparam add_1140_25.INJECT1_1 = "NO";
    CCU2D add_1140_23 (.A0(d6[21]), .B0(d_d6[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[22]), .B1(d_d6[22]), .C1(GND_net), .D1(GND_net), .CIN(n12124), 
          .COUT(n12125), .S0(d7_71__N_1531[21]), .S1(d7_71__N_1531[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1140_23.INIT0 = 16'h5999;
    defparam add_1140_23.INIT1 = 16'h5999;
    defparam add_1140_23.INJECT1_0 = "NO";
    defparam add_1140_23.INJECT1_1 = "NO";
    CCU2D add_1135_37 (.A0(d7[35]), .B0(d_d7[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11484), 
          .S0(d8_71__N_1603[35]), .S1(n6883));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1135_37.INIT0 = 16'h5999;
    defparam add_1135_37.INIT1 = 16'h0000;
    defparam add_1135_37.INJECT1_0 = "NO";
    defparam add_1135_37.INJECT1_1 = "NO";
    CCU2D add_1135_35 (.A0(d7[33]), .B0(d_d7[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[34]), .B1(d_d7[34]), .C1(GND_net), .D1(GND_net), .CIN(n11483), 
          .COUT(n11484), .S0(d8_71__N_1603[33]), .S1(d8_71__N_1603[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1135_35.INIT0 = 16'h5999;
    defparam add_1135_35.INIT1 = 16'h5999;
    defparam add_1135_35.INJECT1_0 = "NO";
    defparam add_1135_35.INJECT1_1 = "NO";
    CCU2D add_1135_33 (.A0(d7[31]), .B0(d_d7[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[32]), .B1(d_d7[32]), .C1(GND_net), .D1(GND_net), .CIN(n11482), 
          .COUT(n11483), .S0(d8_71__N_1603[31]), .S1(d8_71__N_1603[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1135_33.INIT0 = 16'h5999;
    defparam add_1135_33.INIT1 = 16'h5999;
    defparam add_1135_33.INJECT1_0 = "NO";
    defparam add_1135_33.INJECT1_1 = "NO";
    CCU2D add_1135_31 (.A0(d7[29]), .B0(d_d7[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[30]), .B1(d_d7[30]), .C1(GND_net), .D1(GND_net), .CIN(n11481), 
          .COUT(n11482), .S0(d8_71__N_1603[29]), .S1(d8_71__N_1603[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1135_31.INIT0 = 16'h5999;
    defparam add_1135_31.INIT1 = 16'h5999;
    defparam add_1135_31.INJECT1_0 = "NO";
    defparam add_1135_31.INJECT1_1 = "NO";
    CCU2D add_1135_29 (.A0(d7[27]), .B0(d_d7[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[28]), .B1(d_d7[28]), .C1(GND_net), .D1(GND_net), .CIN(n11480), 
          .COUT(n11481), .S0(d8_71__N_1603[27]), .S1(d8_71__N_1603[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1135_29.INIT0 = 16'h5999;
    defparam add_1135_29.INIT1 = 16'h5999;
    defparam add_1135_29.INJECT1_0 = "NO";
    defparam add_1135_29.INJECT1_1 = "NO";
    CCU2D add_1135_27 (.A0(d7[25]), .B0(d_d7[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[26]), .B1(d_d7[26]), .C1(GND_net), .D1(GND_net), .CIN(n11479), 
          .COUT(n11480), .S0(d8_71__N_1603[25]), .S1(d8_71__N_1603[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1135_27.INIT0 = 16'h5999;
    defparam add_1135_27.INIT1 = 16'h5999;
    defparam add_1135_27.INJECT1_0 = "NO";
    defparam add_1135_27.INJECT1_1 = "NO";
    CCU2D add_1135_25 (.A0(d7[23]), .B0(d_d7[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[24]), .B1(d_d7[24]), .C1(GND_net), .D1(GND_net), .CIN(n11478), 
          .COUT(n11479), .S0(d8_71__N_1603[23]), .S1(d8_71__N_1603[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1135_25.INIT0 = 16'h5999;
    defparam add_1135_25.INIT1 = 16'h5999;
    defparam add_1135_25.INJECT1_0 = "NO";
    defparam add_1135_25.INJECT1_1 = "NO";
    CCU2D add_1135_23 (.A0(d7[21]), .B0(d_d7[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[22]), .B1(d_d7[22]), .C1(GND_net), .D1(GND_net), .CIN(n11477), 
          .COUT(n11478), .S0(d8_71__N_1603[21]), .S1(d8_71__N_1603[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1135_23.INIT0 = 16'h5999;
    defparam add_1135_23.INIT1 = 16'h5999;
    defparam add_1135_23.INJECT1_0 = "NO";
    defparam add_1135_23.INJECT1_1 = "NO";
    CCU2D add_1135_21 (.A0(d7[19]), .B0(d_d7[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[20]), .B1(d_d7[20]), .C1(GND_net), .D1(GND_net), .CIN(n11476), 
          .COUT(n11477), .S0(d8_71__N_1603[19]), .S1(d8_71__N_1603[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1135_21.INIT0 = 16'h5999;
    defparam add_1135_21.INIT1 = 16'h5999;
    defparam add_1135_21.INJECT1_0 = "NO";
    defparam add_1135_21.INJECT1_1 = "NO";
    CCU2D add_1135_19 (.A0(d7[17]), .B0(d_d7[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[18]), .B1(d_d7[18]), .C1(GND_net), .D1(GND_net), .CIN(n11475), 
          .COUT(n11476), .S0(d8_71__N_1603[17]), .S1(d8_71__N_1603[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1135_19.INIT0 = 16'h5999;
    defparam add_1135_19.INIT1 = 16'h5999;
    defparam add_1135_19.INJECT1_0 = "NO";
    defparam add_1135_19.INJECT1_1 = "NO";
    CCU2D add_1135_17 (.A0(d7[15]), .B0(d_d7[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[16]), .B1(d_d7[16]), .C1(GND_net), .D1(GND_net), .CIN(n11474), 
          .COUT(n11475), .S0(d8_71__N_1603[15]), .S1(d8_71__N_1603[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1135_17.INIT0 = 16'h5999;
    defparam add_1135_17.INIT1 = 16'h5999;
    defparam add_1135_17.INJECT1_0 = "NO";
    defparam add_1135_17.INJECT1_1 = "NO";
    CCU2D add_1135_15 (.A0(d7[13]), .B0(d_d7[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[14]), .B1(d_d7[14]), .C1(GND_net), .D1(GND_net), .CIN(n11473), 
          .COUT(n11474), .S0(d8_71__N_1603[13]), .S1(d8_71__N_1603[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1135_15.INIT0 = 16'h5999;
    defparam add_1135_15.INIT1 = 16'h5999;
    defparam add_1135_15.INJECT1_0 = "NO";
    defparam add_1135_15.INJECT1_1 = "NO";
    CCU2D add_1135_13 (.A0(d7[11]), .B0(d_d7[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[12]), .B1(d_d7[12]), .C1(GND_net), .D1(GND_net), .CIN(n11472), 
          .COUT(n11473), .S0(d8_71__N_1603[11]), .S1(d8_71__N_1603[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1135_13.INIT0 = 16'h5999;
    defparam add_1135_13.INIT1 = 16'h5999;
    defparam add_1135_13.INJECT1_0 = "NO";
    defparam add_1135_13.INJECT1_1 = "NO";
    CCU2D add_1135_11 (.A0(d7[9]), .B0(d_d7[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[10]), .B1(d_d7[10]), .C1(GND_net), .D1(GND_net), .CIN(n11471), 
          .COUT(n11472), .S0(d8_71__N_1603[9]), .S1(d8_71__N_1603[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1135_11.INIT0 = 16'h5999;
    defparam add_1135_11.INIT1 = 16'h5999;
    defparam add_1135_11.INJECT1_0 = "NO";
    defparam add_1135_11.INJECT1_1 = "NO";
    CCU2D add_1135_9 (.A0(d7[7]), .B0(d_d7[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[8]), .B1(d_d7[8]), .C1(GND_net), .D1(GND_net), .CIN(n11470), 
          .COUT(n11471), .S0(d8_71__N_1603[7]), .S1(d8_71__N_1603[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1135_9.INIT0 = 16'h5999;
    defparam add_1135_9.INIT1 = 16'h5999;
    defparam add_1135_9.INJECT1_0 = "NO";
    defparam add_1135_9.INJECT1_1 = "NO";
    CCU2D add_1135_7 (.A0(d7[5]), .B0(d_d7[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[6]), .B1(d_d7[6]), .C1(GND_net), .D1(GND_net), .CIN(n11469), 
          .COUT(n11470), .S0(d8_71__N_1603[5]), .S1(d8_71__N_1603[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1135_7.INIT0 = 16'h5999;
    defparam add_1135_7.INIT1 = 16'h5999;
    defparam add_1135_7.INJECT1_0 = "NO";
    defparam add_1135_7.INJECT1_1 = "NO";
    CCU2D add_1135_5 (.A0(d7[3]), .B0(d_d7[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[4]), .B1(d_d7[4]), .C1(GND_net), .D1(GND_net), .CIN(n11468), 
          .COUT(n11469), .S0(d8_71__N_1603[3]), .S1(d8_71__N_1603[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1135_5.INIT0 = 16'h5999;
    defparam add_1135_5.INIT1 = 16'h5999;
    defparam add_1135_5.INJECT1_0 = "NO";
    defparam add_1135_5.INJECT1_1 = "NO";
    CCU2D add_1135_3 (.A0(d7[1]), .B0(d_d7[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[2]), .B1(d_d7[2]), .C1(GND_net), .D1(GND_net), .CIN(n11467), 
          .COUT(n11468), .S0(d8_71__N_1603[1]), .S1(d8_71__N_1603[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1135_3.INIT0 = 16'h5999;
    defparam add_1135_3.INIT1 = 16'h5999;
    defparam add_1135_3.INJECT1_0 = "NO";
    defparam add_1135_3.INJECT1_1 = "NO";
    CCU2D add_1135_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d7[0]), .B1(d_d7[0]), .C1(GND_net), .D1(GND_net), .COUT(n11467), 
          .S1(d8_71__N_1603[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1135_1.INIT0 = 16'h0000;
    defparam add_1135_1.INIT1 = 16'h5999;
    defparam add_1135_1.INJECT1_0 = "NO";
    defparam add_1135_1.INJECT1_1 = "NO";
    CCU2D add_1105_37 (.A0(d9[35]), .B0(d_d9[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11348), 
          .S1(n5971));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1105_37.INIT0 = 16'h5999;
    defparam add_1105_37.INIT1 = 16'h0000;
    defparam add_1105_37.INJECT1_0 = "NO";
    defparam add_1105_37.INJECT1_1 = "NO";
    CCU2D add_1105_35 (.A0(d9[33]), .B0(d_d9[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[34]), .B1(d_d9[34]), .C1(GND_net), .D1(GND_net), .CIN(n11347), 
          .COUT(n11348));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1105_35.INIT0 = 16'h5999;
    defparam add_1105_35.INIT1 = 16'h5999;
    defparam add_1105_35.INJECT1_0 = "NO";
    defparam add_1105_35.INJECT1_1 = "NO";
    CCU2D add_1105_33 (.A0(d9[31]), .B0(d_d9[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[32]), .B1(d_d9[32]), .C1(GND_net), .D1(GND_net), .CIN(n11346), 
          .COUT(n11347));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1105_33.INIT0 = 16'h5999;
    defparam add_1105_33.INIT1 = 16'h5999;
    defparam add_1105_33.INJECT1_0 = "NO";
    defparam add_1105_33.INJECT1_1 = "NO";
    CCU2D add_1105_31 (.A0(d9[29]), .B0(d_d9[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[30]), .B1(d_d9[30]), .C1(GND_net), .D1(GND_net), .CIN(n11345), 
          .COUT(n11346));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1105_31.INIT0 = 16'h5999;
    defparam add_1105_31.INIT1 = 16'h5999;
    defparam add_1105_31.INJECT1_0 = "NO";
    defparam add_1105_31.INJECT1_1 = "NO";
    CCU2D add_1105_29 (.A0(d9[27]), .B0(d_d9[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[28]), .B1(d_d9[28]), .C1(GND_net), .D1(GND_net), .CIN(n11344), 
          .COUT(n11345));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1105_29.INIT0 = 16'h5999;
    defparam add_1105_29.INIT1 = 16'h5999;
    defparam add_1105_29.INJECT1_0 = "NO";
    defparam add_1105_29.INJECT1_1 = "NO";
    CCU2D add_1105_27 (.A0(d9[25]), .B0(d_d9[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[26]), .B1(d_d9[26]), .C1(GND_net), .D1(GND_net), .CIN(n11343), 
          .COUT(n11344));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1105_27.INIT0 = 16'h5999;
    defparam add_1105_27.INIT1 = 16'h5999;
    defparam add_1105_27.INJECT1_0 = "NO";
    defparam add_1105_27.INJECT1_1 = "NO";
    CCU2D add_1105_25 (.A0(d9[23]), .B0(d_d9[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[24]), .B1(d_d9[24]), .C1(GND_net), .D1(GND_net), .CIN(n11342), 
          .COUT(n11343));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1105_25.INIT0 = 16'h5999;
    defparam add_1105_25.INIT1 = 16'h5999;
    defparam add_1105_25.INJECT1_0 = "NO";
    defparam add_1105_25.INJECT1_1 = "NO";
    CCU2D add_1105_23 (.A0(d9[21]), .B0(d_d9[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[22]), .B1(d_d9[22]), .C1(GND_net), .D1(GND_net), .CIN(n11341), 
          .COUT(n11342));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1105_23.INIT0 = 16'h5999;
    defparam add_1105_23.INIT1 = 16'h5999;
    defparam add_1105_23.INJECT1_0 = "NO";
    defparam add_1105_23.INJECT1_1 = "NO";
    CCU2D add_1105_21 (.A0(d9[19]), .B0(d_d9[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[20]), .B1(d_d9[20]), .C1(GND_net), .D1(GND_net), .CIN(n11340), 
          .COUT(n11341));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1105_21.INIT0 = 16'h5999;
    defparam add_1105_21.INIT1 = 16'h5999;
    defparam add_1105_21.INJECT1_0 = "NO";
    defparam add_1105_21.INJECT1_1 = "NO";
    CCU2D add_1105_19 (.A0(d9[17]), .B0(d_d9[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[18]), .B1(d_d9[18]), .C1(GND_net), .D1(GND_net), .CIN(n11339), 
          .COUT(n11340));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1105_19.INIT0 = 16'h5999;
    defparam add_1105_19.INIT1 = 16'h5999;
    defparam add_1105_19.INJECT1_0 = "NO";
    defparam add_1105_19.INJECT1_1 = "NO";
    CCU2D add_1105_17 (.A0(d9[15]), .B0(d_d9[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[16]), .B1(d_d9[16]), .C1(GND_net), .D1(GND_net), .CIN(n11338), 
          .COUT(n11339));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1105_17.INIT0 = 16'h5999;
    defparam add_1105_17.INIT1 = 16'h5999;
    defparam add_1105_17.INJECT1_0 = "NO";
    defparam add_1105_17.INJECT1_1 = "NO";
    CCU2D add_1105_15 (.A0(d9[13]), .B0(d_d9[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[14]), .B1(d_d9[14]), .C1(GND_net), .D1(GND_net), .CIN(n11337), 
          .COUT(n11338));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1105_15.INIT0 = 16'h5999;
    defparam add_1105_15.INIT1 = 16'h5999;
    defparam add_1105_15.INJECT1_0 = "NO";
    defparam add_1105_15.INJECT1_1 = "NO";
    CCU2D add_1105_13 (.A0(d9[11]), .B0(d_d9[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[12]), .B1(d_d9[12]), .C1(GND_net), .D1(GND_net), .CIN(n11336), 
          .COUT(n11337));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1105_13.INIT0 = 16'h5999;
    defparam add_1105_13.INIT1 = 16'h5999;
    defparam add_1105_13.INJECT1_0 = "NO";
    defparam add_1105_13.INJECT1_1 = "NO";
    LUT4 i1_2_lut (.A(n375[11]), .B(n54), .Z(count_15__N_1442[11])) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 i4593_2_lut (.A(MixerOutSin[0]), .B(d1[0]), .Z(d1_71__N_418[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4593_2_lut.init = 16'h6666;
    CCU2D add_1140_21 (.A0(d6[19]), .B0(d_d6[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[20]), .B1(d_d6[20]), .C1(GND_net), .D1(GND_net), .CIN(n12123), 
          .COUT(n12124), .S0(d7_71__N_1531[19]), .S1(d7_71__N_1531[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1140_21.INIT0 = 16'h5999;
    defparam add_1140_21.INIT1 = 16'h5999;
    defparam add_1140_21.INJECT1_0 = "NO";
    defparam add_1140_21.INJECT1_1 = "NO";
    LUT4 shift_right_31_i61_3_lut (.A(d10[60]), .B(d10[61]), .C(\CICGain[0] ), 
         .Z(n61_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i61_3_lut.init = 16'hcaca;
    CCU2D add_1140_19 (.A0(d6[17]), .B0(d_d6[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[18]), .B1(d_d6[18]), .C1(GND_net), .D1(GND_net), .CIN(n12122), 
          .COUT(n12123), .S0(d7_71__N_1531[17]), .S1(d7_71__N_1531[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1140_19.INIT0 = 16'h5999;
    defparam add_1140_19.INIT1 = 16'h5999;
    defparam add_1140_19.INJECT1_0 = "NO";
    defparam add_1140_19.INJECT1_1 = "NO";
    CCU2D add_1140_17 (.A0(d6[15]), .B0(d_d6[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[16]), .B1(d_d6[16]), .C1(GND_net), .D1(GND_net), .CIN(n12121), 
          .COUT(n12122), .S0(d7_71__N_1531[15]), .S1(d7_71__N_1531[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1140_17.INIT0 = 16'h5999;
    defparam add_1140_17.INIT1 = 16'h5999;
    defparam add_1140_17.INJECT1_0 = "NO";
    defparam add_1140_17.INJECT1_1 = "NO";
    CCU2D add_1140_15 (.A0(d6[13]), .B0(d_d6[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[14]), .B1(d_d6[14]), .C1(GND_net), .D1(GND_net), .CIN(n12120), 
          .COUT(n12121), .S0(d7_71__N_1531[13]), .S1(d7_71__N_1531[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1140_15.INIT0 = 16'h5999;
    defparam add_1140_15.INIT1 = 16'h5999;
    defparam add_1140_15.INJECT1_0 = "NO";
    defparam add_1140_15.INJECT1_1 = "NO";
    CCU2D add_1140_13 (.A0(d6[11]), .B0(d_d6[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[12]), .B1(d_d6[12]), .C1(GND_net), .D1(GND_net), .CIN(n12119), 
          .COUT(n12120), .S0(d7_71__N_1531[11]), .S1(d7_71__N_1531[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1140_13.INIT0 = 16'h5999;
    defparam add_1140_13.INIT1 = 16'h5999;
    defparam add_1140_13.INJECT1_0 = "NO";
    defparam add_1140_13.INJECT1_1 = "NO";
    CCU2D add_1140_11 (.A0(d6[9]), .B0(d_d6[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[10]), .B1(d_d6[10]), .C1(GND_net), .D1(GND_net), .CIN(n12118), 
          .COUT(n12119), .S0(d7_71__N_1531[9]), .S1(d7_71__N_1531[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1140_11.INIT0 = 16'h5999;
    defparam add_1140_11.INIT1 = 16'h5999;
    defparam add_1140_11.INJECT1_0 = "NO";
    defparam add_1140_11.INJECT1_1 = "NO";
    CCU2D add_1140_9 (.A0(d6[7]), .B0(d_d6[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[8]), .B1(d_d6[8]), .C1(GND_net), .D1(GND_net), .CIN(n12117), 
          .COUT(n12118), .S0(d7_71__N_1531[7]), .S1(d7_71__N_1531[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1140_9.INIT0 = 16'h5999;
    defparam add_1140_9.INIT1 = 16'h5999;
    defparam add_1140_9.INJECT1_0 = "NO";
    defparam add_1140_9.INJECT1_1 = "NO";
    CCU2D add_1140_7 (.A0(d6[5]), .B0(d_d6[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[6]), .B1(d_d6[6]), .C1(GND_net), .D1(GND_net), .CIN(n12116), 
          .COUT(n12117), .S0(d7_71__N_1531[5]), .S1(d7_71__N_1531[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1140_7.INIT0 = 16'h5999;
    defparam add_1140_7.INIT1 = 16'h5999;
    defparam add_1140_7.INJECT1_0 = "NO";
    defparam add_1140_7.INJECT1_1 = "NO";
    CCU2D add_1140_5 (.A0(d6[3]), .B0(d_d6[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[4]), .B1(d_d6[4]), .C1(GND_net), .D1(GND_net), .CIN(n12115), 
          .COUT(n12116), .S0(d7_71__N_1531[3]), .S1(d7_71__N_1531[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1140_5.INIT0 = 16'h5999;
    defparam add_1140_5.INIT1 = 16'h5999;
    defparam add_1140_5.INJECT1_0 = "NO";
    defparam add_1140_5.INJECT1_1 = "NO";
    CCU2D add_1140_3 (.A0(d6[1]), .B0(d_d6[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[2]), .B1(d_d6[2]), .C1(GND_net), .D1(GND_net), .CIN(n12114), 
          .COUT(n12115), .S0(d7_71__N_1531[1]), .S1(d7_71__N_1531[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1140_3.INIT0 = 16'h5999;
    defparam add_1140_3.INIT1 = 16'h5999;
    defparam add_1140_3.INJECT1_0 = "NO";
    defparam add_1140_3.INJECT1_1 = "NO";
    CCU2D add_1140_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d6[0]), .B1(d_d6[0]), .C1(GND_net), .D1(GND_net), .COUT(n12114), 
          .S1(d7_71__N_1531[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1140_1.INIT0 = 16'h0000;
    defparam add_1140_1.INIT1 = 16'h5999;
    defparam add_1140_1.INJECT1_0 = "NO";
    defparam add_1140_1.INJECT1_1 = "NO";
    CCU2D add_1061_22 (.A0(d2[56]), .B0(d3[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[57]), .B1(d3[57]), .C1(GND_net), .D1(GND_net), .CIN(n11907), 
          .COUT(n11908), .S0(n4604[20]), .S1(n4604[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1061_22.INIT0 = 16'h5666;
    defparam add_1061_22.INIT1 = 16'h5666;
    defparam add_1061_22.INJECT1_0 = "NO";
    defparam add_1061_22.INJECT1_1 = "NO";
    CCU2D add_1061_20 (.A0(d2[54]), .B0(d3[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[55]), .B1(d3[55]), .C1(GND_net), .D1(GND_net), .CIN(n11906), 
          .COUT(n11907), .S0(n4604[18]), .S1(n4604[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1061_20.INIT0 = 16'h5666;
    defparam add_1061_20.INIT1 = 16'h5666;
    defparam add_1061_20.INJECT1_0 = "NO";
    defparam add_1061_20.INJECT1_1 = "NO";
    CCU2D add_1061_18 (.A0(d2[52]), .B0(d3[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[53]), .B1(d3[53]), .C1(GND_net), .D1(GND_net), .CIN(n11905), 
          .COUT(n11906), .S0(n4604[16]), .S1(n4604[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1061_18.INIT0 = 16'h5666;
    defparam add_1061_18.INIT1 = 16'h5666;
    defparam add_1061_18.INJECT1_0 = "NO";
    defparam add_1061_18.INJECT1_1 = "NO";
    CCU2D add_1061_16 (.A0(d2[50]), .B0(d3[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[51]), .B1(d3[51]), .C1(GND_net), .D1(GND_net), .CIN(n11904), 
          .COUT(n11905), .S0(n4604[14]), .S1(n4604[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1061_16.INIT0 = 16'h5666;
    defparam add_1061_16.INIT1 = 16'h5666;
    defparam add_1061_16.INJECT1_0 = "NO";
    defparam add_1061_16.INJECT1_1 = "NO";
    CCU2D add_1061_14 (.A0(d2[48]), .B0(d3[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[49]), .B1(d3[49]), .C1(GND_net), .D1(GND_net), .CIN(n11903), 
          .COUT(n11904), .S0(n4604[12]), .S1(n4604[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1061_14.INIT0 = 16'h5666;
    defparam add_1061_14.INIT1 = 16'h5666;
    defparam add_1061_14.INJECT1_0 = "NO";
    defparam add_1061_14.INJECT1_1 = "NO";
    CCU2D add_1061_12 (.A0(d2[46]), .B0(d3[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[47]), .B1(d3[47]), .C1(GND_net), .D1(GND_net), .CIN(n11902), 
          .COUT(n11903), .S0(n4604[10]), .S1(n4604[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1061_12.INIT0 = 16'h5666;
    defparam add_1061_12.INIT1 = 16'h5666;
    defparam add_1061_12.INJECT1_0 = "NO";
    defparam add_1061_12.INJECT1_1 = "NO";
    CCU2D add_1061_10 (.A0(d2[44]), .B0(d3[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[45]), .B1(d3[45]), .C1(GND_net), .D1(GND_net), .CIN(n11901), 
          .COUT(n11902), .S0(n4604[8]), .S1(n4604[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1061_10.INIT0 = 16'h5666;
    defparam add_1061_10.INIT1 = 16'h5666;
    defparam add_1061_10.INJECT1_0 = "NO";
    defparam add_1061_10.INJECT1_1 = "NO";
    CCU2D add_1061_8 (.A0(d2[42]), .B0(d3[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[43]), .B1(d3[43]), .C1(GND_net), .D1(GND_net), .CIN(n11900), 
          .COUT(n11901), .S0(n4604[6]), .S1(n4604[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1061_8.INIT0 = 16'h5666;
    defparam add_1061_8.INIT1 = 16'h5666;
    defparam add_1061_8.INJECT1_0 = "NO";
    defparam add_1061_8.INJECT1_1 = "NO";
    CCU2D add_1061_6 (.A0(d2[40]), .B0(d3[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[41]), .B1(d3[41]), .C1(GND_net), .D1(GND_net), .CIN(n11899), 
          .COUT(n11900), .S0(n4604[4]), .S1(n4604[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1061_6.INIT0 = 16'h5666;
    defparam add_1061_6.INIT1 = 16'h5666;
    defparam add_1061_6.INJECT1_0 = "NO";
    defparam add_1061_6.INJECT1_1 = "NO";
    CCU2D add_1061_4 (.A0(d2[38]), .B0(d3[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[39]), .B1(d3[39]), .C1(GND_net), .D1(GND_net), .CIN(n11898), 
          .COUT(n11899), .S0(n4604[2]), .S1(n4604[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1061_4.INIT0 = 16'h5666;
    defparam add_1061_4.INIT1 = 16'h5666;
    defparam add_1061_4.INJECT1_0 = "NO";
    defparam add_1061_4.INJECT1_1 = "NO";
    CCU2D add_1061_2 (.A0(d2[36]), .B0(d3[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[37]), .B1(d3[37]), .C1(GND_net), .D1(GND_net), .COUT(n11898), 
          .S1(n4604[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1061_2.INIT0 = 16'h7000;
    defparam add_1061_2.INIT1 = 16'h5666;
    defparam add_1061_2.INJECT1_0 = "NO";
    defparam add_1061_2.INJECT1_1 = "NO";
    CCU2D add_1062_37 (.A0(d3[70]), .B0(n4603), .C0(n4604[34]), .D0(d2[70]), 
          .A1(d3[71]), .B1(n4603), .C1(n4604[35]), .D1(d2[71]), .CIN(n11895), 
          .S0(d3_71__N_562[70]), .S1(d3_71__N_562[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1062_37.INIT0 = 16'h74b8;
    defparam add_1062_37.INIT1 = 16'h74b8;
    defparam add_1062_37.INJECT1_0 = "NO";
    defparam add_1062_37.INJECT1_1 = "NO";
    CCU2D add_1062_35 (.A0(d3[68]), .B0(n4603), .C0(n4604[32]), .D0(d2[68]), 
          .A1(d3[69]), .B1(n4603), .C1(n4604[33]), .D1(d2[69]), .CIN(n11894), 
          .COUT(n11895), .S0(d3_71__N_562[68]), .S1(d3_71__N_562[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1062_35.INIT0 = 16'h74b8;
    defparam add_1062_35.INIT1 = 16'h74b8;
    defparam add_1062_35.INJECT1_0 = "NO";
    defparam add_1062_35.INJECT1_1 = "NO";
    CCU2D add_1062_33 (.A0(d3[66]), .B0(n4603), .C0(n4604[30]), .D0(d2[66]), 
          .A1(d3[67]), .B1(n4603), .C1(n4604[31]), .D1(d2[67]), .CIN(n11893), 
          .COUT(n11894), .S0(d3_71__N_562[66]), .S1(d3_71__N_562[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1062_33.INIT0 = 16'h74b8;
    defparam add_1062_33.INIT1 = 16'h74b8;
    defparam add_1062_33.INJECT1_0 = "NO";
    defparam add_1062_33.INJECT1_1 = "NO";
    CCU2D add_1062_31 (.A0(d3[64]), .B0(n4603), .C0(n4604[28]), .D0(d2[64]), 
          .A1(d3[65]), .B1(n4603), .C1(n4604[29]), .D1(d2[65]), .CIN(n11892), 
          .COUT(n11893), .S0(d3_71__N_562[64]), .S1(d3_71__N_562[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1062_31.INIT0 = 16'h74b8;
    defparam add_1062_31.INIT1 = 16'h74b8;
    defparam add_1062_31.INJECT1_0 = "NO";
    defparam add_1062_31.INJECT1_1 = "NO";
    CCU2D add_1062_29 (.A0(d3[62]), .B0(n4603), .C0(n4604[26]), .D0(d2[62]), 
          .A1(d3[63]), .B1(n4603), .C1(n4604[27]), .D1(d2[63]), .CIN(n11891), 
          .COUT(n11892), .S0(d3_71__N_562[62]), .S1(d3_71__N_562[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1062_29.INIT0 = 16'h74b8;
    defparam add_1062_29.INIT1 = 16'h74b8;
    defparam add_1062_29.INJECT1_0 = "NO";
    defparam add_1062_29.INJECT1_1 = "NO";
    CCU2D add_1062_27 (.A0(d3[60]), .B0(n4603), .C0(n4604[24]), .D0(d2[60]), 
          .A1(d3[61]), .B1(n4603), .C1(n4604[25]), .D1(d2[61]), .CIN(n11890), 
          .COUT(n11891), .S0(d3_71__N_562[60]), .S1(d3_71__N_562[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1062_27.INIT0 = 16'h74b8;
    defparam add_1062_27.INIT1 = 16'h74b8;
    defparam add_1062_27.INJECT1_0 = "NO";
    defparam add_1062_27.INJECT1_1 = "NO";
    CCU2D add_1062_25 (.A0(d3[58]), .B0(n4603), .C0(n4604[22]), .D0(d2[58]), 
          .A1(d3[59]), .B1(n4603), .C1(n4604[23]), .D1(d2[59]), .CIN(n11889), 
          .COUT(n11890), .S0(d3_71__N_562[58]), .S1(d3_71__N_562[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1062_25.INIT0 = 16'h74b8;
    defparam add_1062_25.INIT1 = 16'h74b8;
    defparam add_1062_25.INJECT1_0 = "NO";
    defparam add_1062_25.INJECT1_1 = "NO";
    CCU2D add_1062_23 (.A0(d3[56]), .B0(n4603), .C0(n4604[20]), .D0(d2[56]), 
          .A1(d3[57]), .B1(n4603), .C1(n4604[21]), .D1(d2[57]), .CIN(n11888), 
          .COUT(n11889), .S0(d3_71__N_562[56]), .S1(d3_71__N_562[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1062_23.INIT0 = 16'h74b8;
    defparam add_1062_23.INIT1 = 16'h74b8;
    defparam add_1062_23.INJECT1_0 = "NO";
    defparam add_1062_23.INJECT1_1 = "NO";
    CCU2D add_1062_21 (.A0(d3[54]), .B0(n4603), .C0(n4604[18]), .D0(d2[54]), 
          .A1(d3[55]), .B1(n4603), .C1(n4604[19]), .D1(d2[55]), .CIN(n11887), 
          .COUT(n11888), .S0(d3_71__N_562[54]), .S1(d3_71__N_562[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1062_21.INIT0 = 16'h74b8;
    defparam add_1062_21.INIT1 = 16'h74b8;
    defparam add_1062_21.INJECT1_0 = "NO";
    defparam add_1062_21.INJECT1_1 = "NO";
    CCU2D add_1062_19 (.A0(d3[52]), .B0(n4603), .C0(n4604[16]), .D0(d2[52]), 
          .A1(d3[53]), .B1(n4603), .C1(n4604[17]), .D1(d2[53]), .CIN(n11886), 
          .COUT(n11887), .S0(d3_71__N_562[52]), .S1(d3_71__N_562[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1062_19.INIT0 = 16'h74b8;
    defparam add_1062_19.INIT1 = 16'h74b8;
    defparam add_1062_19.INJECT1_0 = "NO";
    defparam add_1062_19.INJECT1_1 = "NO";
    CCU2D add_1062_17 (.A0(d3[50]), .B0(n4603), .C0(n4604[14]), .D0(d2[50]), 
          .A1(d3[51]), .B1(n4603), .C1(n4604[15]), .D1(d2[51]), .CIN(n11885), 
          .COUT(n11886), .S0(d3_71__N_562[50]), .S1(d3_71__N_562[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1062_17.INIT0 = 16'h74b8;
    defparam add_1062_17.INIT1 = 16'h74b8;
    defparam add_1062_17.INJECT1_0 = "NO";
    defparam add_1062_17.INJECT1_1 = "NO";
    CCU2D add_1062_15 (.A0(d3[48]), .B0(n4603), .C0(n4604[12]), .D0(d2[48]), 
          .A1(d3[49]), .B1(n4603), .C1(n4604[13]), .D1(d2[49]), .CIN(n11884), 
          .COUT(n11885), .S0(d3_71__N_562[48]), .S1(d3_71__N_562[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1062_15.INIT0 = 16'h74b8;
    defparam add_1062_15.INIT1 = 16'h74b8;
    defparam add_1062_15.INJECT1_0 = "NO";
    defparam add_1062_15.INJECT1_1 = "NO";
    CCU2D add_1062_13 (.A0(d3[46]), .B0(n4603), .C0(n4604[10]), .D0(d2[46]), 
          .A1(d3[47]), .B1(n4603), .C1(n4604[11]), .D1(d2[47]), .CIN(n11883), 
          .COUT(n11884), .S0(d3_71__N_562[46]), .S1(d3_71__N_562[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1062_13.INIT0 = 16'h74b8;
    defparam add_1062_13.INIT1 = 16'h74b8;
    defparam add_1062_13.INJECT1_0 = "NO";
    defparam add_1062_13.INJECT1_1 = "NO";
    CCU2D add_1062_11 (.A0(d3[44]), .B0(n4603), .C0(n4604[8]), .D0(d2[44]), 
          .A1(d3[45]), .B1(n4603), .C1(n4604[9]), .D1(d2[45]), .CIN(n11882), 
          .COUT(n11883), .S0(d3_71__N_562[44]), .S1(d3_71__N_562[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1062_11.INIT0 = 16'h74b8;
    defparam add_1062_11.INIT1 = 16'h74b8;
    defparam add_1062_11.INJECT1_0 = "NO";
    defparam add_1062_11.INJECT1_1 = "NO";
    CCU2D add_1062_9 (.A0(d3[42]), .B0(n4603), .C0(n4604[6]), .D0(d2[42]), 
          .A1(d3[43]), .B1(n4603), .C1(n4604[7]), .D1(d2[43]), .CIN(n11881), 
          .COUT(n11882), .S0(d3_71__N_562[42]), .S1(d3_71__N_562[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1062_9.INIT0 = 16'h74b8;
    defparam add_1062_9.INIT1 = 16'h74b8;
    defparam add_1062_9.INJECT1_0 = "NO";
    defparam add_1062_9.INJECT1_1 = "NO";
    CCU2D add_1062_7 (.A0(d3[40]), .B0(n4603), .C0(n4604[4]), .D0(d2[40]), 
          .A1(d3[41]), .B1(n4603), .C1(n4604[5]), .D1(d2[41]), .CIN(n11880), 
          .COUT(n11881), .S0(d3_71__N_562[40]), .S1(d3_71__N_562[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1062_7.INIT0 = 16'h74b8;
    defparam add_1062_7.INIT1 = 16'h74b8;
    defparam add_1062_7.INJECT1_0 = "NO";
    defparam add_1062_7.INJECT1_1 = "NO";
    CCU2D add_1062_5 (.A0(d3[38]), .B0(n4603), .C0(n4604[2]), .D0(d2[38]), 
          .A1(d3[39]), .B1(n4603), .C1(n4604[3]), .D1(d2[39]), .CIN(n11879), 
          .COUT(n11880), .S0(d3_71__N_562[38]), .S1(d3_71__N_562[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1062_5.INIT0 = 16'h74b8;
    defparam add_1062_5.INIT1 = 16'h74b8;
    defparam add_1062_5.INJECT1_0 = "NO";
    defparam add_1062_5.INJECT1_1 = "NO";
    CCU2D add_1062_3 (.A0(d3[36]), .B0(n4603), .C0(n4604[0]), .D0(d2[36]), 
          .A1(d3[37]), .B1(n4603), .C1(n4604[1]), .D1(d2[37]), .CIN(n11878), 
          .COUT(n11879), .S0(d3_71__N_562[36]), .S1(d3_71__N_562[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1062_3.INIT0 = 16'h74b8;
    defparam add_1062_3.INIT1 = 16'h74b8;
    defparam add_1062_3.INJECT1_0 = "NO";
    defparam add_1062_3.INJECT1_1 = "NO";
    CCU2D add_1062_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n4603), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11878));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1062_1.INIT0 = 16'hF000;
    defparam add_1062_1.INIT1 = 16'h0555;
    defparam add_1062_1.INJECT1_0 = "NO";
    defparam add_1062_1.INJECT1_1 = "NO";
    CCU2D add_1066_36 (.A0(d3[70]), .B0(d4[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[71]), .B1(d4[71]), .C1(GND_net), .D1(GND_net), .CIN(n11873), 
          .S0(n4756[34]), .S1(n4756[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1066_36.INIT0 = 16'h5666;
    defparam add_1066_36.INIT1 = 16'h5666;
    defparam add_1066_36.INJECT1_0 = "NO";
    defparam add_1066_36.INJECT1_1 = "NO";
    CCU2D add_1066_34 (.A0(d3[68]), .B0(d4[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[69]), .B1(d4[69]), .C1(GND_net), .D1(GND_net), .CIN(n11872), 
          .COUT(n11873), .S0(n4756[32]), .S1(n4756[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1066_34.INIT0 = 16'h5666;
    defparam add_1066_34.INIT1 = 16'h5666;
    defparam add_1066_34.INJECT1_0 = "NO";
    defparam add_1066_34.INJECT1_1 = "NO";
    CCU2D add_1066_32 (.A0(d3[66]), .B0(d4[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[67]), .B1(d4[67]), .C1(GND_net), .D1(GND_net), .CIN(n11871), 
          .COUT(n11872), .S0(n4756[30]), .S1(n4756[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1066_32.INIT0 = 16'h5666;
    defparam add_1066_32.INIT1 = 16'h5666;
    defparam add_1066_32.INJECT1_0 = "NO";
    defparam add_1066_32.INJECT1_1 = "NO";
    CCU2D add_1066_30 (.A0(d3[64]), .B0(d4[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[65]), .B1(d4[65]), .C1(GND_net), .D1(GND_net), .CIN(n11870), 
          .COUT(n11871), .S0(n4756[28]), .S1(n4756[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1066_30.INIT0 = 16'h5666;
    defparam add_1066_30.INIT1 = 16'h5666;
    defparam add_1066_30.INJECT1_0 = "NO";
    defparam add_1066_30.INJECT1_1 = "NO";
    CCU2D add_1066_28 (.A0(d3[62]), .B0(d4[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[63]), .B1(d4[63]), .C1(GND_net), .D1(GND_net), .CIN(n11869), 
          .COUT(n11870), .S0(n4756[26]), .S1(n4756[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1066_28.INIT0 = 16'h5666;
    defparam add_1066_28.INIT1 = 16'h5666;
    defparam add_1066_28.INJECT1_0 = "NO";
    defparam add_1066_28.INJECT1_1 = "NO";
    CCU2D add_1066_26 (.A0(d3[60]), .B0(d4[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[61]), .B1(d4[61]), .C1(GND_net), .D1(GND_net), .CIN(n11868), 
          .COUT(n11869), .S0(n4756[24]), .S1(n4756[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1066_26.INIT0 = 16'h5666;
    defparam add_1066_26.INIT1 = 16'h5666;
    defparam add_1066_26.INJECT1_0 = "NO";
    defparam add_1066_26.INJECT1_1 = "NO";
    CCU2D add_1066_24 (.A0(d3[58]), .B0(d4[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[59]), .B1(d4[59]), .C1(GND_net), .D1(GND_net), .CIN(n11867), 
          .COUT(n11868), .S0(n4756[22]), .S1(n4756[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1066_24.INIT0 = 16'h5666;
    defparam add_1066_24.INIT1 = 16'h5666;
    defparam add_1066_24.INJECT1_0 = "NO";
    defparam add_1066_24.INJECT1_1 = "NO";
    CCU2D add_1066_22 (.A0(d3[56]), .B0(d4[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[57]), .B1(d4[57]), .C1(GND_net), .D1(GND_net), .CIN(n11866), 
          .COUT(n11867), .S0(n4756[20]), .S1(n4756[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1066_22.INIT0 = 16'h5666;
    defparam add_1066_22.INIT1 = 16'h5666;
    defparam add_1066_22.INJECT1_0 = "NO";
    defparam add_1066_22.INJECT1_1 = "NO";
    CCU2D add_1066_20 (.A0(d3[54]), .B0(d4[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[55]), .B1(d4[55]), .C1(GND_net), .D1(GND_net), .CIN(n11865), 
          .COUT(n11866), .S0(n4756[18]), .S1(n4756[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1066_20.INIT0 = 16'h5666;
    defparam add_1066_20.INIT1 = 16'h5666;
    defparam add_1066_20.INJECT1_0 = "NO";
    defparam add_1066_20.INJECT1_1 = "NO";
    CCU2D add_1066_18 (.A0(d3[52]), .B0(d4[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[53]), .B1(d4[53]), .C1(GND_net), .D1(GND_net), .CIN(n11864), 
          .COUT(n11865), .S0(n4756[16]), .S1(n4756[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1066_18.INIT0 = 16'h5666;
    defparam add_1066_18.INIT1 = 16'h5666;
    defparam add_1066_18.INJECT1_0 = "NO";
    defparam add_1066_18.INJECT1_1 = "NO";
    CCU2D add_1066_16 (.A0(d3[50]), .B0(d4[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[51]), .B1(d4[51]), .C1(GND_net), .D1(GND_net), .CIN(n11863), 
          .COUT(n11864), .S0(n4756[14]), .S1(n4756[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1066_16.INIT0 = 16'h5666;
    defparam add_1066_16.INIT1 = 16'h5666;
    defparam add_1066_16.INJECT1_0 = "NO";
    defparam add_1066_16.INJECT1_1 = "NO";
    CCU2D add_1066_14 (.A0(d3[48]), .B0(d4[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[49]), .B1(d4[49]), .C1(GND_net), .D1(GND_net), .CIN(n11862), 
          .COUT(n11863), .S0(n4756[12]), .S1(n4756[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1066_14.INIT0 = 16'h5666;
    defparam add_1066_14.INIT1 = 16'h5666;
    defparam add_1066_14.INJECT1_0 = "NO";
    defparam add_1066_14.INJECT1_1 = "NO";
    CCU2D add_1066_12 (.A0(d3[46]), .B0(d4[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[47]), .B1(d4[47]), .C1(GND_net), .D1(GND_net), .CIN(n11861), 
          .COUT(n11862), .S0(n4756[10]), .S1(n4756[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1066_12.INIT0 = 16'h5666;
    defparam add_1066_12.INIT1 = 16'h5666;
    defparam add_1066_12.INJECT1_0 = "NO";
    defparam add_1066_12.INJECT1_1 = "NO";
    CCU2D add_1066_10 (.A0(d3[44]), .B0(d4[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[45]), .B1(d4[45]), .C1(GND_net), .D1(GND_net), .CIN(n11860), 
          .COUT(n11861), .S0(n4756[8]), .S1(n4756[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1066_10.INIT0 = 16'h5666;
    defparam add_1066_10.INIT1 = 16'h5666;
    defparam add_1066_10.INJECT1_0 = "NO";
    defparam add_1066_10.INJECT1_1 = "NO";
    CCU2D add_1066_8 (.A0(d3[42]), .B0(d4[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[43]), .B1(d4[43]), .C1(GND_net), .D1(GND_net), .CIN(n11859), 
          .COUT(n11860), .S0(n4756[6]), .S1(n4756[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1066_8.INIT0 = 16'h5666;
    defparam add_1066_8.INIT1 = 16'h5666;
    defparam add_1066_8.INJECT1_0 = "NO";
    defparam add_1066_8.INJECT1_1 = "NO";
    CCU2D add_1066_6 (.A0(d3[40]), .B0(d4[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[41]), .B1(d4[41]), .C1(GND_net), .D1(GND_net), .CIN(n11858), 
          .COUT(n11859), .S0(n4756[4]), .S1(n4756[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1066_6.INIT0 = 16'h5666;
    defparam add_1066_6.INIT1 = 16'h5666;
    defparam add_1066_6.INJECT1_0 = "NO";
    defparam add_1066_6.INJECT1_1 = "NO";
    CCU2D add_1066_4 (.A0(d3[38]), .B0(d4[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[39]), .B1(d4[39]), .C1(GND_net), .D1(GND_net), .CIN(n11857), 
          .COUT(n11858), .S0(n4756[2]), .S1(n4756[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1066_4.INIT0 = 16'h5666;
    defparam add_1066_4.INIT1 = 16'h5666;
    defparam add_1066_4.INJECT1_0 = "NO";
    defparam add_1066_4.INJECT1_1 = "NO";
    CCU2D add_1066_2 (.A0(d3[36]), .B0(d4[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[37]), .B1(d4[37]), .C1(GND_net), .D1(GND_net), .COUT(n11857), 
          .S1(n4756[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1066_2.INIT0 = 16'h7000;
    defparam add_1066_2.INIT1 = 16'h5666;
    defparam add_1066_2.INJECT1_0 = "NO";
    defparam add_1066_2.INJECT1_1 = "NO";
    CCU2D add_1067_37 (.A0(d4[70]), .B0(n4755), .C0(n4756[34]), .D0(d3[70]), 
          .A1(d4[71]), .B1(n4755), .C1(n4756[35]), .D1(d3[71]), .CIN(n11854), 
          .S0(d4_71__N_634[70]), .S1(d4_71__N_634[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1067_37.INIT0 = 16'h74b8;
    defparam add_1067_37.INIT1 = 16'h74b8;
    defparam add_1067_37.INJECT1_0 = "NO";
    defparam add_1067_37.INJECT1_1 = "NO";
    CCU2D add_1067_35 (.A0(d4[68]), .B0(n4755), .C0(n4756[32]), .D0(d3[68]), 
          .A1(d4[69]), .B1(n4755), .C1(n4756[33]), .D1(d3[69]), .CIN(n11853), 
          .COUT(n11854), .S0(d4_71__N_634[68]), .S1(d4_71__N_634[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1067_35.INIT0 = 16'h74b8;
    defparam add_1067_35.INIT1 = 16'h74b8;
    defparam add_1067_35.INJECT1_0 = "NO";
    defparam add_1067_35.INJECT1_1 = "NO";
    CCU2D add_1067_33 (.A0(d4[66]), .B0(n4755), .C0(n4756[30]), .D0(d3[66]), 
          .A1(d4[67]), .B1(n4755), .C1(n4756[31]), .D1(d3[67]), .CIN(n11852), 
          .COUT(n11853), .S0(d4_71__N_634[66]), .S1(d4_71__N_634[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1067_33.INIT0 = 16'h74b8;
    defparam add_1067_33.INIT1 = 16'h74b8;
    defparam add_1067_33.INJECT1_0 = "NO";
    defparam add_1067_33.INJECT1_1 = "NO";
    CCU2D add_1067_31 (.A0(d4[64]), .B0(n4755), .C0(n4756[28]), .D0(d3[64]), 
          .A1(d4[65]), .B1(n4755), .C1(n4756[29]), .D1(d3[65]), .CIN(n11851), 
          .COUT(n11852), .S0(d4_71__N_634[64]), .S1(d4_71__N_634[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1067_31.INIT0 = 16'h74b8;
    defparam add_1067_31.INIT1 = 16'h74b8;
    defparam add_1067_31.INJECT1_0 = "NO";
    defparam add_1067_31.INJECT1_1 = "NO";
    LUT4 i4655_2_lut (.A(d1[36]), .B(d2[36]), .Z(n4452[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4655_2_lut.init = 16'h6666;
    FD1S3AX v_comb_66_rep_105 (.D(osc_clk_enable_141), .CK(osc_clk), .Q(osc_clk_enable_260)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_105.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_35 (.A(n13180), .B(n54), .Z(n8425)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_35.init = 16'hbbbb;
    FD1S3AX v_comb_66_rep_104 (.D(osc_clk_enable_141), .CK(osc_clk), .Q(osc_clk_enable_210)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_104.GSR = "ENABLED";
    LUT4 i11_3_lut_4_lut_then_3_lut (.A(\CICGain[0] ), .B(\d10[67] ), .C(\d10[68] ), 
         .Z(n13075)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam i11_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 i1_2_lut_adj_36 (.A(n375[0]), .B(n54), .Z(count_15__N_1442[0])) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_36.init = 16'hbbbb;
    FD1S3AX v_comb_66_rep_111 (.D(osc_clk_enable_141), .CK(osc_clk), .Q(osc_clk_enable_560)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_111.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_112 (.D(osc_clk_enable_141), .CK(osc_clk), .Q(osc_clk_enable_610)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_112.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_103 (.D(osc_clk_enable_141), .CK(osc_clk), .Q(osc_clk_enable_160)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_103.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_102 (.D(osc_clk_enable_141), .CK(osc_clk), .Q(osc_clk_enable_69)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_102.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_110 (.D(osc_clk_enable_141), .CK(osc_clk), .Q(osc_clk_enable_510)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_110.GSR = "ENABLED";
    CCU2D add_1046_37 (.A0(d_tmp[71]), .B0(d_d_tmp[71]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12037), .S0(n4148[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1046_37.INIT0 = 16'h5999;
    defparam add_1046_37.INIT1 = 16'h0000;
    defparam add_1046_37.INJECT1_0 = "NO";
    defparam add_1046_37.INJECT1_1 = "NO";
    CCU2D add_1067_29 (.A0(d4[62]), .B0(n4755), .C0(n4756[26]), .D0(d3[62]), 
          .A1(d4[63]), .B1(n4755), .C1(n4756[27]), .D1(d3[63]), .CIN(n11850), 
          .COUT(n11851), .S0(d4_71__N_634[62]), .S1(d4_71__N_634[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1067_29.INIT0 = 16'h74b8;
    defparam add_1067_29.INIT1 = 16'h74b8;
    defparam add_1067_29.INJECT1_0 = "NO";
    defparam add_1067_29.INJECT1_1 = "NO";
    LUT4 i11_3_lut_4_lut_else_3_lut (.A(\CICGain[0] ), .B(\d10[69] ), .C(\d10[70] ), 
         .Z(n13074)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam i11_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    CCU2D add_1046_35 (.A0(d_tmp[69]), .B0(d_d_tmp[69]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[70]), .B1(d_d_tmp[70]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12036), .COUT(n12037), .S0(n4148[33]), 
          .S1(n4148[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1046_35.INIT0 = 16'h5999;
    defparam add_1046_35.INIT1 = 16'h5999;
    defparam add_1046_35.INJECT1_0 = "NO";
    defparam add_1046_35.INJECT1_1 = "NO";
    CCU2D add_1046_33 (.A0(d_tmp[67]), .B0(d_d_tmp[67]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[68]), .B1(d_d_tmp[68]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12035), .COUT(n12036), .S0(n4148[31]), 
          .S1(n4148[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1046_33.INIT0 = 16'h5999;
    defparam add_1046_33.INIT1 = 16'h5999;
    defparam add_1046_33.INJECT1_0 = "NO";
    defparam add_1046_33.INJECT1_1 = "NO";
    CCU2D add_1046_31 (.A0(d_tmp[65]), .B0(d_d_tmp[65]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[66]), .B1(d_d_tmp[66]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12034), .COUT(n12035), .S0(n4148[29]), 
          .S1(n4148[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1046_31.INIT0 = 16'h5999;
    defparam add_1046_31.INIT1 = 16'h5999;
    defparam add_1046_31.INJECT1_0 = "NO";
    defparam add_1046_31.INJECT1_1 = "NO";
    CCU2D add_1067_27 (.A0(d4[60]), .B0(n4755), .C0(n4756[24]), .D0(d3[60]), 
          .A1(d4[61]), .B1(n4755), .C1(n4756[25]), .D1(d3[61]), .CIN(n11849), 
          .COUT(n11850), .S0(d4_71__N_634[60]), .S1(d4_71__N_634[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1067_27.INIT0 = 16'h74b8;
    defparam add_1067_27.INIT1 = 16'h74b8;
    defparam add_1067_27.INJECT1_0 = "NO";
    defparam add_1067_27.INJECT1_1 = "NO";
    CCU2D add_1067_25 (.A0(d4[58]), .B0(n4755), .C0(n4756[22]), .D0(d3[58]), 
          .A1(d4[59]), .B1(n4755), .C1(n4756[23]), .D1(d3[59]), .CIN(n11848), 
          .COUT(n11849), .S0(d4_71__N_634[58]), .S1(d4_71__N_634[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1067_25.INIT0 = 16'h74b8;
    defparam add_1067_25.INIT1 = 16'h74b8;
    defparam add_1067_25.INJECT1_0 = "NO";
    defparam add_1067_25.INJECT1_1 = "NO";
    CCU2D add_1046_29 (.A0(d_tmp[63]), .B0(d_d_tmp[63]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[64]), .B1(d_d_tmp[64]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12033), .COUT(n12034), .S0(n4148[27]), 
          .S1(n4148[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1046_29.INIT0 = 16'h5999;
    defparam add_1046_29.INIT1 = 16'h5999;
    defparam add_1046_29.INJECT1_0 = "NO";
    defparam add_1046_29.INJECT1_1 = "NO";
    CCU2D add_1046_27 (.A0(d_tmp[61]), .B0(d_d_tmp[61]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[62]), .B1(d_d_tmp[62]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12032), .COUT(n12033), .S0(n4148[25]), 
          .S1(n4148[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1046_27.INIT0 = 16'h5999;
    defparam add_1046_27.INIT1 = 16'h5999;
    defparam add_1046_27.INJECT1_0 = "NO";
    defparam add_1046_27.INJECT1_1 = "NO";
    CCU2D add_1046_25 (.A0(d_tmp[59]), .B0(d_d_tmp[59]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[60]), .B1(d_d_tmp[60]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12031), .COUT(n12032), .S0(n4148[23]), 
          .S1(n4148[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1046_25.INIT0 = 16'h5999;
    defparam add_1046_25.INIT1 = 16'h5999;
    defparam add_1046_25.INJECT1_0 = "NO";
    defparam add_1046_25.INJECT1_1 = "NO";
    CCU2D add_1067_23 (.A0(d4[56]), .B0(n4755), .C0(n4756[20]), .D0(d3[56]), 
          .A1(d4[57]), .B1(n4755), .C1(n4756[21]), .D1(d3[57]), .CIN(n11847), 
          .COUT(n11848), .S0(d4_71__N_634[56]), .S1(d4_71__N_634[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1067_23.INIT0 = 16'h74b8;
    defparam add_1067_23.INIT1 = 16'h74b8;
    defparam add_1067_23.INJECT1_0 = "NO";
    defparam add_1067_23.INJECT1_1 = "NO";
    CCU2D add_1046_23 (.A0(d_tmp[57]), .B0(d_d_tmp[57]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[58]), .B1(d_d_tmp[58]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12030), .COUT(n12031), .S0(n4148[21]), 
          .S1(n4148[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1046_23.INIT0 = 16'h5999;
    defparam add_1046_23.INIT1 = 16'h5999;
    defparam add_1046_23.INJECT1_0 = "NO";
    defparam add_1046_23.INJECT1_1 = "NO";
    CCU2D add_1046_21 (.A0(d_tmp[55]), .B0(d_d_tmp[55]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[56]), .B1(d_d_tmp[56]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12029), .COUT(n12030), .S0(n4148[19]), 
          .S1(n4148[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1046_21.INIT0 = 16'h5999;
    defparam add_1046_21.INIT1 = 16'h5999;
    defparam add_1046_21.INJECT1_0 = "NO";
    defparam add_1046_21.INJECT1_1 = "NO";
    CCU2D add_1046_19 (.A0(d_tmp[53]), .B0(d_d_tmp[53]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[54]), .B1(d_d_tmp[54]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12028), .COUT(n12029), .S0(n4148[17]), 
          .S1(n4148[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1046_19.INIT0 = 16'h5999;
    defparam add_1046_19.INIT1 = 16'h5999;
    defparam add_1046_19.INJECT1_0 = "NO";
    defparam add_1046_19.INJECT1_1 = "NO";
    CCU2D add_1067_21 (.A0(d4[54]), .B0(n4755), .C0(n4756[18]), .D0(d3[54]), 
          .A1(d4[55]), .B1(n4755), .C1(n4756[19]), .D1(d3[55]), .CIN(n11846), 
          .COUT(n11847), .S0(d4_71__N_634[54]), .S1(d4_71__N_634[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1067_21.INIT0 = 16'h74b8;
    defparam add_1067_21.INIT1 = 16'h74b8;
    defparam add_1067_21.INJECT1_0 = "NO";
    defparam add_1067_21.INJECT1_1 = "NO";
    CCU2D add_1067_19 (.A0(d4[52]), .B0(n4755), .C0(n4756[16]), .D0(d3[52]), 
          .A1(d4[53]), .B1(n4755), .C1(n4756[17]), .D1(d3[53]), .CIN(n11845), 
          .COUT(n11846), .S0(d4_71__N_634[52]), .S1(d4_71__N_634[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1067_19.INIT0 = 16'h74b8;
    defparam add_1067_19.INIT1 = 16'h74b8;
    defparam add_1067_19.INJECT1_0 = "NO";
    defparam add_1067_19.INJECT1_1 = "NO";
    CCU2D add_1046_17 (.A0(d_tmp[51]), .B0(d_d_tmp[51]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[52]), .B1(d_d_tmp[52]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12027), .COUT(n12028), .S0(n4148[15]), 
          .S1(n4148[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1046_17.INIT0 = 16'h5999;
    defparam add_1046_17.INIT1 = 16'h5999;
    defparam add_1046_17.INJECT1_0 = "NO";
    defparam add_1046_17.INJECT1_1 = "NO";
    CCU2D add_1046_15 (.A0(d_tmp[49]), .B0(d_d_tmp[49]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[50]), .B1(d_d_tmp[50]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12026), .COUT(n12027), .S0(n4148[13]), 
          .S1(n4148[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1046_15.INIT0 = 16'h5999;
    defparam add_1046_15.INIT1 = 16'h5999;
    defparam add_1046_15.INJECT1_0 = "NO";
    defparam add_1046_15.INJECT1_1 = "NO";
    CCU2D add_1046_13 (.A0(d_tmp[47]), .B0(d_d_tmp[47]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[48]), .B1(d_d_tmp[48]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12025), .COUT(n12026), .S0(n4148[11]), 
          .S1(n4148[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1046_13.INIT0 = 16'h5999;
    defparam add_1046_13.INIT1 = 16'h5999;
    defparam add_1046_13.INJECT1_0 = "NO";
    defparam add_1046_13.INJECT1_1 = "NO";
    CCU2D add_1067_17 (.A0(d4[50]), .B0(n4755), .C0(n4756[14]), .D0(d3[50]), 
          .A1(d4[51]), .B1(n4755), .C1(n4756[15]), .D1(d3[51]), .CIN(n11844), 
          .COUT(n11845), .S0(d4_71__N_634[50]), .S1(d4_71__N_634[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1067_17.INIT0 = 16'h74b8;
    defparam add_1067_17.INIT1 = 16'h74b8;
    defparam add_1067_17.INJECT1_0 = "NO";
    defparam add_1067_17.INJECT1_1 = "NO";
    CCU2D add_1046_11 (.A0(d_tmp[45]), .B0(d_d_tmp[45]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[46]), .B1(d_d_tmp[46]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12024), .COUT(n12025), .S0(n4148[9]), 
          .S1(n4148[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1046_11.INIT0 = 16'h5999;
    defparam add_1046_11.INIT1 = 16'h5999;
    defparam add_1046_11.INJECT1_0 = "NO";
    defparam add_1046_11.INJECT1_1 = "NO";
    CCU2D add_1046_9 (.A0(d_tmp[43]), .B0(d_d_tmp[43]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[44]), .B1(d_d_tmp[44]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12023), .COUT(n12024), .S0(n4148[7]), 
          .S1(n4148[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1046_9.INIT0 = 16'h5999;
    defparam add_1046_9.INIT1 = 16'h5999;
    defparam add_1046_9.INJECT1_0 = "NO";
    defparam add_1046_9.INJECT1_1 = "NO";
    CCU2D add_1046_7 (.A0(d_tmp[41]), .B0(d_d_tmp[41]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[42]), .B1(d_d_tmp[42]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12022), .COUT(n12023), .S0(n4148[5]), 
          .S1(n4148[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1046_7.INIT0 = 16'h5999;
    defparam add_1046_7.INIT1 = 16'h5999;
    defparam add_1046_7.INJECT1_0 = "NO";
    defparam add_1046_7.INJECT1_1 = "NO";
    CCU2D add_1067_15 (.A0(d4[48]), .B0(n4755), .C0(n4756[12]), .D0(d3[48]), 
          .A1(d4[49]), .B1(n4755), .C1(n4756[13]), .D1(d3[49]), .CIN(n11843), 
          .COUT(n11844), .S0(d4_71__N_634[48]), .S1(d4_71__N_634[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1067_15.INIT0 = 16'h74b8;
    defparam add_1067_15.INIT1 = 16'h74b8;
    defparam add_1067_15.INJECT1_0 = "NO";
    defparam add_1067_15.INJECT1_1 = "NO";
    CCU2D add_1067_13 (.A0(d4[46]), .B0(n4755), .C0(n4756[10]), .D0(d3[46]), 
          .A1(d4[47]), .B1(n4755), .C1(n4756[11]), .D1(d3[47]), .CIN(n11842), 
          .COUT(n11843), .S0(d4_71__N_634[46]), .S1(d4_71__N_634[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1067_13.INIT0 = 16'h74b8;
    defparam add_1067_13.INIT1 = 16'h74b8;
    defparam add_1067_13.INJECT1_0 = "NO";
    defparam add_1067_13.INJECT1_1 = "NO";
    CCU2D add_1046_5 (.A0(d_tmp[39]), .B0(d_d_tmp[39]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[40]), .B1(d_d_tmp[40]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12021), .COUT(n12022), .S0(n4148[3]), 
          .S1(n4148[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1046_5.INIT0 = 16'h5999;
    defparam add_1046_5.INIT1 = 16'h5999;
    defparam add_1046_5.INJECT1_0 = "NO";
    defparam add_1046_5.INJECT1_1 = "NO";
    CCU2D add_1046_3 (.A0(d_tmp[37]), .B0(d_d_tmp[37]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[38]), .B1(d_d_tmp[38]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12020), .COUT(n12021), .S0(n4148[1]), 
          .S1(n4148[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1046_3.INIT0 = 16'h5999;
    defparam add_1046_3.INIT1 = 16'h5999;
    defparam add_1046_3.INJECT1_0 = "NO";
    defparam add_1046_3.INJECT1_1 = "NO";
    CCU2D add_1046_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[36]), .B1(d_d_tmp[36]), .C1(GND_net), .D1(GND_net), 
          .COUT(n12020), .S1(n4148[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1046_1.INIT0 = 16'hF000;
    defparam add_1046_1.INIT1 = 16'h5999;
    defparam add_1046_1.INJECT1_0 = "NO";
    defparam add_1046_1.INJECT1_1 = "NO";
    CCU2D add_1047_37 (.A0(d_d_tmp[70]), .B0(n4147), .C0(n4148[34]), .D0(d_tmp[70]), 
          .A1(d_d_tmp[71]), .B1(n4147), .C1(n4148[35]), .D1(d_tmp[71]), 
          .CIN(n12018), .S0(d6_71__N_1459[70]), .S1(d6_71__N_1459[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1047_37.INIT0 = 16'hb874;
    defparam add_1047_37.INIT1 = 16'hb874;
    defparam add_1047_37.INJECT1_0 = "NO";
    defparam add_1047_37.INJECT1_1 = "NO";
    CCU2D add_1047_35 (.A0(d_d_tmp[68]), .B0(n4147), .C0(n4148[32]), .D0(d_tmp[68]), 
          .A1(d_d_tmp[69]), .B1(n4147), .C1(n4148[33]), .D1(d_tmp[69]), 
          .CIN(n12017), .COUT(n12018), .S0(d6_71__N_1459[68]), .S1(d6_71__N_1459[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1047_35.INIT0 = 16'hb874;
    defparam add_1047_35.INIT1 = 16'hb874;
    defparam add_1047_35.INJECT1_0 = "NO";
    defparam add_1047_35.INJECT1_1 = "NO";
    LUT4 i13_4_lut_rep_99 (.A(n21_adj_2495), .B(n26), .C(n15), .D(n16), 
         .Z(n13180)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i13_4_lut_rep_99.init = 16'h8000;
    CCU2D add_1047_33 (.A0(d_d_tmp[66]), .B0(n4147), .C0(n4148[30]), .D0(d_tmp[66]), 
          .A1(d_d_tmp[67]), .B1(n4147), .C1(n4148[31]), .D1(d_tmp[67]), 
          .CIN(n12016), .COUT(n12017), .S0(d6_71__N_1459[66]), .S1(d6_71__N_1459[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1047_33.INIT0 = 16'hb874;
    defparam add_1047_33.INIT1 = 16'hb874;
    defparam add_1047_33.INJECT1_0 = "NO";
    defparam add_1047_33.INJECT1_1 = "NO";
    CCU2D add_1047_31 (.A0(d_d_tmp[64]), .B0(n4147), .C0(n4148[28]), .D0(d_tmp[64]), 
          .A1(d_d_tmp[65]), .B1(n4147), .C1(n4148[29]), .D1(d_tmp[65]), 
          .CIN(n12015), .COUT(n12016), .S0(d6_71__N_1459[64]), .S1(d6_71__N_1459[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1047_31.INIT0 = 16'hb874;
    defparam add_1047_31.INIT1 = 16'hb874;
    defparam add_1047_31.INJECT1_0 = "NO";
    defparam add_1047_31.INJECT1_1 = "NO";
    CCU2D add_1047_29 (.A0(d_d_tmp[62]), .B0(n4147), .C0(n4148[26]), .D0(d_tmp[62]), 
          .A1(d_d_tmp[63]), .B1(n4147), .C1(n4148[27]), .D1(d_tmp[63]), 
          .CIN(n12014), .COUT(n12015), .S0(d6_71__N_1459[62]), .S1(d6_71__N_1459[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1047_29.INIT0 = 16'hb874;
    defparam add_1047_29.INIT1 = 16'hb874;
    defparam add_1047_29.INJECT1_0 = "NO";
    defparam add_1047_29.INJECT1_1 = "NO";
    CCU2D add_1047_27 (.A0(d_d_tmp[60]), .B0(n4147), .C0(n4148[24]), .D0(d_tmp[60]), 
          .A1(d_d_tmp[61]), .B1(n4147), .C1(n4148[25]), .D1(d_tmp[61]), 
          .CIN(n12013), .COUT(n12014), .S0(d6_71__N_1459[60]), .S1(d6_71__N_1459[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1047_27.INIT0 = 16'hb874;
    defparam add_1047_27.INIT1 = 16'hb874;
    defparam add_1047_27.INJECT1_0 = "NO";
    defparam add_1047_27.INJECT1_1 = "NO";
    CCU2D add_1047_25 (.A0(d_d_tmp[58]), .B0(n4147), .C0(n4148[22]), .D0(d_tmp[58]), 
          .A1(d_d_tmp[59]), .B1(n4147), .C1(n4148[23]), .D1(d_tmp[59]), 
          .CIN(n12012), .COUT(n12013), .S0(d6_71__N_1459[58]), .S1(d6_71__N_1459[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1047_25.INIT0 = 16'hb874;
    defparam add_1047_25.INIT1 = 16'hb874;
    defparam add_1047_25.INJECT1_0 = "NO";
    defparam add_1047_25.INJECT1_1 = "NO";
    CCU2D add_1047_23 (.A0(d_d_tmp[56]), .B0(n4147), .C0(n4148[20]), .D0(d_tmp[56]), 
          .A1(d_d_tmp[57]), .B1(n4147), .C1(n4148[21]), .D1(d_tmp[57]), 
          .CIN(n12011), .COUT(n12012), .S0(d6_71__N_1459[56]), .S1(d6_71__N_1459[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1047_23.INIT0 = 16'hb874;
    defparam add_1047_23.INIT1 = 16'hb874;
    defparam add_1047_23.INJECT1_0 = "NO";
    defparam add_1047_23.INJECT1_1 = "NO";
    CCU2D add_1047_21 (.A0(d_d_tmp[54]), .B0(n4147), .C0(n4148[18]), .D0(d_tmp[54]), 
          .A1(d_d_tmp[55]), .B1(n4147), .C1(n4148[19]), .D1(d_tmp[55]), 
          .CIN(n12010), .COUT(n12011), .S0(d6_71__N_1459[54]), .S1(d6_71__N_1459[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1047_21.INIT0 = 16'hb874;
    defparam add_1047_21.INIT1 = 16'hb874;
    defparam add_1047_21.INJECT1_0 = "NO";
    defparam add_1047_21.INJECT1_1 = "NO";
    CCU2D add_1047_19 (.A0(d_d_tmp[52]), .B0(n4147), .C0(n4148[16]), .D0(d_tmp[52]), 
          .A1(d_d_tmp[53]), .B1(n4147), .C1(n4148[17]), .D1(d_tmp[53]), 
          .CIN(n12009), .COUT(n12010), .S0(d6_71__N_1459[52]), .S1(d6_71__N_1459[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1047_19.INIT0 = 16'hb874;
    defparam add_1047_19.INIT1 = 16'hb874;
    defparam add_1047_19.INJECT1_0 = "NO";
    defparam add_1047_19.INJECT1_1 = "NO";
    CCU2D add_1047_17 (.A0(d_d_tmp[50]), .B0(n4147), .C0(n4148[14]), .D0(d_tmp[50]), 
          .A1(d_d_tmp[51]), .B1(n4147), .C1(n4148[15]), .D1(d_tmp[51]), 
          .CIN(n12008), .COUT(n12009), .S0(d6_71__N_1459[50]), .S1(d6_71__N_1459[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1047_17.INIT0 = 16'hb874;
    defparam add_1047_17.INIT1 = 16'hb874;
    defparam add_1047_17.INJECT1_0 = "NO";
    defparam add_1047_17.INJECT1_1 = "NO";
    CCU2D add_1047_15 (.A0(d_d_tmp[48]), .B0(n4147), .C0(n4148[12]), .D0(d_tmp[48]), 
          .A1(d_d_tmp[49]), .B1(n4147), .C1(n4148[13]), .D1(d_tmp[49]), 
          .CIN(n12007), .COUT(n12008), .S0(d6_71__N_1459[48]), .S1(d6_71__N_1459[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1047_15.INIT0 = 16'hb874;
    defparam add_1047_15.INIT1 = 16'hb874;
    defparam add_1047_15.INJECT1_0 = "NO";
    defparam add_1047_15.INJECT1_1 = "NO";
    CCU2D add_1047_13 (.A0(d_d_tmp[46]), .B0(n4147), .C0(n4148[10]), .D0(d_tmp[46]), 
          .A1(d_d_tmp[47]), .B1(n4147), .C1(n4148[11]), .D1(d_tmp[47]), 
          .CIN(n12006), .COUT(n12007), .S0(d6_71__N_1459[46]), .S1(d6_71__N_1459[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1047_13.INIT0 = 16'hb874;
    defparam add_1047_13.INIT1 = 16'hb874;
    defparam add_1047_13.INJECT1_0 = "NO";
    defparam add_1047_13.INJECT1_1 = "NO";
    CCU2D add_1047_11 (.A0(d_d_tmp[44]), .B0(n4147), .C0(n4148[8]), .D0(d_tmp[44]), 
          .A1(d_d_tmp[45]), .B1(n4147), .C1(n4148[9]), .D1(d_tmp[45]), 
          .CIN(n12005), .COUT(n12006), .S0(d6_71__N_1459[44]), .S1(d6_71__N_1459[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1047_11.INIT0 = 16'hb874;
    defparam add_1047_11.INIT1 = 16'hb874;
    defparam add_1047_11.INJECT1_0 = "NO";
    defparam add_1047_11.INJECT1_1 = "NO";
    CCU2D add_1067_11 (.A0(d4[44]), .B0(n4755), .C0(n4756[8]), .D0(d3[44]), 
          .A1(d4[45]), .B1(n4755), .C1(n4756[9]), .D1(d3[45]), .CIN(n11841), 
          .COUT(n11842), .S0(d4_71__N_634[44]), .S1(d4_71__N_634[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1067_11.INIT0 = 16'h74b8;
    defparam add_1067_11.INIT1 = 16'h74b8;
    defparam add_1067_11.INJECT1_0 = "NO";
    defparam add_1067_11.INJECT1_1 = "NO";
    CCU2D add_1047_9 (.A0(d_d_tmp[42]), .B0(n4147), .C0(n4148[6]), .D0(d_tmp[42]), 
          .A1(d_d_tmp[43]), .B1(n4147), .C1(n4148[7]), .D1(d_tmp[43]), 
          .CIN(n12004), .COUT(n12005), .S0(d6_71__N_1459[42]), .S1(d6_71__N_1459[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1047_9.INIT0 = 16'hb874;
    defparam add_1047_9.INIT1 = 16'hb874;
    defparam add_1047_9.INJECT1_0 = "NO";
    defparam add_1047_9.INJECT1_1 = "NO";
    CCU2D add_1047_7 (.A0(d_d_tmp[40]), .B0(n4147), .C0(n4148[4]), .D0(d_tmp[40]), 
          .A1(d_d_tmp[41]), .B1(n4147), .C1(n4148[5]), .D1(d_tmp[41]), 
          .CIN(n12003), .COUT(n12004), .S0(d6_71__N_1459[40]), .S1(d6_71__N_1459[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1047_7.INIT0 = 16'hb874;
    defparam add_1047_7.INIT1 = 16'hb874;
    defparam add_1047_7.INJECT1_0 = "NO";
    defparam add_1047_7.INJECT1_1 = "NO";
    CCU2D add_1047_5 (.A0(d_d_tmp[38]), .B0(n4147), .C0(n4148[2]), .D0(d_tmp[38]), 
          .A1(d_d_tmp[39]), .B1(n4147), .C1(n4148[3]), .D1(d_tmp[39]), 
          .CIN(n12002), .COUT(n12003), .S0(d6_71__N_1459[38]), .S1(d6_71__N_1459[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1047_5.INIT0 = 16'hb874;
    defparam add_1047_5.INIT1 = 16'hb874;
    defparam add_1047_5.INJECT1_0 = "NO";
    defparam add_1047_5.INJECT1_1 = "NO";
    CCU2D add_1047_3 (.A0(d_d_tmp[36]), .B0(n4147), .C0(n4148[0]), .D0(d_tmp[36]), 
          .A1(d_d_tmp[37]), .B1(n4147), .C1(n4148[1]), .D1(d_tmp[37]), 
          .CIN(n12001), .COUT(n12002), .S0(d6_71__N_1459[36]), .S1(d6_71__N_1459[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1047_3.INIT0 = 16'hb874;
    defparam add_1047_3.INIT1 = 16'hb874;
    defparam add_1047_3.INJECT1_0 = "NO";
    defparam add_1047_3.INJECT1_1 = "NO";
    CCU2D add_1047_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n4147), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n12001));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1047_1.INIT0 = 16'hF000;
    defparam add_1047_1.INIT1 = 16'h0555;
    defparam add_1047_1.INJECT1_0 = "NO";
    defparam add_1047_1.INJECT1_1 = "NO";
    CCU2D add_1051_36 (.A0(MixerOutSin[11]), .B0(d1[70]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[71]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11996), .S0(n4300[34]), .S1(n4300[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1051_36.INIT0 = 16'h5666;
    defparam add_1051_36.INIT1 = 16'h5666;
    defparam add_1051_36.INJECT1_0 = "NO";
    defparam add_1051_36.INJECT1_1 = "NO";
    CCU2D add_1067_9 (.A0(d4[42]), .B0(n4755), .C0(n4756[6]), .D0(d3[42]), 
          .A1(d4[43]), .B1(n4755), .C1(n4756[7]), .D1(d3[43]), .CIN(n11840), 
          .COUT(n11841), .S0(d4_71__N_634[42]), .S1(d4_71__N_634[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1067_9.INIT0 = 16'h74b8;
    defparam add_1067_9.INIT1 = 16'h74b8;
    defparam add_1067_9.INJECT1_0 = "NO";
    defparam add_1067_9.INJECT1_1 = "NO";
    CCU2D add_1051_34 (.A0(MixerOutSin[11]), .B0(d1[68]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[69]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11995), .COUT(n11996), .S0(n4300[32]), 
          .S1(n4300[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1051_34.INIT0 = 16'h5666;
    defparam add_1051_34.INIT1 = 16'h5666;
    defparam add_1051_34.INJECT1_0 = "NO";
    defparam add_1051_34.INJECT1_1 = "NO";
    CCU2D add_1051_32 (.A0(MixerOutSin[11]), .B0(d1[66]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[67]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11994), .COUT(n11995), .S0(n4300[30]), 
          .S1(n4300[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1051_32.INIT0 = 16'h5666;
    defparam add_1051_32.INIT1 = 16'h5666;
    defparam add_1051_32.INJECT1_0 = "NO";
    defparam add_1051_32.INJECT1_1 = "NO";
    CCU2D add_1051_30 (.A0(MixerOutSin[11]), .B0(d1[64]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[65]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11993), .COUT(n11994), .S0(n4300[28]), 
          .S1(n4300[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1051_30.INIT0 = 16'h5666;
    defparam add_1051_30.INIT1 = 16'h5666;
    defparam add_1051_30.INJECT1_0 = "NO";
    defparam add_1051_30.INJECT1_1 = "NO";
    CCU2D add_1051_28 (.A0(MixerOutSin[11]), .B0(d1[62]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[63]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11992), .COUT(n11993), .S0(n4300[26]), 
          .S1(n4300[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1051_28.INIT0 = 16'h5666;
    defparam add_1051_28.INIT1 = 16'h5666;
    defparam add_1051_28.INJECT1_0 = "NO";
    defparam add_1051_28.INJECT1_1 = "NO";
    CCU2D add_1051_26 (.A0(MixerOutSin[11]), .B0(d1[60]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[61]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11991), .COUT(n11992), .S0(n4300[24]), 
          .S1(n4300[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1051_26.INIT0 = 16'h5666;
    defparam add_1051_26.INIT1 = 16'h5666;
    defparam add_1051_26.INJECT1_0 = "NO";
    defparam add_1051_26.INJECT1_1 = "NO";
    CCU2D add_1067_7 (.A0(d4[40]), .B0(n4755), .C0(n4756[4]), .D0(d3[40]), 
          .A1(d4[41]), .B1(n4755), .C1(n4756[5]), .D1(d3[41]), .CIN(n11839), 
          .COUT(n11840), .S0(d4_71__N_634[40]), .S1(d4_71__N_634[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1067_7.INIT0 = 16'h74b8;
    defparam add_1067_7.INIT1 = 16'h74b8;
    defparam add_1067_7.INJECT1_0 = "NO";
    defparam add_1067_7.INJECT1_1 = "NO";
    CCU2D add_1051_24 (.A0(MixerOutSin[11]), .B0(d1[58]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[59]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11990), .COUT(n11991), .S0(n4300[22]), 
          .S1(n4300[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1051_24.INIT0 = 16'h5666;
    defparam add_1051_24.INIT1 = 16'h5666;
    defparam add_1051_24.INJECT1_0 = "NO";
    defparam add_1051_24.INJECT1_1 = "NO";
    CCU2D add_1051_22 (.A0(MixerOutSin[11]), .B0(d1[56]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[57]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11989), .COUT(n11990), .S0(n4300[20]), 
          .S1(n4300[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1051_22.INIT0 = 16'h5666;
    defparam add_1051_22.INIT1 = 16'h5666;
    defparam add_1051_22.INJECT1_0 = "NO";
    defparam add_1051_22.INJECT1_1 = "NO";
    CCU2D add_1051_20 (.A0(MixerOutSin[11]), .B0(d1[54]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[55]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11988), .COUT(n11989), .S0(n4300[18]), 
          .S1(n4300[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1051_20.INIT0 = 16'h5666;
    defparam add_1051_20.INIT1 = 16'h5666;
    defparam add_1051_20.INJECT1_0 = "NO";
    defparam add_1051_20.INJECT1_1 = "NO";
    CCU2D add_1051_18 (.A0(MixerOutSin[11]), .B0(d1[52]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[53]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11987), .COUT(n11988), .S0(n4300[16]), 
          .S1(n4300[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1051_18.INIT0 = 16'h5666;
    defparam add_1051_18.INIT1 = 16'h5666;
    defparam add_1051_18.INJECT1_0 = "NO";
    defparam add_1051_18.INJECT1_1 = "NO";
    LUT4 i11_3_lut_4_lut_else_3_lut_adj_37 (.A(\CICGain[0] ), .B(d10[69]), 
         .C(d10[70]), .Z(n13077)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam i11_3_lut_4_lut_else_3_lut_adj_37.init = 16'hd8d8;
    CCU2D add_1106_9 (.A0(d9[43]), .B0(d_d9[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[44]), .B1(d_d9[44]), .C1(GND_net), .D1(GND_net), .CIN(n11533), 
          .COUT(n11534));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1106_9.INIT0 = 16'h5999;
    defparam add_1106_9.INIT1 = 16'h5999;
    defparam add_1106_9.INJECT1_0 = "NO";
    defparam add_1106_9.INJECT1_1 = "NO";
    LUT4 mux_1244_i2_3_lut (.A(n5972[21]), .B(n6010[21]), .C(n5971), .Z(d10_71__N_1747[57])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1244_i2_3_lut.init = 16'hcaca;
    CCU2D add_1106_29 (.A0(d9[63]), .B0(d_d9[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[64]), .B1(d_d9[64]), .C1(GND_net), .D1(GND_net), .CIN(n11543), 
          .COUT(n11544), .S0(n5972[27]), .S1(n5972[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1106_29.INIT0 = 16'h5999;
    defparam add_1106_29.INIT1 = 16'h5999;
    defparam add_1106_29.INJECT1_0 = "NO";
    defparam add_1106_29.INJECT1_1 = "NO";
    LUT4 mux_1244_i3_3_lut (.A(n5972[22]), .B(n6010[22]), .C(n5971), .Z(d10_71__N_1747[58])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1244_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1244_i4_3_lut (.A(n5972[23]), .B(n6010[23]), .C(n5971), .Z(d10_71__N_1747[59])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1244_i4_3_lut.init = 16'hcaca;
    FD1S3AX v_comb_66_rep_114 (.D(osc_clk_enable_141), .CK(osc_clk), .Q(osc_clk_enable_710)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_114.GSR = "ENABLED";
    CCU2D add_1106_25 (.A0(d9[59]), .B0(d_d9[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[60]), .B1(d_d9[60]), .C1(GND_net), .D1(GND_net), .CIN(n11541), 
          .COUT(n11542), .S0(n5972[23]), .S1(n5972[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1106_25.INIT0 = 16'h5999;
    defparam add_1106_25.INIT1 = 16'h5999;
    defparam add_1106_25.INJECT1_0 = "NO";
    defparam add_1106_25.INJECT1_1 = "NO";
    LUT4 i5418_then_3_lut (.A(\CICGain[1] ), .B(d10[59]), .C(d10[57]), 
         .Z(n13081)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i5418_then_3_lut.init = 16'he4e4;
    CCU2D add_1106_27 (.A0(d9[61]), .B0(d_d9[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[62]), .B1(d_d9[62]), .C1(GND_net), .D1(GND_net), .CIN(n11542), 
          .COUT(n11543), .S0(n5972[25]), .S1(n5972[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1106_27.INIT0 = 16'h5999;
    defparam add_1106_27.INIT1 = 16'h5999;
    defparam add_1106_27.INJECT1_0 = "NO";
    defparam add_1106_27.INJECT1_1 = "NO";
    LUT4 i5418_else_3_lut (.A(n61_c), .B(\CICGain[1] ), .C(d10[58]), .Z(n13080)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i5418_else_3_lut.init = 16'he2e2;
    CCU2D add_1051_16 (.A0(MixerOutSin[11]), .B0(d1[50]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[51]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11986), .COUT(n11987), .S0(n4300[14]), 
          .S1(n4300[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1051_16.INIT0 = 16'h5666;
    defparam add_1051_16.INIT1 = 16'h5666;
    defparam add_1051_16.INJECT1_0 = "NO";
    defparam add_1051_16.INJECT1_1 = "NO";
    CCU2D add_1051_14 (.A0(MixerOutSin[11]), .B0(d1[48]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[49]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11985), .COUT(n11986), .S0(n4300[12]), 
          .S1(n4300[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1051_14.INIT0 = 16'h5666;
    defparam add_1051_14.INIT1 = 16'h5666;
    defparam add_1051_14.INJECT1_0 = "NO";
    defparam add_1051_14.INJECT1_1 = "NO";
    CCU2D add_1051_12 (.A0(MixerOutSin[11]), .B0(d1[46]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[47]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11984), .COUT(n11985), .S0(n4300[10]), 
          .S1(n4300[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1051_12.INIT0 = 16'h5666;
    defparam add_1051_12.INIT1 = 16'h5666;
    defparam add_1051_12.INJECT1_0 = "NO";
    defparam add_1051_12.INJECT1_1 = "NO";
    CCU2D add_1051_10 (.A0(MixerOutSin[11]), .B0(d1[44]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[45]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11983), .COUT(n11984), .S0(n4300[8]), 
          .S1(n4300[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1051_10.INIT0 = 16'h5666;
    defparam add_1051_10.INIT1 = 16'h5666;
    defparam add_1051_10.INJECT1_0 = "NO";
    defparam add_1051_10.INJECT1_1 = "NO";
    CCU2D add_1051_8 (.A0(MixerOutSin[11]), .B0(d1[42]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[43]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11982), .COUT(n11983), .S0(n4300[6]), 
          .S1(n4300[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1051_8.INIT0 = 16'h5666;
    defparam add_1051_8.INIT1 = 16'h5666;
    defparam add_1051_8.INJECT1_0 = "NO";
    defparam add_1051_8.INJECT1_1 = "NO";
    CCU2D add_1051_6 (.A0(MixerOutSin[11]), .B0(d1[40]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[41]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11981), .COUT(n11982), .S0(n4300[4]), 
          .S1(n4300[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1051_6.INIT0 = 16'h5666;
    defparam add_1051_6.INIT1 = 16'h5666;
    defparam add_1051_6.INJECT1_0 = "NO";
    defparam add_1051_6.INJECT1_1 = "NO";
    CCU2D add_1051_4 (.A0(MixerOutSin[11]), .B0(d1[38]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[39]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11980), .COUT(n11981), .S0(n4300[2]), 
          .S1(n4300[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1051_4.INIT0 = 16'h5666;
    defparam add_1051_4.INIT1 = 16'h5666;
    defparam add_1051_4.INJECT1_0 = "NO";
    defparam add_1051_4.INJECT1_1 = "NO";
    CCU2D add_1051_2 (.A0(MixerOutSin[11]), .B0(d1[36]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[37]), .C1(GND_net), 
          .D1(GND_net), .COUT(n11980), .S1(n4300[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1051_2.INIT0 = 16'h7000;
    defparam add_1051_2.INIT1 = 16'h5666;
    defparam add_1051_2.INJECT1_0 = "NO";
    defparam add_1051_2.INJECT1_1 = "NO";
    CCU2D add_1067_5 (.A0(d4[38]), .B0(n4755), .C0(n4756[2]), .D0(d3[38]), 
          .A1(d4[39]), .B1(n4755), .C1(n4756[3]), .D1(d3[39]), .CIN(n11838), 
          .COUT(n11839), .S0(d4_71__N_634[38]), .S1(d4_71__N_634[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1067_5.INIT0 = 16'h74b8;
    defparam add_1067_5.INIT1 = 16'h74b8;
    defparam add_1067_5.INJECT1_0 = "NO";
    defparam add_1067_5.INJECT1_1 = "NO";
    LUT4 mux_1244_i5_3_lut (.A(n5972[24]), .B(n6010[24]), .C(n5971), .Z(d10_71__N_1747[60])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1244_i5_3_lut.init = 16'hcaca;
    LUT4 i5428_then_3_lut (.A(\CICGain[1] ), .B(d10[60]), .C(d10[58]), 
         .Z(n13084)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i5428_then_3_lut.init = 16'he4e4;
    CCU2D add_1067_3 (.A0(d4[36]), .B0(n4755), .C0(n4756[0]), .D0(d3[36]), 
          .A1(d4[37]), .B1(n4755), .C1(n4756[1]), .D1(d3[37]), .CIN(n11837), 
          .COUT(n11838), .S0(d4_71__N_634[36]), .S1(d4_71__N_634[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1067_3.INIT0 = 16'h74b8;
    defparam add_1067_3.INIT1 = 16'h74b8;
    defparam add_1067_3.INJECT1_0 = "NO";
    defparam add_1067_3.INJECT1_1 = "NO";
    LUT4 mux_1244_i6_3_lut (.A(n5972[25]), .B(n6010[25]), .C(n5971), .Z(d10_71__N_1747[61])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1244_i6_3_lut.init = 16'hcaca;
    LUT4 i5428_else_3_lut (.A(n62_c), .B(\CICGain[1] ), .C(d10[59]), .Z(n13083)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i5428_else_3_lut.init = 16'he2e2;
    CCU2D add_1067_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n4755), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11837));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1067_1.INIT0 = 16'hF000;
    defparam add_1067_1.INIT1 = 16'h0555;
    defparam add_1067_1.INJECT1_0 = "NO";
    defparam add_1067_1.INJECT1_1 = "NO";
    LUT4 mux_1244_i7_3_lut (.A(n5972[26]), .B(n6010[26]), .C(n5971), .Z(d10_71__N_1747[62])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1244_i7_3_lut.init = 16'hcaca;
    LUT4 i4597_2_lut (.A(d1[0]), .B(d2[0]), .Z(d2_71__N_490[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4597_2_lut.init = 16'h6666;
    LUT4 i4598_2_lut (.A(d2[0]), .B(d3[0]), .Z(d3_71__N_562[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4598_2_lut.init = 16'h6666;
    LUT4 i4599_2_lut (.A(d3[0]), .B(d4[0]), .Z(d4_71__N_634[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4599_2_lut.init = 16'h6666;
    LUT4 mux_1244_i8_3_lut (.A(n5972[27]), .B(n6010[27]), .C(n5971), .Z(d10_71__N_1747[63])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1244_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1244_i9_3_lut (.A(n5972[28]), .B(n6010[28]), .C(n5971), .Z(d10_71__N_1747[64])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1244_i9_3_lut.init = 16'hcaca;
    CCU2D add_1071_36 (.A0(d4[70]), .B0(d5[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[71]), .B1(d5[71]), .C1(GND_net), .D1(GND_net), .CIN(n11832), 
          .S0(n4908[34]), .S1(n4908[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1071_36.INIT0 = 16'h5666;
    defparam add_1071_36.INIT1 = 16'h5666;
    defparam add_1071_36.INJECT1_0 = "NO";
    defparam add_1071_36.INJECT1_1 = "NO";
    LUT4 shift_right_31_i138_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n68_c), .D(d10[66]), .Z(n138)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i138_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i67_3_lut_rep_97 (.A(d10[66]), .B(d10[67]), .C(\CICGain[0] ), 
         .Z(n13176)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i67_3_lut_rep_97.init = 16'hcaca;
    LUT4 shift_right_31_i137_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n13176), .D(d10[65]), .Z(n137)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i137_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i133_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63_c), .D(d10[61]), .Z(n133)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i133_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i136_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66_c), .D(d10[64]), .Z(n136)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i136_3_lut_4_lut.init = 16'hf960;
    LUT4 i11_3_lut_4_lut_then_3_lut_3_lut (.A(d10[67]), .B(\CICGain[0] ), 
         .C(d10[68]), .Z(n13078)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam i11_3_lut_4_lut_then_3_lut_3_lut.init = 16'hb8b8;
    LUT4 mux_1244_i10_3_lut (.A(n5972[29]), .B(n6010[29]), .C(n5971), 
         .Z(d10_71__N_1747[65])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1244_i10_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i132_3_lut_4_lut_adj_38 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n62_c), .D(d10[60]), .Z(n132_adj_2488)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i132_3_lut_4_lut_adj_38.init = 16'hf960;
    CCU2D add_1071_34 (.A0(d4[68]), .B0(d5[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[69]), .B1(d5[69]), .C1(GND_net), .D1(GND_net), .CIN(n11831), 
          .COUT(n11832), .S0(n4908[32]), .S1(n4908[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1071_34.INIT0 = 16'h5666;
    defparam add_1071_34.INIT1 = 16'h5666;
    defparam add_1071_34.INJECT1_0 = "NO";
    defparam add_1071_34.INJECT1_1 = "NO";
    LUT4 i13_4_lut_rep_100 (.A(n21_adj_2495), .B(n26), .C(n15), .D(n16), 
         .Z(osc_clk_enable_141)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i13_4_lut_rep_100.init = 16'h8000;
    PFUMX i5440 (.BLUT(n13083), .ALUT(n13084), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[1]));
    LUT4 shift_right_31_i140_3_lut_4_lut_adj_39 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n70), .D(\d10[68] ), .Z(n140_adj_2514)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i140_3_lut_4_lut_adj_39.init = 16'hf960;
    CCU2D add_1071_32 (.A0(d4[66]), .B0(d5[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[67]), .B1(d5[67]), .C1(GND_net), .D1(GND_net), .CIN(n11830), 
          .COUT(n11831), .S0(n4908[30]), .S1(n4908[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1071_32.INIT0 = 16'h5666;
    defparam add_1071_32.INIT1 = 16'h5666;
    defparam add_1071_32.INJECT1_0 = "NO";
    defparam add_1071_32.INJECT1_1 = "NO";
    LUT4 i4600_2_lut (.A(d4[0]), .B(d5[0]), .Z(d5_71__N_706[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4600_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_adj_40 (.A(n54), .B(d_clk_tmp), .Z(n8403)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(50[14:19])
    defparam i1_2_lut_adj_40.init = 16'h8888;
    LUT4 shift_right_31_i137_3_lut_4_lut_adj_41 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n67), .D(\d10[65] ), .Z(n137_adj_2507)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i137_3_lut_4_lut_adj_41.init = 16'hf960;
    CCU2D add_1071_30 (.A0(d4[64]), .B0(d5[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[65]), .B1(d5[65]), .C1(GND_net), .D1(GND_net), .CIN(n11829), 
          .COUT(n11830), .S0(n4908[28]), .S1(n4908[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1071_30.INIT0 = 16'h5666;
    defparam add_1071_30.INIT1 = 16'h5666;
    defparam add_1071_30.INJECT1_0 = "NO";
    defparam add_1071_30.INJECT1_1 = "NO";
    CCU2D add_1071_28 (.A0(d4[62]), .B0(d5[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[63]), .B1(d5[63]), .C1(GND_net), .D1(GND_net), .CIN(n11828), 
          .COUT(n11829), .S0(n4908[26]), .S1(n4908[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1071_28.INIT0 = 16'h5666;
    defparam add_1071_28.INIT1 = 16'h5666;
    defparam add_1071_28.INJECT1_0 = "NO";
    defparam add_1071_28.INJECT1_1 = "NO";
    CCU2D add_1071_26 (.A0(d4[60]), .B0(d5[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[61]), .B1(d5[61]), .C1(GND_net), .D1(GND_net), .CIN(n11827), 
          .COUT(n11828), .S0(n4908[24]), .S1(n4908[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1071_26.INIT0 = 16'h5666;
    defparam add_1071_26.INIT1 = 16'h5666;
    defparam add_1071_26.INJECT1_0 = "NO";
    defparam add_1071_26.INJECT1_1 = "NO";
    CCU2D add_1071_24 (.A0(d4[58]), .B0(d5[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[59]), .B1(d5[59]), .C1(GND_net), .D1(GND_net), .CIN(n11826), 
          .COUT(n11827), .S0(n4908[22]), .S1(n4908[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1071_24.INIT0 = 16'h5666;
    defparam add_1071_24.INIT1 = 16'h5666;
    defparam add_1071_24.INJECT1_0 = "NO";
    defparam add_1071_24.INJECT1_1 = "NO";
    CCU2D add_1071_22 (.A0(d4[56]), .B0(d5[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[57]), .B1(d5[57]), .C1(GND_net), .D1(GND_net), .CIN(n11825), 
          .COUT(n11826), .S0(n4908[20]), .S1(n4908[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1071_22.INIT0 = 16'h5666;
    defparam add_1071_22.INIT1 = 16'h5666;
    defparam add_1071_22.INJECT1_0 = "NO";
    defparam add_1071_22.INJECT1_1 = "NO";
    CCU2D add_1071_20 (.A0(d4[54]), .B0(d5[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[55]), .B1(d5[55]), .C1(GND_net), .D1(GND_net), .CIN(n11824), 
          .COUT(n11825), .S0(n4908[18]), .S1(n4908[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1071_20.INIT0 = 16'h5666;
    defparam add_1071_20.INIT1 = 16'h5666;
    defparam add_1071_20.INJECT1_0 = "NO";
    defparam add_1071_20.INJECT1_1 = "NO";
    PFUMX i5438 (.BLUT(n13080), .ALUT(n13081), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[0]));
    CCU2D add_1071_18 (.A0(d4[52]), .B0(d5[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[53]), .B1(d5[53]), .C1(GND_net), .D1(GND_net), .CIN(n11823), 
          .COUT(n11824), .S0(n4908[16]), .S1(n4908[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1071_18.INIT0 = 16'h5666;
    defparam add_1071_18.INIT1 = 16'h5666;
    defparam add_1071_18.INJECT1_0 = "NO";
    defparam add_1071_18.INJECT1_1 = "NO";
    CCU2D add_1071_16 (.A0(d4[50]), .B0(d5[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[51]), .B1(d5[51]), .C1(GND_net), .D1(GND_net), .CIN(n11822), 
          .COUT(n11823), .S0(n4908[14]), .S1(n4908[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1071_16.INIT0 = 16'h5666;
    defparam add_1071_16.INIT1 = 16'h5666;
    defparam add_1071_16.INJECT1_0 = "NO";
    defparam add_1071_16.INJECT1_1 = "NO";
    LUT4 i13_4_lut_adj_42 (.A(n25), .B(n23), .C(n19), .D(n20), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_42.init = 16'hfffe;
    CCU2D add_1071_14 (.A0(d4[48]), .B0(d5[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[49]), .B1(d5[49]), .C1(GND_net), .D1(GND_net), .CIN(n11821), 
          .COUT(n11822), .S0(n4908[12]), .S1(n4908[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1071_14.INIT0 = 16'h5666;
    defparam add_1071_14.INIT1 = 16'h5666;
    defparam add_1071_14.INJECT1_0 = "NO";
    defparam add_1071_14.INJECT1_1 = "NO";
    CCU2D add_1071_12 (.A0(d4[46]), .B0(d5[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[47]), .B1(d5[47]), .C1(GND_net), .D1(GND_net), .CIN(n11820), 
          .COUT(n11821), .S0(n4908[10]), .S1(n4908[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1071_12.INIT0 = 16'h5666;
    defparam add_1071_12.INIT1 = 16'h5666;
    defparam add_1071_12.INJECT1_0 = "NO";
    defparam add_1071_12.INJECT1_1 = "NO";
    LUT4 i11_4_lut (.A(n21), .B(count[8]), .C(n16_adj_2489), .D(count[3]), 
         .Z(n25)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i11_4_lut.init = 16'hfffe;
    CCU2D add_1071_10 (.A0(d4[44]), .B0(d5[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[45]), .B1(d5[45]), .C1(GND_net), .D1(GND_net), .CIN(n11819), 
          .COUT(n11820), .S0(n4908[8]), .S1(n4908[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1071_10.INIT0 = 16'h5666;
    defparam add_1071_10.INIT1 = 16'h5666;
    defparam add_1071_10.INJECT1_0 = "NO";
    defparam add_1071_10.INJECT1_1 = "NO";
    CCU2D add_1071_8 (.A0(d4[42]), .B0(d5[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[43]), .B1(d5[43]), .C1(GND_net), .D1(GND_net), .CIN(n11818), 
          .COUT(n11819), .S0(n4908[6]), .S1(n4908[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1071_8.INIT0 = 16'h5666;
    defparam add_1071_8.INIT1 = 16'h5666;
    defparam add_1071_8.INJECT1_0 = "NO";
    defparam add_1071_8.INJECT1_1 = "NO";
    LUT4 shift_right_31_i138_3_lut_4_lut_adj_43 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n68), .D(\d10[66] ), .Z(n138_adj_2511)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i138_3_lut_4_lut_adj_43.init = 16'hf960;
    CCU2D add_1071_6 (.A0(d4[40]), .B0(d5[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[41]), .B1(d5[41]), .C1(GND_net), .D1(GND_net), .CIN(n11817), 
          .COUT(n11818), .S0(n4908[4]), .S1(n4908[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1071_6.INIT0 = 16'h5666;
    defparam add_1071_6.INIT1 = 16'h5666;
    defparam add_1071_6.INJECT1_0 = "NO";
    defparam add_1071_6.INJECT1_1 = "NO";
    CCU2D add_1071_4 (.A0(d4[38]), .B0(d5[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[39]), .B1(d5[39]), .C1(GND_net), .D1(GND_net), .CIN(n11816), 
          .COUT(n11817), .S0(n4908[2]), .S1(n4908[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1071_4.INIT0 = 16'h5666;
    defparam add_1071_4.INIT1 = 16'h5666;
    defparam add_1071_4.INJECT1_0 = "NO";
    defparam add_1071_4.INJECT1_1 = "NO";
    PFUMX i5436 (.BLUT(n13077), .ALUT(n13078), .C0(\CICGain[1] ), .Z(d_out_11__N_1819[10]));
    CCU2D add_1071_2 (.A0(d4[36]), .B0(d5[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[37]), .B1(d5[37]), .C1(GND_net), .D1(GND_net), .COUT(n11816), 
          .S1(n4908[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1071_2.INIT0 = 16'h7000;
    defparam add_1071_2.INIT1 = 16'h5666;
    defparam add_1071_2.INJECT1_0 = "NO";
    defparam add_1071_2.INJECT1_1 = "NO";
    LUT4 mux_1244_i11_3_lut (.A(n5972[30]), .B(n6010[30]), .C(n5971), 
         .Z(d10_71__N_1747[66])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1244_i11_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i135_3_lut_4_lut_adj_44 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65), .D(\d10[63] ), .Z(n135_adj_2502)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i135_3_lut_4_lut_adj_44.init = 16'hf960;
    LUT4 mux_1244_i12_3_lut (.A(n5972[31]), .B(n6010[31]), .C(n5971), 
         .Z(d10_71__N_1747[67])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1244_i12_3_lut.init = 16'hcaca;
    CCU2D add_1072_37 (.A0(d5[70]), .B0(n4907), .C0(n4908[34]), .D0(d4[70]), 
          .A1(d5[71]), .B1(n4907), .C1(n4908[35]), .D1(d4[71]), .CIN(n11813), 
          .S0(d5_71__N_706[70]), .S1(d5_71__N_706[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1072_37.INIT0 = 16'h74b8;
    defparam add_1072_37.INIT1 = 16'h74b8;
    defparam add_1072_37.INJECT1_0 = "NO";
    defparam add_1072_37.INJECT1_1 = "NO";
    LUT4 mux_1244_i13_3_lut (.A(n5972[32]), .B(n6010[32]), .C(n5971), 
         .Z(d10_71__N_1747[68])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1244_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1244_i14_3_lut (.A(n5972[33]), .B(n6010[33]), .C(n5971), 
         .Z(d10_71__N_1747[69])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1244_i14_3_lut.init = 16'hcaca;
    CCU2D add_1072_35 (.A0(d5[68]), .B0(n4907), .C0(n4908[32]), .D0(d4[68]), 
          .A1(d5[69]), .B1(n4907), .C1(n4908[33]), .D1(d4[69]), .CIN(n11812), 
          .COUT(n11813), .S0(d5_71__N_706[68]), .S1(d5_71__N_706[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1072_35.INIT0 = 16'h74b8;
    defparam add_1072_35.INIT1 = 16'h74b8;
    defparam add_1072_35.INJECT1_0 = "NO";
    defparam add_1072_35.INJECT1_1 = "NO";
    CCU2D add_1072_33 (.A0(d5[66]), .B0(n4907), .C0(n4908[30]), .D0(d4[66]), 
          .A1(d5[67]), .B1(n4907), .C1(n4908[31]), .D1(d4[67]), .CIN(n11811), 
          .COUT(n11812), .S0(d5_71__N_706[66]), .S1(d5_71__N_706[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1072_33.INIT0 = 16'h74b8;
    defparam add_1072_33.INIT1 = 16'h74b8;
    defparam add_1072_33.INJECT1_0 = "NO";
    defparam add_1072_33.INJECT1_1 = "NO";
    CCU2D add_1052_37 (.A0(d1[70]), .B0(n4299), .C0(n4300[34]), .D0(MixerOutSin[11]), 
          .A1(d1[71]), .B1(n4299), .C1(n4300[35]), .D1(MixerOutSin[11]), 
          .CIN(n11977), .S0(d1_71__N_418[70]), .S1(d1_71__N_418[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1052_37.INIT0 = 16'h74b8;
    defparam add_1052_37.INIT1 = 16'h74b8;
    defparam add_1052_37.INJECT1_0 = "NO";
    defparam add_1052_37.INJECT1_1 = "NO";
    PFUMX i5434 (.BLUT(n13074), .ALUT(n13075), .C0(\CICGain[1] ), .Z(\d_out_11__N_1819[10] ));
    LUT4 shift_right_31_i136_3_lut_4_lut_adj_45 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66), .D(\d10[64] ), .Z(n136_adj_2505)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i136_3_lut_4_lut_adj_45.init = 16'hf960;
    CCU2D add_1072_31 (.A0(d5[64]), .B0(n4907), .C0(n4908[28]), .D0(d4[64]), 
          .A1(d5[65]), .B1(n4907), .C1(n4908[29]), .D1(d4[65]), .CIN(n11810), 
          .COUT(n11811), .S0(d5_71__N_706[64]), .S1(d5_71__N_706[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1072_31.INIT0 = 16'h74b8;
    defparam add_1072_31.INIT1 = 16'h74b8;
    defparam add_1072_31.INJECT1_0 = "NO";
    defparam add_1072_31.INJECT1_1 = "NO";
    CCU2D add_1072_29 (.A0(d5[62]), .B0(n4907), .C0(n4908[26]), .D0(d4[62]), 
          .A1(d5[63]), .B1(n4907), .C1(n4908[27]), .D1(d4[63]), .CIN(n11809), 
          .COUT(n11810), .S0(d5_71__N_706[62]), .S1(d5_71__N_706[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1072_29.INIT0 = 16'h74b8;
    defparam add_1072_29.INIT1 = 16'h74b8;
    defparam add_1072_29.INJECT1_0 = "NO";
    defparam add_1072_29.INJECT1_1 = "NO";
    CCU2D add_1052_35 (.A0(d1[68]), .B0(n4299), .C0(n4300[32]), .D0(MixerOutSin[11]), 
          .A1(d1[69]), .B1(n4299), .C1(n4300[33]), .D1(MixerOutSin[11]), 
          .CIN(n11976), .COUT(n11977), .S0(d1_71__N_418[68]), .S1(d1_71__N_418[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1052_35.INIT0 = 16'h74b8;
    defparam add_1052_35.INIT1 = 16'h74b8;
    defparam add_1052_35.INJECT1_0 = "NO";
    defparam add_1052_35.INJECT1_1 = "NO";
    CCU2D add_1052_33 (.A0(d1[66]), .B0(n4299), .C0(n4300[30]), .D0(MixerOutSin[11]), 
          .A1(d1[67]), .B1(n4299), .C1(n4300[31]), .D1(MixerOutSin[11]), 
          .CIN(n11975), .COUT(n11976), .S0(d1_71__N_418[66]), .S1(d1_71__N_418[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1052_33.INIT0 = 16'h74b8;
    defparam add_1052_33.INIT1 = 16'h74b8;
    defparam add_1052_33.INJECT1_0 = "NO";
    defparam add_1052_33.INJECT1_1 = "NO";
    LUT4 mux_1244_i15_3_lut (.A(n5972[34]), .B(n6010[34]), .C(n5971), 
         .Z(d10_71__N_1747[70])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1244_i15_3_lut.init = 16'hcaca;
    CCU2D add_1072_27 (.A0(d5[60]), .B0(n4907), .C0(n4908[24]), .D0(d4[60]), 
          .A1(d5[61]), .B1(n4907), .C1(n4908[25]), .D1(d4[61]), .CIN(n11808), 
          .COUT(n11809), .S0(d5_71__N_706[60]), .S1(d5_71__N_706[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1072_27.INIT0 = 16'h74b8;
    defparam add_1072_27.INIT1 = 16'h74b8;
    defparam add_1072_27.INJECT1_0 = "NO";
    defparam add_1072_27.INJECT1_1 = "NO";
    CCU2D add_1072_25 (.A0(d5[58]), .B0(n4907), .C0(n4908[22]), .D0(d4[58]), 
          .A1(d5[59]), .B1(n4907), .C1(n4908[23]), .D1(d4[59]), .CIN(n11807), 
          .COUT(n11808), .S0(d5_71__N_706[58]), .S1(d5_71__N_706[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1072_25.INIT0 = 16'h74b8;
    defparam add_1072_25.INIT1 = 16'h74b8;
    defparam add_1072_25.INJECT1_0 = "NO";
    defparam add_1072_25.INJECT1_1 = "NO";
    CCU2D add_1072_23 (.A0(d5[56]), .B0(n4907), .C0(n4908[20]), .D0(d4[56]), 
          .A1(d5[57]), .B1(n4907), .C1(n4908[21]), .D1(d4[57]), .CIN(n11806), 
          .COUT(n11807), .S0(d5_71__N_706[56]), .S1(d5_71__N_706[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1072_23.INIT0 = 16'h74b8;
    defparam add_1072_23.INIT1 = 16'h74b8;
    defparam add_1072_23.INJECT1_0 = "NO";
    defparam add_1072_23.INJECT1_1 = "NO";
    CCU2D add_1072_21 (.A0(d5[54]), .B0(n4907), .C0(n4908[18]), .D0(d4[54]), 
          .A1(d5[55]), .B1(n4907), .C1(n4908[19]), .D1(d4[55]), .CIN(n11805), 
          .COUT(n11806), .S0(d5_71__N_706[54]), .S1(d5_71__N_706[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1072_21.INIT0 = 16'h74b8;
    defparam add_1072_21.INIT1 = 16'h74b8;
    defparam add_1072_21.INJECT1_0 = "NO";
    defparam add_1072_21.INJECT1_1 = "NO";
    CCU2D add_1072_19 (.A0(d5[52]), .B0(n4907), .C0(n4908[16]), .D0(d4[52]), 
          .A1(d5[53]), .B1(n4907), .C1(n4908[17]), .D1(d4[53]), .CIN(n11804), 
          .COUT(n11805), .S0(d5_71__N_706[52]), .S1(d5_71__N_706[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1072_19.INIT0 = 16'h74b8;
    defparam add_1072_19.INIT1 = 16'h74b8;
    defparam add_1072_19.INJECT1_0 = "NO";
    defparam add_1072_19.INJECT1_1 = "NO";
    CCU2D add_1072_17 (.A0(d5[50]), .B0(n4907), .C0(n4908[14]), .D0(d4[50]), 
          .A1(d5[51]), .B1(n4907), .C1(n4908[15]), .D1(d4[51]), .CIN(n11803), 
          .COUT(n11804), .S0(d5_71__N_706[50]), .S1(d5_71__N_706[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1072_17.INIT0 = 16'h74b8;
    defparam add_1072_17.INIT1 = 16'h74b8;
    defparam add_1072_17.INJECT1_0 = "NO";
    defparam add_1072_17.INJECT1_1 = "NO";
    CCU2D add_1072_15 (.A0(d5[48]), .B0(n4907), .C0(n4908[12]), .D0(d4[48]), 
          .A1(d5[49]), .B1(n4907), .C1(n4908[13]), .D1(d4[49]), .CIN(n11802), 
          .COUT(n11803), .S0(d5_71__N_706[48]), .S1(d5_71__N_706[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1072_15.INIT0 = 16'h74b8;
    defparam add_1072_15.INIT1 = 16'h74b8;
    defparam add_1072_15.INJECT1_0 = "NO";
    defparam add_1072_15.INJECT1_1 = "NO";
    CCU2D add_1072_13 (.A0(d5[46]), .B0(n4907), .C0(n4908[10]), .D0(d4[46]), 
          .A1(d5[47]), .B1(n4907), .C1(n4908[11]), .D1(d4[47]), .CIN(n11801), 
          .COUT(n11802), .S0(d5_71__N_706[46]), .S1(d5_71__N_706[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1072_13.INIT0 = 16'h74b8;
    defparam add_1072_13.INIT1 = 16'h74b8;
    defparam add_1072_13.INJECT1_0 = "NO";
    defparam add_1072_13.INJECT1_1 = "NO";
    CCU2D add_1072_11 (.A0(d5[44]), .B0(n4907), .C0(n4908[8]), .D0(d4[44]), 
          .A1(d5[45]), .B1(n4907), .C1(n4908[9]), .D1(d4[45]), .CIN(n11800), 
          .COUT(n11801), .S0(d5_71__N_706[44]), .S1(d5_71__N_706[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1072_11.INIT0 = 16'h74b8;
    defparam add_1072_11.INIT1 = 16'h74b8;
    defparam add_1072_11.INJECT1_0 = "NO";
    defparam add_1072_11.INJECT1_1 = "NO";
    LUT4 mux_1244_i16_3_lut (.A(n5972[35]), .B(n6010[35]), .C(n5971), 
         .Z(d10_71__N_1747[71])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1244_i16_3_lut.init = 16'hcaca;
    CCU2D add_1072_9 (.A0(d5[42]), .B0(n4907), .C0(n4908[6]), .D0(d4[42]), 
          .A1(d5[43]), .B1(n4907), .C1(n4908[7]), .D1(d4[43]), .CIN(n11799), 
          .COUT(n11800), .S0(d5_71__N_706[42]), .S1(d5_71__N_706[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1072_9.INIT0 = 16'h74b8;
    defparam add_1072_9.INIT1 = 16'h74b8;
    defparam add_1072_9.INJECT1_0 = "NO";
    defparam add_1072_9.INJECT1_1 = "NO";
    LUT4 shift_right_31_i133_3_lut_4_lut_adj_46 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63), .D(\d10[61] ), .Z(n133_adj_2497)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i133_3_lut_4_lut_adj_46.init = 16'hf960;
    CCU2D add_1072_7 (.A0(d5[40]), .B0(n4907), .C0(n4908[4]), .D0(d4[40]), 
          .A1(d5[41]), .B1(n4907), .C1(n4908[5]), .D1(d4[41]), .CIN(n11798), 
          .COUT(n11799), .S0(d5_71__N_706[40]), .S1(d5_71__N_706[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1072_7.INIT0 = 16'h74b8;
    defparam add_1072_7.INIT1 = 16'h74b8;
    defparam add_1072_7.INJECT1_0 = "NO";
    defparam add_1072_7.INJECT1_1 = "NO";
    CCU2D add_1072_5 (.A0(d5[38]), .B0(n4907), .C0(n4908[2]), .D0(d4[38]), 
          .A1(d5[39]), .B1(n4907), .C1(n4908[3]), .D1(d4[39]), .CIN(n11797), 
          .COUT(n11798), .S0(d5_71__N_706[38]), .S1(d5_71__N_706[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1072_5.INIT0 = 16'h74b8;
    defparam add_1072_5.INIT1 = 16'h74b8;
    defparam add_1072_5.INJECT1_0 = "NO";
    defparam add_1072_5.INJECT1_1 = "NO";
    FD1S3AX v_comb_66_rep_107 (.D(osc_clk_enable_141), .CK(osc_clk), .Q(osc_clk_enable_360)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=171, LSE_RLINE=177 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_107.GSR = "ENABLED";
    CCU2D add_1072_3 (.A0(d5[36]), .B0(n4907), .C0(n4908[0]), .D0(d4[36]), 
          .A1(d5[37]), .B1(n4907), .C1(n4908[1]), .D1(d4[37]), .CIN(n11796), 
          .COUT(n11797), .S0(d5_71__N_706[36]), .S1(d5_71__N_706[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1072_3.INIT0 = 16'h74b8;
    defparam add_1072_3.INIT1 = 16'h74b8;
    defparam add_1072_3.INJECT1_0 = "NO";
    defparam add_1072_3.INJECT1_1 = "NO";
    CCU2D add_1072_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n4907), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11796));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1072_1.INIT0 = 16'hF000;
    defparam add_1072_1.INIT1 = 16'h0555;
    defparam add_1072_1.INJECT1_0 = "NO";
    defparam add_1072_1.INJECT1_1 = "NO";
    CCU2D add_1052_31 (.A0(d1[64]), .B0(n4299), .C0(n4300[28]), .D0(MixerOutSin[11]), 
          .A1(d1[65]), .B1(n4299), .C1(n4300[29]), .D1(MixerOutSin[11]), 
          .CIN(n11974), .COUT(n11975), .S0(d1_71__N_418[64]), .S1(d1_71__N_418[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1052_31.INIT0 = 16'h74b8;
    defparam add_1052_31.INIT1 = 16'h74b8;
    defparam add_1052_31.INJECT1_0 = "NO";
    defparam add_1052_31.INJECT1_1 = "NO";
    CCU2D add_1052_29 (.A0(d1[62]), .B0(n4299), .C0(n4300[26]), .D0(MixerOutSin[11]), 
          .A1(d1[63]), .B1(n4299), .C1(n4300[27]), .D1(MixerOutSin[11]), 
          .CIN(n11973), .COUT(n11974), .S0(d1_71__N_418[62]), .S1(d1_71__N_418[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1052_29.INIT0 = 16'h74b8;
    defparam add_1052_29.INIT1 = 16'h74b8;
    defparam add_1052_29.INJECT1_0 = "NO";
    defparam add_1052_29.INJECT1_1 = "NO";
    CCU2D add_1052_27 (.A0(d1[60]), .B0(n4299), .C0(n4300[24]), .D0(MixerOutSin[11]), 
          .A1(d1[61]), .B1(n4299), .C1(n4300[25]), .D1(MixerOutSin[11]), 
          .CIN(n11972), .COUT(n11973), .S0(d1_71__N_418[60]), .S1(d1_71__N_418[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1052_27.INIT0 = 16'h74b8;
    defparam add_1052_27.INIT1 = 16'h74b8;
    defparam add_1052_27.INJECT1_0 = "NO";
    defparam add_1052_27.INJECT1_1 = "NO";
    CCU2D add_1052_25 (.A0(d1[58]), .B0(n4299), .C0(n4300[22]), .D0(MixerOutSin[11]), 
          .A1(d1[59]), .B1(n4299), .C1(n4300[23]), .D1(MixerOutSin[11]), 
          .CIN(n11971), .COUT(n11972), .S0(d1_71__N_418[58]), .S1(d1_71__N_418[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1052_25.INIT0 = 16'h74b8;
    defparam add_1052_25.INIT1 = 16'h74b8;
    defparam add_1052_25.INJECT1_0 = "NO";
    defparam add_1052_25.INJECT1_1 = "NO";
    CCU2D add_1052_23 (.A0(d1[56]), .B0(n4299), .C0(n4300[20]), .D0(MixerOutSin[11]), 
          .A1(d1[57]), .B1(n4299), .C1(n4300[21]), .D1(MixerOutSin[11]), 
          .CIN(n11970), .COUT(n11971), .S0(d1_71__N_418[56]), .S1(d1_71__N_418[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1052_23.INIT0 = 16'h74b8;
    defparam add_1052_23.INIT1 = 16'h74b8;
    defparam add_1052_23.INJECT1_0 = "NO";
    defparam add_1052_23.INJECT1_1 = "NO";
    LUT4 shift_right_31_i134_3_lut_4_lut_adj_47 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64), .D(\d10[62] ), .Z(n134_adj_2500)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i134_3_lut_4_lut_adj_47.init = 16'hf960;
    CCU2D add_1052_21 (.A0(d1[54]), .B0(n4299), .C0(n4300[18]), .D0(MixerOutSin[11]), 
          .A1(d1[55]), .B1(n4299), .C1(n4300[19]), .D1(MixerOutSin[11]), 
          .CIN(n11969), .COUT(n11970), .S0(d1_71__N_418[54]), .S1(d1_71__N_418[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1052_21.INIT0 = 16'h74b8;
    defparam add_1052_21.INIT1 = 16'h74b8;
    defparam add_1052_21.INJECT1_0 = "NO";
    defparam add_1052_21.INJECT1_1 = "NO";
    LUT4 shift_right_31_i131_3_lut_4_lut_adj_48 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n61), .D(\d10[59] ), .Z(n131_adj_2491)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i131_3_lut_4_lut_adj_48.init = 16'hf960;
    CCU2D add_1052_19 (.A0(d1[52]), .B0(n4299), .C0(n4300[16]), .D0(MixerOutSin[11]), 
          .A1(d1[53]), .B1(n4299), .C1(n4300[17]), .D1(MixerOutSin[11]), 
          .CIN(n11968), .COUT(n11969), .S0(d1_71__N_418[52]), .S1(d1_71__N_418[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1052_19.INIT0 = 16'h74b8;
    defparam add_1052_19.INIT1 = 16'h74b8;
    defparam add_1052_19.INJECT1_0 = "NO";
    defparam add_1052_19.INJECT1_1 = "NO";
    CCU2D add_1052_17 (.A0(d1[50]), .B0(n4299), .C0(n4300[14]), .D0(MixerOutSin[11]), 
          .A1(d1[51]), .B1(n4299), .C1(n4300[15]), .D1(MixerOutSin[11]), 
          .CIN(n11967), .COUT(n11968), .S0(d1_71__N_418[50]), .S1(d1_71__N_418[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1052_17.INIT0 = 16'h74b8;
    defparam add_1052_17.INIT1 = 16'h74b8;
    defparam add_1052_17.INJECT1_0 = "NO";
    defparam add_1052_17.INJECT1_1 = "NO";
    CCU2D add_1052_15 (.A0(d1[48]), .B0(n4299), .C0(n4300[12]), .D0(MixerOutSin[11]), 
          .A1(d1[49]), .B1(n4299), .C1(n4300[13]), .D1(MixerOutSin[11]), 
          .CIN(n11966), .COUT(n11967), .S0(d1_71__N_418[48]), .S1(d1_71__N_418[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1052_15.INIT0 = 16'h74b8;
    defparam add_1052_15.INIT1 = 16'h74b8;
    defparam add_1052_15.INJECT1_0 = "NO";
    defparam add_1052_15.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module nco_sig
//

module nco_sig (osc_clk, \phase_accum[56] , \phase_accum[57] , \phase_accum[58] , 
            \phase_accum[59] , \phase_accum[60] , \phase_accum[61] , \phase_accum[62] , 
            \phase_accum[63] , phase_inc_carrGen1, GND_net, sinGen_c) /* synthesis syn_module_defined=1 */ ;
    input osc_clk;
    output \phase_accum[56] ;
    output \phase_accum[57] ;
    output \phase_accum[58] ;
    output \phase_accum[59] ;
    output \phase_accum[60] ;
    output \phase_accum[61] ;
    output \phase_accum[62] ;
    output \phase_accum[63] ;
    input [63:0]phase_inc_carrGen1;
    input GND_net;
    output sinGen_c;
    
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(69[8:15])
    wire [63:0]phase_accum;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(29[19:30])
    wire [63:0]phase_accum_63__N_146;
    
    wire n10692, n10691, n10690, n10689, n10688, n10687, n10686, 
        n10685, n10684, n10683, n10682, n10681, n10680, n10679, 
        n10678, n10677, n10676, n10675, n10674, n10673, n10672, 
        n10671, n10670, n10669, n10668, n10667, n10666, n10665, 
        n10664, n10663, n10662;
    
    FD1S3AX phase_accum_i0 (.D(phase_accum_63__N_146[0]), .CK(osc_clk), 
            .Q(phase_accum[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i0.GSR = "ENABLED";
    FD1S3AX phase_accum_i1 (.D(phase_accum_63__N_146[1]), .CK(osc_clk), 
            .Q(phase_accum[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i1.GSR = "ENABLED";
    FD1S3AX phase_accum_i2 (.D(phase_accum_63__N_146[2]), .CK(osc_clk), 
            .Q(phase_accum[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i2.GSR = "ENABLED";
    FD1S3AX phase_accum_i3 (.D(phase_accum_63__N_146[3]), .CK(osc_clk), 
            .Q(phase_accum[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i3.GSR = "ENABLED";
    FD1S3AX phase_accum_i4 (.D(phase_accum_63__N_146[4]), .CK(osc_clk), 
            .Q(phase_accum[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i4.GSR = "ENABLED";
    FD1S3AX phase_accum_i5 (.D(phase_accum_63__N_146[5]), .CK(osc_clk), 
            .Q(phase_accum[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i5.GSR = "ENABLED";
    FD1S3AX phase_accum_i6 (.D(phase_accum_63__N_146[6]), .CK(osc_clk), 
            .Q(phase_accum[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i6.GSR = "ENABLED";
    FD1S3AX phase_accum_i7 (.D(phase_accum_63__N_146[7]), .CK(osc_clk), 
            .Q(phase_accum[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i7.GSR = "ENABLED";
    FD1S3AX phase_accum_i8 (.D(phase_accum_63__N_146[8]), .CK(osc_clk), 
            .Q(phase_accum[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i8.GSR = "ENABLED";
    FD1S3AX phase_accum_i9 (.D(phase_accum_63__N_146[9]), .CK(osc_clk), 
            .Q(phase_accum[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i9.GSR = "ENABLED";
    FD1S3AX phase_accum_i10 (.D(phase_accum_63__N_146[10]), .CK(osc_clk), 
            .Q(phase_accum[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i10.GSR = "ENABLED";
    FD1S3AX phase_accum_i11 (.D(phase_accum_63__N_146[11]), .CK(osc_clk), 
            .Q(phase_accum[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i11.GSR = "ENABLED";
    FD1S3AX phase_accum_i12 (.D(phase_accum_63__N_146[12]), .CK(osc_clk), 
            .Q(phase_accum[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i12.GSR = "ENABLED";
    FD1S3AX phase_accum_i13 (.D(phase_accum_63__N_146[13]), .CK(osc_clk), 
            .Q(phase_accum[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i13.GSR = "ENABLED";
    FD1S3AX phase_accum_i14 (.D(phase_accum_63__N_146[14]), .CK(osc_clk), 
            .Q(phase_accum[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i14.GSR = "ENABLED";
    FD1S3AX phase_accum_i15 (.D(phase_accum_63__N_146[15]), .CK(osc_clk), 
            .Q(phase_accum[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i15.GSR = "ENABLED";
    FD1S3AX phase_accum_i16 (.D(phase_accum_63__N_146[16]), .CK(osc_clk), 
            .Q(phase_accum[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i16.GSR = "ENABLED";
    FD1S3AX phase_accum_i17 (.D(phase_accum_63__N_146[17]), .CK(osc_clk), 
            .Q(phase_accum[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i17.GSR = "ENABLED";
    FD1S3AX phase_accum_i18 (.D(phase_accum_63__N_146[18]), .CK(osc_clk), 
            .Q(phase_accum[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i18.GSR = "ENABLED";
    FD1S3AX phase_accum_i19 (.D(phase_accum_63__N_146[19]), .CK(osc_clk), 
            .Q(phase_accum[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i19.GSR = "ENABLED";
    FD1S3AX phase_accum_i20 (.D(phase_accum_63__N_146[20]), .CK(osc_clk), 
            .Q(phase_accum[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i20.GSR = "ENABLED";
    FD1S3AX phase_accum_i21 (.D(phase_accum_63__N_146[21]), .CK(osc_clk), 
            .Q(phase_accum[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i21.GSR = "ENABLED";
    FD1S3AX phase_accum_i22 (.D(phase_accum_63__N_146[22]), .CK(osc_clk), 
            .Q(phase_accum[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i22.GSR = "ENABLED";
    FD1S3AX phase_accum_i23 (.D(phase_accum_63__N_146[23]), .CK(osc_clk), 
            .Q(phase_accum[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i23.GSR = "ENABLED";
    FD1S3AX phase_accum_i24 (.D(phase_accum_63__N_146[24]), .CK(osc_clk), 
            .Q(phase_accum[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i24.GSR = "ENABLED";
    FD1S3AX phase_accum_i25 (.D(phase_accum_63__N_146[25]), .CK(osc_clk), 
            .Q(phase_accum[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i25.GSR = "ENABLED";
    FD1S3AX phase_accum_i26 (.D(phase_accum_63__N_146[26]), .CK(osc_clk), 
            .Q(phase_accum[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i26.GSR = "ENABLED";
    FD1S3AX phase_accum_i27 (.D(phase_accum_63__N_146[27]), .CK(osc_clk), 
            .Q(phase_accum[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i27.GSR = "ENABLED";
    FD1S3AX phase_accum_i28 (.D(phase_accum_63__N_146[28]), .CK(osc_clk), 
            .Q(phase_accum[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i28.GSR = "ENABLED";
    FD1S3AX phase_accum_i29 (.D(phase_accum_63__N_146[29]), .CK(osc_clk), 
            .Q(phase_accum[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i29.GSR = "ENABLED";
    FD1S3AX phase_accum_i30 (.D(phase_accum_63__N_146[30]), .CK(osc_clk), 
            .Q(phase_accum[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i30.GSR = "ENABLED";
    FD1S3AX phase_accum_i31 (.D(phase_accum_63__N_146[31]), .CK(osc_clk), 
            .Q(phase_accum[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i31.GSR = "ENABLED";
    FD1S3AX phase_accum_i32 (.D(phase_accum_63__N_146[32]), .CK(osc_clk), 
            .Q(phase_accum[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i32.GSR = "ENABLED";
    FD1S3AX phase_accum_i33 (.D(phase_accum_63__N_146[33]), .CK(osc_clk), 
            .Q(phase_accum[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i33.GSR = "ENABLED";
    FD1S3AX phase_accum_i34 (.D(phase_accum_63__N_146[34]), .CK(osc_clk), 
            .Q(phase_accum[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i34.GSR = "ENABLED";
    FD1S3AX phase_accum_i35 (.D(phase_accum_63__N_146[35]), .CK(osc_clk), 
            .Q(phase_accum[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i35.GSR = "ENABLED";
    FD1S3AX phase_accum_i36 (.D(phase_accum_63__N_146[36]), .CK(osc_clk), 
            .Q(phase_accum[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i36.GSR = "ENABLED";
    FD1S3AX phase_accum_i37 (.D(phase_accum_63__N_146[37]), .CK(osc_clk), 
            .Q(phase_accum[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i37.GSR = "ENABLED";
    FD1S3AX phase_accum_i38 (.D(phase_accum_63__N_146[38]), .CK(osc_clk), 
            .Q(phase_accum[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i38.GSR = "ENABLED";
    FD1S3AX phase_accum_i39 (.D(phase_accum_63__N_146[39]), .CK(osc_clk), 
            .Q(phase_accum[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i39.GSR = "ENABLED";
    FD1S3AX phase_accum_i40 (.D(phase_accum_63__N_146[40]), .CK(osc_clk), 
            .Q(phase_accum[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i40.GSR = "ENABLED";
    FD1S3AX phase_accum_i41 (.D(phase_accum_63__N_146[41]), .CK(osc_clk), 
            .Q(phase_accum[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i41.GSR = "ENABLED";
    FD1S3AX phase_accum_i42 (.D(phase_accum_63__N_146[42]), .CK(osc_clk), 
            .Q(phase_accum[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i42.GSR = "ENABLED";
    FD1S3AX phase_accum_i43 (.D(phase_accum_63__N_146[43]), .CK(osc_clk), 
            .Q(phase_accum[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i43.GSR = "ENABLED";
    FD1S3AX phase_accum_i44 (.D(phase_accum_63__N_146[44]), .CK(osc_clk), 
            .Q(phase_accum[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i44.GSR = "ENABLED";
    FD1S3AX phase_accum_i45 (.D(phase_accum_63__N_146[45]), .CK(osc_clk), 
            .Q(phase_accum[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i45.GSR = "ENABLED";
    FD1S3AX phase_accum_i46 (.D(phase_accum_63__N_146[46]), .CK(osc_clk), 
            .Q(phase_accum[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i46.GSR = "ENABLED";
    FD1S3AX phase_accum_i47 (.D(phase_accum_63__N_146[47]), .CK(osc_clk), 
            .Q(phase_accum[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i47.GSR = "ENABLED";
    FD1S3AX phase_accum_i48 (.D(phase_accum_63__N_146[48]), .CK(osc_clk), 
            .Q(phase_accum[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i48.GSR = "ENABLED";
    FD1S3AX phase_accum_i49 (.D(phase_accum_63__N_146[49]), .CK(osc_clk), 
            .Q(phase_accum[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i49.GSR = "ENABLED";
    FD1S3AX phase_accum_i50 (.D(phase_accum_63__N_146[50]), .CK(osc_clk), 
            .Q(phase_accum[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i50.GSR = "ENABLED";
    FD1S3AX phase_accum_i51 (.D(phase_accum_63__N_146[51]), .CK(osc_clk), 
            .Q(phase_accum[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i51.GSR = "ENABLED";
    FD1S3AX phase_accum_i52 (.D(phase_accum_63__N_146[52]), .CK(osc_clk), 
            .Q(phase_accum[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i52.GSR = "ENABLED";
    FD1S3AX phase_accum_i53 (.D(phase_accum_63__N_146[53]), .CK(osc_clk), 
            .Q(phase_accum[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i53.GSR = "ENABLED";
    FD1S3AX phase_accum_i54 (.D(phase_accum_63__N_146[54]), .CK(osc_clk), 
            .Q(phase_accum[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i54.GSR = "ENABLED";
    FD1S3AX phase_accum_i55 (.D(phase_accum_63__N_146[55]), .CK(osc_clk), 
            .Q(phase_accum[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i55.GSR = "ENABLED";
    FD1S3AX phase_accum_i56 (.D(phase_accum_63__N_146[56]), .CK(osc_clk), 
            .Q(\phase_accum[56] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i56.GSR = "ENABLED";
    FD1S3AX phase_accum_i57 (.D(phase_accum_63__N_146[57]), .CK(osc_clk), 
            .Q(\phase_accum[57] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i57.GSR = "ENABLED";
    FD1S3AX phase_accum_i58 (.D(phase_accum_63__N_146[58]), .CK(osc_clk), 
            .Q(\phase_accum[58] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i58.GSR = "ENABLED";
    FD1S3AX phase_accum_i59 (.D(phase_accum_63__N_146[59]), .CK(osc_clk), 
            .Q(\phase_accum[59] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i59.GSR = "ENABLED";
    FD1S3AX phase_accum_i60 (.D(phase_accum_63__N_146[60]), .CK(osc_clk), 
            .Q(\phase_accum[60] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i60.GSR = "ENABLED";
    FD1S3AX phase_accum_i61 (.D(phase_accum_63__N_146[61]), .CK(osc_clk), 
            .Q(\phase_accum[61] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i61.GSR = "ENABLED";
    FD1S3AX phase_accum_i62 (.D(phase_accum_63__N_146[62]), .CK(osc_clk), 
            .Q(\phase_accum[62] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i62.GSR = "ENABLED";
    FD1S3AX phase_accum_i63 (.D(phase_accum_63__N_146[63]), .CK(osc_clk), 
            .Q(\phase_accum[63] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=151, LSE_RLINE=157 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i63.GSR = "ENABLED";
    CCU2D phase_accum_63__I_0_12_64 (.A0(\phase_accum[62] ), .B0(phase_inc_carrGen1[62]), 
          .C0(GND_net), .D0(GND_net), .A1(\phase_accum[63] ), .B1(phase_inc_carrGen1[63]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10692), .S0(phase_accum_63__N_146[62]), 
          .S1(phase_accum_63__N_146[63]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_64.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_64.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_64.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_64.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_62 (.A0(\phase_accum[60] ), .B0(phase_inc_carrGen1[60]), 
          .C0(GND_net), .D0(GND_net), .A1(\phase_accum[61] ), .B1(phase_inc_carrGen1[61]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10691), .COUT(n10692), .S0(phase_accum_63__N_146[60]), 
          .S1(phase_accum_63__N_146[61]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_62.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_62.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_62.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_62.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_60 (.A0(\phase_accum[58] ), .B0(phase_inc_carrGen1[58]), 
          .C0(GND_net), .D0(GND_net), .A1(\phase_accum[59] ), .B1(phase_inc_carrGen1[59]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10690), .COUT(n10691), .S0(phase_accum_63__N_146[58]), 
          .S1(phase_accum_63__N_146[59]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_60.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_60.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_60.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_60.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_58 (.A0(\phase_accum[56] ), .B0(phase_inc_carrGen1[56]), 
          .C0(GND_net), .D0(GND_net), .A1(\phase_accum[57] ), .B1(phase_inc_carrGen1[57]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10689), .COUT(n10690), .S0(phase_accum_63__N_146[56]), 
          .S1(phase_accum_63__N_146[57]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_58.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_58.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_58.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_58.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_56 (.A0(phase_accum[54]), .B0(phase_inc_carrGen1[54]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[55]), .B1(phase_inc_carrGen1[55]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10688), .COUT(n10689), .S0(phase_accum_63__N_146[54]), 
          .S1(phase_accum_63__N_146[55]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_56.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_56.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_56.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_56.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_54 (.A0(phase_accum[52]), .B0(phase_inc_carrGen1[52]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[53]), .B1(phase_inc_carrGen1[53]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10687), .COUT(n10688), .S0(phase_accum_63__N_146[52]), 
          .S1(phase_accum_63__N_146[53]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_54.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_54.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_54.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_54.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_52 (.A0(phase_accum[50]), .B0(phase_inc_carrGen1[50]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[51]), .B1(phase_inc_carrGen1[51]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10686), .COUT(n10687), .S0(phase_accum_63__N_146[50]), 
          .S1(phase_accum_63__N_146[51]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_52.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_52.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_52.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_52.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_50 (.A0(phase_accum[48]), .B0(phase_inc_carrGen1[48]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[49]), .B1(phase_inc_carrGen1[49]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10685), .COUT(n10686), .S0(phase_accum_63__N_146[48]), 
          .S1(phase_accum_63__N_146[49]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_50.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_50.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_50.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_50.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_48 (.A0(phase_accum[46]), .B0(phase_inc_carrGen1[46]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[47]), .B1(phase_inc_carrGen1[47]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10684), .COUT(n10685), .S0(phase_accum_63__N_146[46]), 
          .S1(phase_accum_63__N_146[47]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_48.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_48.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_48.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_48.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_46 (.A0(phase_accum[44]), .B0(phase_inc_carrGen1[44]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[45]), .B1(phase_inc_carrGen1[45]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10683), .COUT(n10684), .S0(phase_accum_63__N_146[44]), 
          .S1(phase_accum_63__N_146[45]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_46.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_46.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_46.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_46.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_44 (.A0(phase_accum[42]), .B0(phase_inc_carrGen1[42]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[43]), .B1(phase_inc_carrGen1[43]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10682), .COUT(n10683), .S0(phase_accum_63__N_146[42]), 
          .S1(phase_accum_63__N_146[43]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_44.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_44.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_44.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_44.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_42 (.A0(phase_accum[40]), .B0(phase_inc_carrGen1[40]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[41]), .B1(phase_inc_carrGen1[41]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10681), .COUT(n10682), .S0(phase_accum_63__N_146[40]), 
          .S1(phase_accum_63__N_146[41]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_42.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_42.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_42.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_42.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_40 (.A0(phase_accum[38]), .B0(phase_inc_carrGen1[38]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[39]), .B1(phase_inc_carrGen1[39]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10680), .COUT(n10681), .S0(phase_accum_63__N_146[38]), 
          .S1(phase_accum_63__N_146[39]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_40.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_40.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_40.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_40.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_38 (.A0(phase_accum[36]), .B0(phase_inc_carrGen1[36]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[37]), .B1(phase_inc_carrGen1[37]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10679), .COUT(n10680), .S0(phase_accum_63__N_146[36]), 
          .S1(phase_accum_63__N_146[37]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_38.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_38.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_38.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_38.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_36 (.A0(phase_accum[34]), .B0(phase_inc_carrGen1[34]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[35]), .B1(phase_inc_carrGen1[35]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10678), .COUT(n10679), .S0(phase_accum_63__N_146[34]), 
          .S1(phase_accum_63__N_146[35]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_36.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_36.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_36.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_36.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_34 (.A0(phase_accum[32]), .B0(phase_inc_carrGen1[32]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[33]), .B1(phase_inc_carrGen1[33]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10677), .COUT(n10678), .S0(phase_accum_63__N_146[32]), 
          .S1(phase_accum_63__N_146[33]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_34.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_34.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_34.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_34.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_32 (.A0(phase_accum[30]), .B0(phase_inc_carrGen1[30]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[31]), .B1(phase_inc_carrGen1[31]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10676), .COUT(n10677), .S0(phase_accum_63__N_146[30]), 
          .S1(phase_accum_63__N_146[31]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_32.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_32.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_32.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_32.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_30 (.A0(phase_accum[28]), .B0(phase_inc_carrGen1[28]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[29]), .B1(phase_inc_carrGen1[29]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10675), .COUT(n10676), .S0(phase_accum_63__N_146[28]), 
          .S1(phase_accum_63__N_146[29]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_30.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_30.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_30.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_30.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_28 (.A0(phase_accum[26]), .B0(phase_inc_carrGen1[26]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[27]), .B1(phase_inc_carrGen1[27]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10674), .COUT(n10675), .S0(phase_accum_63__N_146[26]), 
          .S1(phase_accum_63__N_146[27]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_28.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_28.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_28.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_28.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_26 (.A0(phase_accum[24]), .B0(phase_inc_carrGen1[24]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[25]), .B1(phase_inc_carrGen1[25]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10673), .COUT(n10674), .S0(phase_accum_63__N_146[24]), 
          .S1(phase_accum_63__N_146[25]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_26.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_26.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_26.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_26.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_24 (.A0(phase_accum[22]), .B0(phase_inc_carrGen1[22]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[23]), .B1(phase_inc_carrGen1[23]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10672), .COUT(n10673), .S0(phase_accum_63__N_146[22]), 
          .S1(phase_accum_63__N_146[23]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_24.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_24.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_24.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_24.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_22 (.A0(phase_accum[20]), .B0(phase_inc_carrGen1[20]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[21]), .B1(phase_inc_carrGen1[21]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10671), .COUT(n10672), .S0(phase_accum_63__N_146[20]), 
          .S1(phase_accum_63__N_146[21]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_22.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_22.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_22.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_22.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_20 (.A0(phase_accum[18]), .B0(phase_inc_carrGen1[18]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[19]), .B1(phase_inc_carrGen1[19]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10670), .COUT(n10671), .S0(phase_accum_63__N_146[18]), 
          .S1(phase_accum_63__N_146[19]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_20.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_20.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_20.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_20.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_18 (.A0(phase_accum[16]), .B0(phase_inc_carrGen1[16]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[17]), .B1(phase_inc_carrGen1[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10669), .COUT(n10670), .S0(phase_accum_63__N_146[16]), 
          .S1(phase_accum_63__N_146[17]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_18.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_18.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_18.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_18.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_16 (.A0(phase_accum[14]), .B0(phase_inc_carrGen1[14]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[15]), .B1(phase_inc_carrGen1[15]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10668), .COUT(n10669), .S0(phase_accum_63__N_146[14]), 
          .S1(phase_accum_63__N_146[15]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_16.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_16.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_16.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_16.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_14 (.A0(phase_accum[12]), .B0(phase_inc_carrGen1[12]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[13]), .B1(phase_inc_carrGen1[13]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10667), .COUT(n10668), .S0(phase_accum_63__N_146[12]), 
          .S1(phase_accum_63__N_146[13]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_14.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_14.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_14.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_14.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_12 (.A0(phase_accum[10]), .B0(phase_inc_carrGen1[10]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[11]), .B1(phase_inc_carrGen1[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10666), .COUT(n10667), .S0(phase_accum_63__N_146[10]), 
          .S1(phase_accum_63__N_146[11]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_12.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_12.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_12.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_12.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_10 (.A0(phase_accum[8]), .B0(phase_inc_carrGen1[8]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[9]), .B1(phase_inc_carrGen1[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10665), .COUT(n10666), .S0(phase_accum_63__N_146[8]), 
          .S1(phase_accum_63__N_146[9]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_10.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_10.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_10.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_10.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_8 (.A0(phase_accum[6]), .B0(phase_inc_carrGen1[6]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[7]), .B1(phase_inc_carrGen1[7]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10664), .COUT(n10665), .S0(phase_accum_63__N_146[6]), 
          .S1(phase_accum_63__N_146[7]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_8.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_8.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_8.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_8.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_6 (.A0(phase_accum[4]), .B0(phase_inc_carrGen1[4]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[5]), .B1(phase_inc_carrGen1[5]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10663), .COUT(n10664), .S0(phase_accum_63__N_146[4]), 
          .S1(phase_accum_63__N_146[5]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_6.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_6.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_6.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_6.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_4 (.A0(phase_accum[2]), .B0(phase_inc_carrGen1[2]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[3]), .B1(phase_inc_carrGen1[3]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10662), .COUT(n10663), .S0(phase_accum_63__N_146[2]), 
          .S1(phase_accum_63__N_146[3]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_4.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_4.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_4.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_4.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_2 (.A0(phase_accum[0]), .B0(phase_inc_carrGen1[0]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[1]), .B1(phase_inc_carrGen1[1]), 
          .C1(GND_net), .D1(GND_net), .COUT(n10662), .S1(phase_accum_63__N_146[1]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_2.INIT0 = 16'h7000;
    defparam phase_accum_63__I_0_12_2.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_2.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_2.INJECT1_1 = "NO";
    LUT4 phase_accum_63__I_0_13_1_lut (.A(\phase_accum[63] ), .Z(sinGen_c)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(32[18:56])
    defparam phase_accum_63__I_0_13_1_lut.init = 16'h5555;
    LUT4 i4594_2_lut (.A(phase_accum[0]), .B(phase_inc_carrGen1[0]), .Z(phase_accum_63__N_146[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4594_2_lut.init = 16'h6666;
    
endmodule
//
// Verilog Description of module \CIC(width=72,decimation_ratio=4096)_U1 
//

module \CIC(width=72,decimation_ratio=4096)_U1  (GND_net, MixerOutCos, osc_clk, 
            CIC1_outCos, \d10[61] , \d10[62] , \CICGain[0] , n62, 
            \d10[63] , n63, \d10[64] , n64, \d10[65] , n65, \d10[66] , 
            n66, \d10[60] , n61, \d10[67] , n67, \d10[68] , n68, 
            \d10[69] , \d10[70] , n70, \d10[59] , \d10[71] , \d_out_11__N_1819[2] , 
            \d_out_11__N_1819[3] , \d_out_11__N_1819[4] , \d_out_11__N_1819[5] , 
            \d_out_11__N_1819[6] , \d_out_11__N_1819[7] , \d_out_11__N_1819[8] , 
            \d_out_11__N_1819[9] , \d_out_11__N_1819[10] , \d_out_11__N_1819[11] , 
            \CICGain[1] ) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input [11:0]MixerOutCos;
    input osc_clk;
    output [11:0]CIC1_outCos;
    output \d10[61] ;
    output \d10[62] ;
    input \CICGain[0] ;
    output n62;
    output \d10[63] ;
    output n63;
    output \d10[64] ;
    output n64;
    output \d10[65] ;
    output n65;
    output \d10[66] ;
    output n66;
    output \d10[60] ;
    output n61;
    output \d10[67] ;
    output n67;
    output \d10[68] ;
    output n68;
    output \d10[69] ;
    output \d10[70] ;
    output n70;
    output \d10[59] ;
    output \d10[71] ;
    input \d_out_11__N_1819[2] ;
    input \d_out_11__N_1819[3] ;
    input \d_out_11__N_1819[4] ;
    input \d_out_11__N_1819[5] ;
    input \d_out_11__N_1819[6] ;
    input \d_out_11__N_1819[7] ;
    input \d_out_11__N_1819[8] ;
    input \d_out_11__N_1819[9] ;
    input \d_out_11__N_1819[10] ;
    input \d_out_11__N_1819[11] ;
    input \CICGain[1] ;
    
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(69[8:15])
    
    wire n11737;
    wire [71:0]d1;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(35[26:28])
    wire [71:0]d2;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(36[26:28])
    wire [35:0]n5212;
    
    wire n11738, n11736, n11735, n11599;
    wire [71:0]d5;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(39[26:28])
    
    wire n5667;
    wire [35:0]n5668;
    wire [71:0]d4;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(38[26:28])
    wire [71:0]d5_71__N_706;
    
    wire n11600;
    wire [35:0]n6732;
    wire [35:0]n6770;
    
    wire n6731;
    wire [71:0]d10_71__N_1747;
    
    wire n11756, n5059;
    wire [35:0]n5060;
    wire [71:0]d1_71__N_418;
    
    wire n11757, n11755, n11750;
    wire [71:0]d_tmp;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(30[26:31])
    
    wire osc_clk_enable_757;
    wire [71:0]d_d_tmp;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(30[33:40])
    
    wire osc_clk_enable_797;
    wire [71:0]d2_71__N_490;
    wire [71:0]d3;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(37[26:28])
    wire [71:0]d3_71__N_562;
    wire [71:0]d4_71__N_634;
    wire [71:0]d6;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(43[26:28])
    wire [71:0]d6_71__N_1459;
    
    wire v_comb;
    wire [71:0]d_d6;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(43[30:34])
    wire [71:0]d7;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(44[26:28])
    wire [71:0]d7_71__N_1531;
    wire [71:0]d_d7;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(44[30:34])
    wire [71:0]d8;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(45[26:28])
    wire [71:0]d8_71__N_1603;
    wire [71:0]d_d8;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(45[30:34])
    wire [71:0]d9;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(46[26:28])
    wire [71:0]d9_71__N_1675;
    wire [71:0]d_d9;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(46[30:34])
    wire [71:0]d_out_11__N_1819;
    
    wire n11598, n11744, n11745, n11602, n11603, n11743, n11742, 
        n11741, n11740, n11674, n5363;
    wire [35:0]n5364;
    
    wire n11675, n11739, n11734, n11673, n11730, n5211, n11731, 
        n11597, n11717, n11718, n11716, n11714, n11708, n11709, 
        n11715, n11707, n11668;
    wire [35:0]n5516;
    
    wire n11667, n11330;
    wire [35:0]n6124;
    wire [15:0]count;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(50[14:19])
    wire [15:0]count_15__N_1442;
    
    wire n11666, n11665, n11664, n11608, n11663, n11607, n11706, 
        n11702, n11703, n11596, n11693, n11689, n11690, n11688, 
        n11606, n12778, n12503, n12780, n13196, n11687, n11683, 
        n11684, n11677, n11678, n11662, n11676, n11682, n11681, 
        n11686, n11680, n11679, n11685, n11595, n11719, n11720;
    wire [15:0]n375;
    
    wire n31, n22, n18, n11594, n11593, n11592, n19, n15, n11591, 
        n11729, n11604, n11605, n11728, n11727, n11726, n11725, 
        n11724, n11601, n11329, n11328, n11327, n11326, n11325, 
        n11324, n11323, n11322, n11321, n11696, n11697, n11320, 
        n11319, n11318, n11661, n11660, n11695, n11659, n11701, 
        n11694, n11700, n11705, n11699, n11698, n7, n11704, n11749, 
        n11748, n11723, n11658, n11721, n11722, n11747, n11746, 
        n11657, n11656, n11655, n11654, n11653, n11652, n11317, 
        n11649, n5515, n11648, n11647, n11646, n11645, n11644, 
        n11643, n11642, n11641, n11640, n11639, n11638, n11637, 
        n11636, n11635, n11634, n11633, n11632, n11627, n11626, 
        n11625, n11624, n11623, n11622, n11621, n11620, n11619, 
        n11618, n11617, n11616, n11615, n11614, n11613, n11612, 
        n11611, count_15__N_1458, osc_clk_enable_847, osc_clk_enable_897, 
        osc_clk_enable_947, osc_clk_enable_997, osc_clk_enable_1047, osc_clk_enable_1097, 
        osc_clk_enable_1147, osc_clk_enable_1197, osc_clk_enable_1247, 
        osc_clk_enable_1297, osc_clk_enable_1347, osc_clk_enable_1397;
    wire [71:0]d10;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(47[26:29])
    
    wire n11316, n11315, n11314, n11313, n11311, n6123, n11310, 
        n11309, n11308, n11307, n11306, n11305, n11304, n11303, 
        n11302, n11301, n11300, n11299, n11298, n11297, n11296, 
        n11295, n11294, n11290;
    wire [35:0]n6276;
    
    wire n11289, n11288, n11287, n11286, n11285, n11284, n11283, 
        n11282, n11281, n11280, n11279, n11278, n11277, n11276, 
        n11275, n11274, n11273, n11271, n6275, n11270, n11269, 
        n11268, n11267, n11266, n11265, n11264, n11263, n11262, 
        n11261, n11260, n11259, n11258, n11257, n11256, n11255, 
        n11254, n11250;
    wire [35:0]n6428;
    
    wire n11249, n11248, n11247, n11246, n11245, n11244, n11243, 
        n11242, n11241, n11240, n11239, n11238, n11237, n11236, 
        n11235, n11234, n11233, n11231, n6427, n11230, n11229, 
        n11228, n11227, n11226, n11225, n11224, n11223, n11222, 
        n11221, n11220, n11219, n11218, n11217, n11216, n11215, 
        n11214, n11210;
    wire [35:0]n6580;
    
    wire n11209, n11208, n11207, n11206, n11205, n11204, n11203, 
        n11202, n11201, n11200, n11199, n11198, n11197, n11196, 
        n11195, n11194, n11193, n11191, n6579, n11190, n11189, 
        n11188, n11187, n11186, n11185, n11184, n11183, n11182, 
        n11181, n11180, n11179, n11178, n11177, n11176, n11175, 
        n11174, n11170, n11169, n11168, n11167, n11166, n11165, 
        n11164, n11163, n11162, n11161, n11160, n11159, n11158, 
        n11157, n11156, n11155, n11154, n11153, n11152, n11151, 
        n11150, n11149, n11148, n11147, n11146, n11145, n11144, 
        n11143, n11142, n11141, n11140, n11139, n11138, n11137, 
        n11136, n11135, n8436, n10938, n10937, n10936, n10935, 
        n10934, n10933, n10932, n10931, n10912, n10911, n10910, 
        n10909, n10908, n10907, n10906, n10905, n10904, n10903, 
        n10902, n10901, n10900, n10899, n10898, n10897, n10896, 
        n10895, n10893, n10892, n10891, n10890, n10889, n10888, 
        n10887, n10886, n10885, n10884, n10883, n10882, n10881, 
        n10880, n10879, n10878, n10877, n10876, n10874, n10873, 
        n10872, n10871, n10870, n10869, n10868, n10867, n10866, 
        n10865, n10864, n10863, n10862, n10861, n10860, n10859, 
        n10858, n10857, n10855, n10854, n10853, n10852, n10851, 
        n10850, n10849, n10848, n10847, n10846, n10845, n10844, 
        n10843, n10842, n10841, n10840, n10839, n10838, n10798, 
        n10797, n10796, n10795, n10794, n10793, n10792, n10791, 
        n10790, n10789, n10788, n10787, n10786, n10785, n10784, 
        n10783, n10782, n10781, n11452, n11451, n11450, n11449, 
        n11448, n11447, n11446, n11445, n11444, n11443, n11442, 
        n11441, n11440, n11439, n11438, n11437, n11436, n11435, 
        n11434, n11433, n11432, n11431, n11430, n11429, n11428, 
        n11427, n11426, n11425, n11424, n11423, n11422, n11421, 
        n11420, n11419, n11418, n11417, n11416, n11415, n11414, 
        n11413, n11412, n11411, n11410, n11409, n11408, n11407, 
        n11406, n11405, n11404, n11403, n11402, n11401, n11400, 
        n11399, n11398, n11397, n11396, n11395, n11394, n11393, 
        n11392, n11391, n11390, n11389, n11388, n11387, n11386, 
        n11385, n11384, n11383, n11382, n11381, n11380, n11379, 
        n11378, n11377, n11376, n11375, n11374, n11373, n11372, 
        n11371, n11370, n11369, n11368, n11367, n11366, n11365, 
        n11364, n11363, n12, n8, n11758, n11761, n11762, n11772, 
        n11771, n11770, n11769, n11768, n11767, n11766, n13089, 
        n13090, n13087, n13086, n11765, n11764, n11760, n11759, 
        n11763, n11791, n11790, n11789, n11788, n11787, n11786, 
        n11785, n11784, n11783, n11782, n11781, n11780, n11779, 
        n11778, n11777, n11776, n11775;
    
    CCU2D add_1081_10 (.A0(d1[44]), .B0(d2[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[45]), .B1(d2[45]), .C1(GND_net), .D1(GND_net), .CIN(n11737), 
          .COUT(n11738), .S0(n5212[8]), .S1(n5212[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1081_10.INIT0 = 16'h5666;
    defparam add_1081_10.INIT1 = 16'h5666;
    defparam add_1081_10.INJECT1_0 = "NO";
    defparam add_1081_10.INJECT1_1 = "NO";
    CCU2D add_1081_8 (.A0(d1[42]), .B0(d2[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[43]), .B1(d2[43]), .C1(GND_net), .D1(GND_net), .CIN(n11736), 
          .COUT(n11737), .S0(n5212[6]), .S1(n5212[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1081_8.INIT0 = 16'h5666;
    defparam add_1081_8.INIT1 = 16'h5666;
    defparam add_1081_8.INJECT1_0 = "NO";
    defparam add_1081_8.INJECT1_1 = "NO";
    CCU2D add_1081_6 (.A0(d1[40]), .B0(d2[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[41]), .B1(d2[41]), .C1(GND_net), .D1(GND_net), .CIN(n11735), 
          .COUT(n11736), .S0(n5212[4]), .S1(n5212[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1081_6.INIT0 = 16'h5666;
    defparam add_1081_6.INIT1 = 16'h5666;
    defparam add_1081_6.INJECT1_0 = "NO";
    defparam add_1081_6.INJECT1_1 = "NO";
    CCU2D add_1097_19 (.A0(d5[52]), .B0(n5667), .C0(n5668[16]), .D0(d4[52]), 
          .A1(d5[53]), .B1(n5667), .C1(n5668[17]), .D1(d4[53]), .CIN(n11599), 
          .COUT(n11600), .S0(d5_71__N_706[52]), .S1(d5_71__N_706[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1097_19.INIT0 = 16'h74b8;
    defparam add_1097_19.INIT1 = 16'h74b8;
    defparam add_1097_19.INJECT1_0 = "NO";
    defparam add_1097_19.INJECT1_1 = "NO";
    LUT4 mux_1243_i15_3_lut (.A(n6732[34]), .B(n6770[34]), .C(n6731), 
         .Z(d10_71__N_1747[70])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1243_i15_3_lut.init = 16'hcaca;
    CCU2D add_1077_5 (.A0(d1[38]), .B0(n5059), .C0(n5060[2]), .D0(MixerOutCos[11]), 
          .A1(d1[39]), .B1(n5059), .C1(n5060[3]), .D1(MixerOutCos[11]), 
          .CIN(n11756), .COUT(n11757), .S0(d1_71__N_418[38]), .S1(d1_71__N_418[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1077_5.INIT0 = 16'h74b8;
    defparam add_1077_5.INIT1 = 16'h74b8;
    defparam add_1077_5.INJECT1_0 = "NO";
    defparam add_1077_5.INJECT1_1 = "NO";
    CCU2D add_1077_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5059), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11755));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1077_1.INIT0 = 16'hF000;
    defparam add_1077_1.INIT1 = 16'h0555;
    defparam add_1077_1.INJECT1_0 = "NO";
    defparam add_1077_1.INJECT1_1 = "NO";
    CCU2D add_1077_3 (.A0(d1[36]), .B0(n5059), .C0(n5060[0]), .D0(MixerOutCos[11]), 
          .A1(d1[37]), .B1(n5059), .C1(n5060[1]), .D1(MixerOutCos[11]), 
          .CIN(n11755), .COUT(n11756), .S0(d1_71__N_418[36]), .S1(d1_71__N_418[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1077_3.INIT0 = 16'h74b8;
    defparam add_1077_3.INIT1 = 16'h74b8;
    defparam add_1077_3.INJECT1_0 = "NO";
    defparam add_1077_3.INJECT1_1 = "NO";
    CCU2D add_1081_36 (.A0(d1[70]), .B0(d2[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[71]), .B1(d2[71]), .C1(GND_net), .D1(GND_net), .CIN(n11750), 
          .S0(n5212[34]), .S1(n5212[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1081_36.INIT0 = 16'h5666;
    defparam add_1081_36.INIT1 = 16'h5666;
    defparam add_1081_36.INJECT1_0 = "NO";
    defparam add_1081_36.INJECT1_1 = "NO";
    LUT4 i4605_2_lut (.A(d4[0]), .B(d5[0]), .Z(d5_71__N_706[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4605_2_lut.init = 16'h6666;
    FD1P3AX d_tmp_i0_i0 (.D(d5[0]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i0 (.D(d_tmp[0]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i0.GSR = "ENABLED";
    LUT4 mux_1243_i16_3_lut (.A(n6732[35]), .B(n6770[35]), .C(n6731), 
         .Z(d10_71__N_1747[71])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1243_i16_3_lut.init = 16'hcaca;
    FD1S3AX d2_i0 (.D(d2_71__N_490[0]), .CK(osc_clk), .Q(d2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i0.GSR = "ENABLED";
    FD1S3AX d3_i0 (.D(d3_71__N_562[0]), .CK(osc_clk), .Q(d3[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i0.GSR = "ENABLED";
    FD1S3AX d4_i0 (.D(d4_71__N_634[0]), .CK(osc_clk), .Q(d4[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i0.GSR = "ENABLED";
    FD1S3AX d5_i0 (.D(d5_71__N_706[0]), .CK(osc_clk), .Q(d5[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i0.GSR = "ENABLED";
    FD1P3AX d6_i0_i0 (.D(d6_71__N_1459[0]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i0.GSR = "ENABLED";
    FD1S3AX v_comb_66 (.D(osc_clk_enable_757), .CK(osc_clk), .Q(v_comb)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i0 (.D(d6[0]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i0.GSR = "ENABLED";
    FD1P3AX d7_i0_i0 (.D(d7_71__N_1531[0]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i0.GSR = "ENABLED";
    LUT4 i4643_2_lut (.A(MixerOutCos[11]), .B(d1[36]), .Z(n5060[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4643_2_lut.init = 16'h6666;
    FD1P3AX d_d7_i0_i0 (.D(d7[0]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d8_i0_i0 (.D(d8_71__N_1603[0]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i0 (.D(d8[0]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d9_i0_i0 (.D(d9_71__N_1675[0]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i0 (.D(d9[0]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_out_i0_i0 (.D(d_out_11__N_1819[0]), .SP(osc_clk_enable_797), 
            .CK(osc_clk), .Q(CIC1_outCos[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i0.GSR = "ENABLED";
    FD1S3AX d1_i0 (.D(d1_71__N_418[0]), .CK(osc_clk), .Q(d1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i0.GSR = "ENABLED";
    CCU2D add_1097_17 (.A0(d5[50]), .B0(n5667), .C0(n5668[14]), .D0(d4[50]), 
          .A1(d5[51]), .B1(n5667), .C1(n5668[15]), .D1(d4[51]), .CIN(n11598), 
          .COUT(n11599), .S0(d5_71__N_706[50]), .S1(d5_71__N_706[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1097_17.INIT0 = 16'h74b8;
    defparam add_1097_17.INIT1 = 16'h74b8;
    defparam add_1097_17.INJECT1_0 = "NO";
    defparam add_1097_17.INJECT1_1 = "NO";
    CCU2D add_1081_24 (.A0(d1[58]), .B0(d2[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[59]), .B1(d2[59]), .C1(GND_net), .D1(GND_net), .CIN(n11744), 
          .COUT(n11745), .S0(n5212[22]), .S1(n5212[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1081_24.INIT0 = 16'h5666;
    defparam add_1081_24.INIT1 = 16'h5666;
    defparam add_1081_24.INJECT1_0 = "NO";
    defparam add_1081_24.INJECT1_1 = "NO";
    CCU2D add_1097_25 (.A0(d5[58]), .B0(n5667), .C0(n5668[22]), .D0(d4[58]), 
          .A1(d5[59]), .B1(n5667), .C1(n5668[23]), .D1(d4[59]), .CIN(n11602), 
          .COUT(n11603), .S0(d5_71__N_706[58]), .S1(d5_71__N_706[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1097_25.INIT0 = 16'h74b8;
    defparam add_1097_25.INIT1 = 16'h74b8;
    defparam add_1097_25.INJECT1_0 = "NO";
    defparam add_1097_25.INJECT1_1 = "NO";
    CCU2D add_1081_22 (.A0(d1[56]), .B0(d2[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[57]), .B1(d2[57]), .C1(GND_net), .D1(GND_net), .CIN(n11743), 
          .COUT(n11744), .S0(n5212[20]), .S1(n5212[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1081_22.INIT0 = 16'h5666;
    defparam add_1081_22.INIT1 = 16'h5666;
    defparam add_1081_22.INJECT1_0 = "NO";
    defparam add_1081_22.INJECT1_1 = "NO";
    CCU2D add_1081_20 (.A0(d1[54]), .B0(d2[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[55]), .B1(d2[55]), .C1(GND_net), .D1(GND_net), .CIN(n11742), 
          .COUT(n11743), .S0(n5212[18]), .S1(n5212[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1081_20.INIT0 = 16'h5666;
    defparam add_1081_20.INIT1 = 16'h5666;
    defparam add_1081_20.INJECT1_0 = "NO";
    defparam add_1081_20.INJECT1_1 = "NO";
    CCU2D add_1081_18 (.A0(d1[52]), .B0(d2[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[53]), .B1(d2[53]), .C1(GND_net), .D1(GND_net), .CIN(n11741), 
          .COUT(n11742), .S0(n5212[16]), .S1(n5212[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1081_18.INIT0 = 16'h5666;
    defparam add_1081_18.INIT1 = 16'h5666;
    defparam add_1081_18.INJECT1_0 = "NO";
    defparam add_1081_18.INJECT1_1 = "NO";
    CCU2D add_1081_16 (.A0(d1[50]), .B0(d2[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[51]), .B1(d2[51]), .C1(GND_net), .D1(GND_net), .CIN(n11740), 
          .COUT(n11741), .S0(n5212[14]), .S1(n5212[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1081_16.INIT0 = 16'h5666;
    defparam add_1081_16.INIT1 = 16'h5666;
    defparam add_1081_16.INJECT1_0 = "NO";
    defparam add_1081_16.INJECT1_1 = "NO";
    CCU2D add_1087_5 (.A0(d3[38]), .B0(n5363), .C0(n5364[2]), .D0(d2[38]), 
          .A1(d3[39]), .B1(n5363), .C1(n5364[3]), .D1(d2[39]), .CIN(n11674), 
          .COUT(n11675), .S0(d3_71__N_562[38]), .S1(d3_71__N_562[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1087_5.INIT0 = 16'h74b8;
    defparam add_1087_5.INIT1 = 16'h74b8;
    defparam add_1087_5.INJECT1_0 = "NO";
    defparam add_1087_5.INJECT1_1 = "NO";
    CCU2D add_1081_14 (.A0(d1[48]), .B0(d2[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[49]), .B1(d2[49]), .C1(GND_net), .D1(GND_net), .CIN(n11739), 
          .COUT(n11740), .S0(n5212[12]), .S1(n5212[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1081_14.INIT0 = 16'h5666;
    defparam add_1081_14.INIT1 = 16'h5666;
    defparam add_1081_14.INJECT1_0 = "NO";
    defparam add_1081_14.INJECT1_1 = "NO";
    CCU2D add_1081_4 (.A0(d1[38]), .B0(d2[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[39]), .B1(d2[39]), .C1(GND_net), .D1(GND_net), .CIN(n11734), 
          .COUT(n11735), .S0(n5212[2]), .S1(n5212[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1081_4.INIT0 = 16'h5666;
    defparam add_1081_4.INIT1 = 16'h5666;
    defparam add_1081_4.INJECT1_0 = "NO";
    defparam add_1081_4.INJECT1_1 = "NO";
    CCU2D add_1087_3 (.A0(d3[36]), .B0(n5363), .C0(n5364[0]), .D0(d2[36]), 
          .A1(d3[37]), .B1(n5363), .C1(n5364[1]), .D1(d2[37]), .CIN(n11673), 
          .COUT(n11674), .S0(d3_71__N_562[36]), .S1(d3_71__N_562[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1087_3.INIT0 = 16'h74b8;
    defparam add_1087_3.INIT1 = 16'h74b8;
    defparam add_1087_3.INJECT1_0 = "NO";
    defparam add_1087_3.INJECT1_1 = "NO";
    CCU2D add_1087_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5363), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11673));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1087_1.INIT0 = 16'hF000;
    defparam add_1087_1.INIT1 = 16'h0555;
    defparam add_1087_1.INJECT1_0 = "NO";
    defparam add_1087_1.INJECT1_1 = "NO";
    CCU2D add_1081_12 (.A0(d1[46]), .B0(d2[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[47]), .B1(d2[47]), .C1(GND_net), .D1(GND_net), .CIN(n11738), 
          .COUT(n11739), .S0(n5212[10]), .S1(n5212[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1081_12.INIT0 = 16'h5666;
    defparam add_1081_12.INIT1 = 16'h5666;
    defparam add_1081_12.INJECT1_0 = "NO";
    defparam add_1081_12.INJECT1_1 = "NO";
    CCU2D add_1082_35 (.A0(d2[68]), .B0(n5211), .C0(n5212[32]), .D0(d1[68]), 
          .A1(d2[69]), .B1(n5211), .C1(n5212[33]), .D1(d1[69]), .CIN(n11730), 
          .COUT(n11731), .S0(d2_71__N_490[68]), .S1(d2_71__N_490[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1082_35.INIT0 = 16'h74b8;
    defparam add_1082_35.INIT1 = 16'h74b8;
    defparam add_1082_35.INJECT1_0 = "NO";
    defparam add_1082_35.INJECT1_1 = "NO";
    CCU2D add_1097_15 (.A0(d5[48]), .B0(n5667), .C0(n5668[12]), .D0(d4[48]), 
          .A1(d5[49]), .B1(n5667), .C1(n5668[13]), .D1(d4[49]), .CIN(n11597), 
          .COUT(n11598), .S0(d5_71__N_706[48]), .S1(d5_71__N_706[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1097_15.INIT0 = 16'h74b8;
    defparam add_1097_15.INIT1 = 16'h74b8;
    defparam add_1097_15.INJECT1_0 = "NO";
    defparam add_1097_15.INJECT1_1 = "NO";
    CCU2D add_1082_9 (.A0(d2[42]), .B0(n5211), .C0(n5212[6]), .D0(d1[42]), 
          .A1(d2[43]), .B1(n5211), .C1(n5212[7]), .D1(d1[43]), .CIN(n11717), 
          .COUT(n11718), .S0(d2_71__N_490[42]), .S1(d2_71__N_490[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1082_9.INIT0 = 16'h74b8;
    defparam add_1082_9.INIT1 = 16'h74b8;
    defparam add_1082_9.INJECT1_0 = "NO";
    defparam add_1082_9.INJECT1_1 = "NO";
    CCU2D add_1082_7 (.A0(d2[40]), .B0(n5211), .C0(n5212[4]), .D0(d1[40]), 
          .A1(d2[41]), .B1(n5211), .C1(n5212[5]), .D1(d1[41]), .CIN(n11716), 
          .COUT(n11717), .S0(d2_71__N_490[40]), .S1(d2_71__N_490[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1082_7.INIT0 = 16'h74b8;
    defparam add_1082_7.INIT1 = 16'h74b8;
    defparam add_1082_7.INJECT1_0 = "NO";
    defparam add_1082_7.INJECT1_1 = "NO";
    CCU2D add_1082_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5211), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11714));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1082_1.INIT0 = 16'hF000;
    defparam add_1082_1.INIT1 = 16'h0555;
    defparam add_1082_1.INJECT1_0 = "NO";
    defparam add_1082_1.INJECT1_1 = "NO";
    CCU2D add_1086_34 (.A0(d2[68]), .B0(d3[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[69]), .B1(d3[69]), .C1(GND_net), .D1(GND_net), .CIN(n11708), 
          .COUT(n11709), .S0(n5364[32]), .S1(n5364[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1086_34.INIT0 = 16'h5666;
    defparam add_1086_34.INIT1 = 16'h5666;
    defparam add_1086_34.INJECT1_0 = "NO";
    defparam add_1086_34.INJECT1_1 = "NO";
    CCU2D add_1082_5 (.A0(d2[38]), .B0(n5211), .C0(n5212[2]), .D0(d1[38]), 
          .A1(d2[39]), .B1(n5211), .C1(n5212[3]), .D1(d1[39]), .CIN(n11715), 
          .COUT(n11716), .S0(d2_71__N_490[38]), .S1(d2_71__N_490[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1082_5.INIT0 = 16'h74b8;
    defparam add_1082_5.INIT1 = 16'h74b8;
    defparam add_1082_5.INJECT1_0 = "NO";
    defparam add_1082_5.INJECT1_1 = "NO";
    CCU2D add_1086_36 (.A0(d2[70]), .B0(d3[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[71]), .B1(d3[71]), .C1(GND_net), .D1(GND_net), .CIN(n11709), 
          .S0(n5364[34]), .S1(n5364[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1086_36.INIT0 = 16'h5666;
    defparam add_1086_36.INIT1 = 16'h5666;
    defparam add_1086_36.INJECT1_0 = "NO";
    defparam add_1086_36.INJECT1_1 = "NO";
    CCU2D add_1086_32 (.A0(d2[66]), .B0(d3[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[67]), .B1(d3[67]), .C1(GND_net), .D1(GND_net), .CIN(n11707), 
          .COUT(n11708), .S0(n5364[30]), .S1(n5364[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1086_32.INIT0 = 16'h5666;
    defparam add_1086_32.INIT1 = 16'h5666;
    defparam add_1086_32.INJECT1_0 = "NO";
    defparam add_1086_32.INJECT1_1 = "NO";
    CCU2D add_1082_3 (.A0(d2[36]), .B0(n5211), .C0(n5212[0]), .D0(d1[36]), 
          .A1(d2[37]), .B1(n5211), .C1(n5212[1]), .D1(d1[37]), .CIN(n11714), 
          .COUT(n11715), .S0(d2_71__N_490[36]), .S1(d2_71__N_490[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1082_3.INIT0 = 16'h74b8;
    defparam add_1082_3.INIT1 = 16'h74b8;
    defparam add_1082_3.INJECT1_0 = "NO";
    defparam add_1082_3.INJECT1_1 = "NO";
    CCU2D add_1091_36 (.A0(d3[70]), .B0(d4[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[71]), .B1(d4[71]), .C1(GND_net), .D1(GND_net), .CIN(n11668), 
          .S0(n5516[34]), .S1(n5516[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1091_36.INIT0 = 16'h5666;
    defparam add_1091_36.INIT1 = 16'h5666;
    defparam add_1091_36.INJECT1_0 = "NO";
    defparam add_1091_36.INJECT1_1 = "NO";
    CCU2D add_1091_34 (.A0(d3[68]), .B0(d4[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[69]), .B1(d4[69]), .C1(GND_net), .D1(GND_net), .CIN(n11667), 
          .COUT(n11668), .S0(n5516[32]), .S1(n5516[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1091_34.INIT0 = 16'h5666;
    defparam add_1091_34.INIT1 = 16'h5666;
    defparam add_1091_34.INJECT1_0 = "NO";
    defparam add_1091_34.INJECT1_1 = "NO";
    CCU2D add_1111_37 (.A0(d_tmp[71]), .B0(d_d_tmp[71]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11330), .S0(n6124[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1111_37.INIT0 = 16'h5999;
    defparam add_1111_37.INIT1 = 16'h0000;
    defparam add_1111_37.INJECT1_0 = "NO";
    defparam add_1111_37.INJECT1_1 = "NO";
    FD1S3IX count__i0 (.D(count_15__N_1442[0]), .CK(osc_clk), .CD(osc_clk_enable_757), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i0.GSR = "ENABLED";
    CCU2D add_1091_32 (.A0(d3[66]), .B0(d4[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[67]), .B1(d4[67]), .C1(GND_net), .D1(GND_net), .CIN(n11666), 
          .COUT(n11667), .S0(n5516[30]), .S1(n5516[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1091_32.INIT0 = 16'h5666;
    defparam add_1091_32.INIT1 = 16'h5666;
    defparam add_1091_32.INJECT1_0 = "NO";
    defparam add_1091_32.INJECT1_1 = "NO";
    CCU2D add_1091_30 (.A0(d3[64]), .B0(d4[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[65]), .B1(d4[65]), .C1(GND_net), .D1(GND_net), .CIN(n11665), 
          .COUT(n11666), .S0(n5516[28]), .S1(n5516[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1091_30.INIT0 = 16'h5666;
    defparam add_1091_30.INIT1 = 16'h5666;
    defparam add_1091_30.INJECT1_0 = "NO";
    defparam add_1091_30.INJECT1_1 = "NO";
    CCU2D add_1091_28 (.A0(d3[62]), .B0(d4[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[63]), .B1(d4[63]), .C1(GND_net), .D1(GND_net), .CIN(n11664), 
          .COUT(n11665), .S0(n5516[26]), .S1(n5516[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1091_28.INIT0 = 16'h5666;
    defparam add_1091_28.INIT1 = 16'h5666;
    defparam add_1091_28.INJECT1_0 = "NO";
    defparam add_1091_28.INJECT1_1 = "NO";
    CCU2D add_1097_37 (.A0(d5[70]), .B0(n5667), .C0(n5668[34]), .D0(d4[70]), 
          .A1(d5[71]), .B1(n5667), .C1(n5668[35]), .D1(d4[71]), .CIN(n11608), 
          .S0(d5_71__N_706[70]), .S1(d5_71__N_706[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1097_37.INIT0 = 16'h74b8;
    defparam add_1097_37.INIT1 = 16'h74b8;
    defparam add_1097_37.INJECT1_0 = "NO";
    defparam add_1097_37.INJECT1_1 = "NO";
    CCU2D add_1091_26 (.A0(d3[60]), .B0(d4[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[61]), .B1(d4[61]), .C1(GND_net), .D1(GND_net), .CIN(n11663), 
          .COUT(n11664), .S0(n5516[24]), .S1(n5516[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1091_26.INIT0 = 16'h5666;
    defparam add_1091_26.INIT1 = 16'h5666;
    defparam add_1091_26.INJECT1_0 = "NO";
    defparam add_1091_26.INJECT1_1 = "NO";
    CCU2D add_1097_35 (.A0(d5[68]), .B0(n5667), .C0(n5668[32]), .D0(d4[68]), 
          .A1(d5[69]), .B1(n5667), .C1(n5668[33]), .D1(d4[69]), .CIN(n11607), 
          .COUT(n11608), .S0(d5_71__N_706[68]), .S1(d5_71__N_706[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1097_35.INIT0 = 16'h74b8;
    defparam add_1097_35.INIT1 = 16'h74b8;
    defparam add_1097_35.INJECT1_0 = "NO";
    defparam add_1097_35.INJECT1_1 = "NO";
    CCU2D add_1086_30 (.A0(d2[64]), .B0(d3[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[65]), .B1(d3[65]), .C1(GND_net), .D1(GND_net), .CIN(n11706), 
          .COUT(n11707), .S0(n5364[28]), .S1(n5364[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1086_30.INIT0 = 16'h5666;
    defparam add_1086_30.INIT1 = 16'h5666;
    defparam add_1086_30.INJECT1_0 = "NO";
    defparam add_1086_30.INJECT1_1 = "NO";
    CCU2D add_1086_22 (.A0(d2[56]), .B0(d3[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[57]), .B1(d3[57]), .C1(GND_net), .D1(GND_net), .CIN(n11702), 
          .COUT(n11703), .S0(n5364[20]), .S1(n5364[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1086_22.INIT0 = 16'h5666;
    defparam add_1086_22.INIT1 = 16'h5666;
    defparam add_1086_22.INJECT1_0 = "NO";
    defparam add_1086_22.INJECT1_1 = "NO";
    CCU2D add_1097_13 (.A0(d5[46]), .B0(n5667), .C0(n5668[10]), .D0(d4[46]), 
          .A1(d5[47]), .B1(n5667), .C1(n5668[11]), .D1(d4[47]), .CIN(n11596), 
          .COUT(n11597), .S0(d5_71__N_706[46]), .S1(d5_71__N_706[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1097_13.INIT0 = 16'h74b8;
    defparam add_1097_13.INIT1 = 16'h74b8;
    defparam add_1097_13.INJECT1_0 = "NO";
    defparam add_1097_13.INJECT1_1 = "NO";
    CCU2D add_1086_2 (.A0(d2[36]), .B0(d3[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[37]), .B1(d3[37]), .C1(GND_net), .D1(GND_net), .COUT(n11693), 
          .S1(n5364[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1086_2.INIT0 = 16'h7000;
    defparam add_1086_2.INIT1 = 16'h5666;
    defparam add_1086_2.INJECT1_0 = "NO";
    defparam add_1086_2.INJECT1_1 = "NO";
    CCU2D add_1087_35 (.A0(d3[68]), .B0(n5363), .C0(n5364[32]), .D0(d2[68]), 
          .A1(d3[69]), .B1(n5363), .C1(n5364[33]), .D1(d2[69]), .CIN(n11689), 
          .COUT(n11690), .S0(d3_71__N_562[68]), .S1(d3_71__N_562[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1087_35.INIT0 = 16'h74b8;
    defparam add_1087_35.INIT1 = 16'h74b8;
    defparam add_1087_35.INJECT1_0 = "NO";
    defparam add_1087_35.INJECT1_1 = "NO";
    CCU2D add_1087_33 (.A0(d3[66]), .B0(n5363), .C0(n5364[30]), .D0(d2[66]), 
          .A1(d3[67]), .B1(n5363), .C1(n5364[31]), .D1(d2[67]), .CIN(n11688), 
          .COUT(n11689), .S0(d3_71__N_562[66]), .S1(d3_71__N_562[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1087_33.INIT0 = 16'h74b8;
    defparam add_1087_33.INIT1 = 16'h74b8;
    defparam add_1087_33.INJECT1_0 = "NO";
    defparam add_1087_33.INJECT1_1 = "NO";
    CCU2D add_1097_33 (.A0(d5[66]), .B0(n5667), .C0(n5668[30]), .D0(d4[66]), 
          .A1(d5[67]), .B1(n5667), .C1(n5668[31]), .D1(d4[67]), .CIN(n11606), 
          .COUT(n11607), .S0(d5_71__N_706[66]), .S1(d5_71__N_706[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1097_33.INIT0 = 16'h74b8;
    defparam add_1097_33.INIT1 = 16'h74b8;
    defparam add_1097_33.INJECT1_0 = "NO";
    defparam add_1097_33.INJECT1_1 = "NO";
    CCU2D add_1087_37 (.A0(d3[70]), .B0(n5363), .C0(n5364[34]), .D0(d2[70]), 
          .A1(d3[71]), .B1(n5363), .C1(n5364[35]), .D1(d2[71]), .CIN(n11690), 
          .S0(d3_71__N_562[70]), .S1(d3_71__N_562[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1087_37.INIT0 = 16'h74b8;
    defparam add_1087_37.INIT1 = 16'h74b8;
    defparam add_1087_37.INJECT1_0 = "NO";
    defparam add_1087_37.INJECT1_1 = "NO";
    LUT4 shift_right_31_i62_3_lut (.A(\d10[61] ), .B(\d10[62] ), .C(\CICGain[0] ), 
         .Z(n62)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i62_3_lut.init = 16'hcaca;
    LUT4 i5330_4_lut_rep_115 (.A(n12778), .B(n12503), .C(n12780), .D(count[3]), 
         .Z(n13196)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i5330_4_lut_rep_115.init = 16'h2000;
    CCU2D add_1087_31 (.A0(d3[64]), .B0(n5363), .C0(n5364[28]), .D0(d2[64]), 
          .A1(d3[65]), .B1(n5363), .C1(n5364[29]), .D1(d2[65]), .CIN(n11687), 
          .COUT(n11688), .S0(d3_71__N_562[64]), .S1(d3_71__N_562[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1087_31.INIT0 = 16'h74b8;
    defparam add_1087_31.INIT1 = 16'h74b8;
    defparam add_1087_31.INJECT1_0 = "NO";
    defparam add_1087_31.INJECT1_1 = "NO";
    CCU2D add_1087_23 (.A0(d3[56]), .B0(n5363), .C0(n5364[20]), .D0(d2[56]), 
          .A1(d3[57]), .B1(n5363), .C1(n5364[21]), .D1(d2[57]), .CIN(n11683), 
          .COUT(n11684), .S0(d3_71__N_562[56]), .S1(d3_71__N_562[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1087_23.INIT0 = 16'h74b8;
    defparam add_1087_23.INIT1 = 16'h74b8;
    defparam add_1087_23.INJECT1_0 = "NO";
    defparam add_1087_23.INJECT1_1 = "NO";
    CCU2D add_1087_11 (.A0(d3[44]), .B0(n5363), .C0(n5364[8]), .D0(d2[44]), 
          .A1(d3[45]), .B1(n5363), .C1(n5364[9]), .D1(d2[45]), .CIN(n11677), 
          .COUT(n11678), .S0(d3_71__N_562[44]), .S1(d3_71__N_562[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1087_11.INIT0 = 16'h74b8;
    defparam add_1087_11.INIT1 = 16'h74b8;
    defparam add_1087_11.INJECT1_0 = "NO";
    defparam add_1087_11.INJECT1_1 = "NO";
    CCU2D add_1091_24 (.A0(d3[58]), .B0(d4[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[59]), .B1(d4[59]), .C1(GND_net), .D1(GND_net), .CIN(n11662), 
          .COUT(n11663), .S0(n5516[22]), .S1(n5516[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1091_24.INIT0 = 16'h5666;
    defparam add_1091_24.INIT1 = 16'h5666;
    defparam add_1091_24.INJECT1_0 = "NO";
    defparam add_1091_24.INJECT1_1 = "NO";
    CCU2D add_1087_9 (.A0(d3[42]), .B0(n5363), .C0(n5364[6]), .D0(d2[42]), 
          .A1(d3[43]), .B1(n5363), .C1(n5364[7]), .D1(d2[43]), .CIN(n11676), 
          .COUT(n11677), .S0(d3_71__N_562[42]), .S1(d3_71__N_562[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1087_9.INIT0 = 16'h74b8;
    defparam add_1087_9.INIT1 = 16'h74b8;
    defparam add_1087_9.INJECT1_0 = "NO";
    defparam add_1087_9.INJECT1_1 = "NO";
    CCU2D add_1087_21 (.A0(d3[54]), .B0(n5363), .C0(n5364[18]), .D0(d2[54]), 
          .A1(d3[55]), .B1(n5363), .C1(n5364[19]), .D1(d2[55]), .CIN(n11682), 
          .COUT(n11683), .S0(d3_71__N_562[54]), .S1(d3_71__N_562[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1087_21.INIT0 = 16'h74b8;
    defparam add_1087_21.INIT1 = 16'h74b8;
    defparam add_1087_21.INJECT1_0 = "NO";
    defparam add_1087_21.INJECT1_1 = "NO";
    CCU2D add_1087_7 (.A0(d3[40]), .B0(n5363), .C0(n5364[4]), .D0(d2[40]), 
          .A1(d3[41]), .B1(n5363), .C1(n5364[5]), .D1(d2[41]), .CIN(n11675), 
          .COUT(n11676), .S0(d3_71__N_562[40]), .S1(d3_71__N_562[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1087_7.INIT0 = 16'h74b8;
    defparam add_1087_7.INIT1 = 16'h74b8;
    defparam add_1087_7.INJECT1_0 = "NO";
    defparam add_1087_7.INJECT1_1 = "NO";
    CCU2D add_1087_19 (.A0(d3[52]), .B0(n5363), .C0(n5364[16]), .D0(d2[52]), 
          .A1(d3[53]), .B1(n5363), .C1(n5364[17]), .D1(d2[53]), .CIN(n11681), 
          .COUT(n11682), .S0(d3_71__N_562[52]), .S1(d3_71__N_562[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1087_19.INIT0 = 16'h74b8;
    defparam add_1087_19.INIT1 = 16'h74b8;
    defparam add_1087_19.INJECT1_0 = "NO";
    defparam add_1087_19.INJECT1_1 = "NO";
    CCU2D add_1087_29 (.A0(d3[62]), .B0(n5363), .C0(n5364[26]), .D0(d2[62]), 
          .A1(d3[63]), .B1(n5363), .C1(n5364[27]), .D1(d2[63]), .CIN(n11686), 
          .COUT(n11687), .S0(d3_71__N_562[62]), .S1(d3_71__N_562[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1087_29.INIT0 = 16'h74b8;
    defparam add_1087_29.INIT1 = 16'h74b8;
    defparam add_1087_29.INJECT1_0 = "NO";
    defparam add_1087_29.INJECT1_1 = "NO";
    CCU2D add_1087_17 (.A0(d3[50]), .B0(n5363), .C0(n5364[14]), .D0(d2[50]), 
          .A1(d3[51]), .B1(n5363), .C1(n5364[15]), .D1(d2[51]), .CIN(n11680), 
          .COUT(n11681), .S0(d3_71__N_562[50]), .S1(d3_71__N_562[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1087_17.INIT0 = 16'h74b8;
    defparam add_1087_17.INIT1 = 16'h74b8;
    defparam add_1087_17.INJECT1_0 = "NO";
    defparam add_1087_17.INJECT1_1 = "NO";
    CCU2D add_1087_15 (.A0(d3[48]), .B0(n5363), .C0(n5364[12]), .D0(d2[48]), 
          .A1(d3[49]), .B1(n5363), .C1(n5364[13]), .D1(d2[49]), .CIN(n11679), 
          .COUT(n11680), .S0(d3_71__N_562[48]), .S1(d3_71__N_562[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1087_15.INIT0 = 16'h74b8;
    defparam add_1087_15.INIT1 = 16'h74b8;
    defparam add_1087_15.INJECT1_0 = "NO";
    defparam add_1087_15.INJECT1_1 = "NO";
    CCU2D add_1087_27 (.A0(d3[60]), .B0(n5363), .C0(n5364[24]), .D0(d2[60]), 
          .A1(d3[61]), .B1(n5363), .C1(n5364[25]), .D1(d2[61]), .CIN(n11685), 
          .COUT(n11686), .S0(d3_71__N_562[60]), .S1(d3_71__N_562[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1087_27.INIT0 = 16'h74b8;
    defparam add_1087_27.INIT1 = 16'h74b8;
    defparam add_1087_27.INJECT1_0 = "NO";
    defparam add_1087_27.INJECT1_1 = "NO";
    CCU2D add_1087_13 (.A0(d3[46]), .B0(n5363), .C0(n5364[10]), .D0(d2[46]), 
          .A1(d3[47]), .B1(n5363), .C1(n5364[11]), .D1(d2[47]), .CIN(n11678), 
          .COUT(n11679), .S0(d3_71__N_562[46]), .S1(d3_71__N_562[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1087_13.INIT0 = 16'h74b8;
    defparam add_1087_13.INIT1 = 16'h74b8;
    defparam add_1087_13.INJECT1_0 = "NO";
    defparam add_1087_13.INJECT1_1 = "NO";
    CCU2D add_1087_25 (.A0(d3[58]), .B0(n5363), .C0(n5364[22]), .D0(d2[58]), 
          .A1(d3[59]), .B1(n5363), .C1(n5364[23]), .D1(d2[59]), .CIN(n11684), 
          .COUT(n11685), .S0(d3_71__N_562[58]), .S1(d3_71__N_562[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1087_25.INIT0 = 16'h74b8;
    defparam add_1087_25.INIT1 = 16'h74b8;
    defparam add_1087_25.INJECT1_0 = "NO";
    defparam add_1087_25.INJECT1_1 = "NO";
    CCU2D add_1097_11 (.A0(d5[44]), .B0(n5667), .C0(n5668[8]), .D0(d4[44]), 
          .A1(d5[45]), .B1(n5667), .C1(n5668[9]), .D1(d4[45]), .CIN(n11595), 
          .COUT(n11596), .S0(d5_71__N_706[44]), .S1(d5_71__N_706[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1097_11.INIT0 = 16'h74b8;
    defparam add_1097_11.INIT1 = 16'h74b8;
    defparam add_1097_11.INJECT1_0 = "NO";
    defparam add_1097_11.INJECT1_1 = "NO";
    CCU2D add_1082_13 (.A0(d2[46]), .B0(n5211), .C0(n5212[10]), .D0(d1[46]), 
          .A1(d2[47]), .B1(n5211), .C1(n5212[11]), .D1(d1[47]), .CIN(n11719), 
          .COUT(n11720), .S0(d2_71__N_490[46]), .S1(d2_71__N_490[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1082_13.INIT0 = 16'h74b8;
    defparam add_1082_13.INIT1 = 16'h74b8;
    defparam add_1082_13.INJECT1_0 = "NO";
    defparam add_1082_13.INJECT1_1 = "NO";
    CCU2D add_1081_2 (.A0(d1[36]), .B0(d2[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[37]), .B1(d2[37]), .C1(GND_net), .D1(GND_net), .COUT(n11734), 
          .S1(n5212[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1081_2.INIT0 = 16'h7000;
    defparam add_1081_2.INIT1 = 16'h5666;
    defparam add_1081_2.INJECT1_0 = "NO";
    defparam add_1081_2.INJECT1_1 = "NO";
    LUT4 i2554_2_lut (.A(n375[0]), .B(n31), .Z(count_15__N_1442[0])) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(86[13] 89[16])
    defparam i2554_2_lut.init = 16'hbbbb;
    LUT4 i11_4_lut (.A(count[9]), .B(n22), .C(n18), .D(count[4]), .Z(n31)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i11_4_lut.init = 16'hfffe;
    CCU2D add_1097_9 (.A0(d5[42]), .B0(n5667), .C0(n5668[6]), .D0(d4[42]), 
          .A1(d5[43]), .B1(n5667), .C1(n5668[7]), .D1(d4[43]), .CIN(n11594), 
          .COUT(n11595), .S0(d5_71__N_706[42]), .S1(d5_71__N_706[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1097_9.INIT0 = 16'h74b8;
    defparam add_1097_9.INIT1 = 16'h74b8;
    defparam add_1097_9.INJECT1_0 = "NO";
    defparam add_1097_9.INJECT1_1 = "NO";
    CCU2D add_1097_7 (.A0(d5[40]), .B0(n5667), .C0(n5668[4]), .D0(d4[40]), 
          .A1(d5[41]), .B1(n5667), .C1(n5668[5]), .D1(d4[41]), .CIN(n11593), 
          .COUT(n11594), .S0(d5_71__N_706[40]), .S1(d5_71__N_706[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1097_7.INIT0 = 16'h74b8;
    defparam add_1097_7.INIT1 = 16'h74b8;
    defparam add_1097_7.INJECT1_0 = "NO";
    defparam add_1097_7.INJECT1_1 = "NO";
    CCU2D add_1097_5 (.A0(d5[38]), .B0(n5667), .C0(n5668[2]), .D0(d4[38]), 
          .A1(d5[39]), .B1(n5667), .C1(n5668[3]), .D1(d4[39]), .CIN(n11592), 
          .COUT(n11593), .S0(d5_71__N_706[38]), .S1(d5_71__N_706[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1097_5.INIT0 = 16'h74b8;
    defparam add_1097_5.INIT1 = 16'h74b8;
    defparam add_1097_5.INJECT1_0 = "NO";
    defparam add_1097_5.INJECT1_1 = "NO";
    LUT4 shift_right_31_i63_3_lut (.A(\d10[62] ), .B(\d10[63] ), .C(\CICGain[0] ), 
         .Z(n63)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i63_3_lut.init = 16'hcaca;
    LUT4 i10_4_lut (.A(n19), .B(n15), .C(n12503), .D(count[2]), .Z(n22)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i10_4_lut.init = 16'hfffe;
    CCU2D add_1097_3 (.A0(d5[36]), .B0(n5667), .C0(n5668[0]), .D0(d4[36]), 
          .A1(d5[37]), .B1(n5667), .C1(n5668[1]), .D1(d4[37]), .CIN(n11591), 
          .COUT(n11592), .S0(d5_71__N_706[36]), .S1(d5_71__N_706[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1097_3.INIT0 = 16'h74b8;
    defparam add_1097_3.INIT1 = 16'h74b8;
    defparam add_1097_3.INJECT1_0 = "NO";
    defparam add_1097_3.INJECT1_1 = "NO";
    CCU2D add_1097_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5667), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11591));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1097_1.INIT0 = 16'hF000;
    defparam add_1097_1.INIT1 = 16'h0555;
    defparam add_1097_1.INJECT1_0 = "NO";
    defparam add_1097_1.INJECT1_1 = "NO";
    LUT4 i6_2_lut (.A(count[3]), .B(count[0]), .Z(n18)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 shift_right_31_i64_3_lut (.A(\d10[63] ), .B(\d10[64] ), .C(\CICGain[0] ), 
         .Z(n64)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i64_3_lut.init = 16'hcaca;
    LUT4 i7_4_lut (.A(count[10]), .B(count[1]), .C(count[5]), .D(count[6]), 
         .Z(n19)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[8]), .B(count[7]), .Z(n15)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i3_2_lut.init = 16'heeee;
    LUT4 shift_right_31_i65_3_lut (.A(\d10[64] ), .B(\d10[65] ), .C(\CICGain[0] ), 
         .Z(n65)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i65_3_lut.init = 16'hcaca;
    LUT4 i4631_2_lut (.A(d4[36]), .B(d5[36]), .Z(n5668[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4631_2_lut.init = 16'h6666;
    CCU2D add_1082_37 (.A0(d2[70]), .B0(n5211), .C0(n5212[34]), .D0(d1[70]), 
          .A1(d2[71]), .B1(n5211), .C1(n5212[35]), .D1(d1[71]), .CIN(n11731), 
          .S0(d2_71__N_490[70]), .S1(d2_71__N_490[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1082_37.INIT0 = 16'h74b8;
    defparam add_1082_37.INIT1 = 16'h74b8;
    defparam add_1082_37.INJECT1_0 = "NO";
    defparam add_1082_37.INJECT1_1 = "NO";
    CCU2D add_1082_33 (.A0(d2[66]), .B0(n5211), .C0(n5212[30]), .D0(d1[66]), 
          .A1(d2[67]), .B1(n5211), .C1(n5212[31]), .D1(d1[67]), .CIN(n11729), 
          .COUT(n11730), .S0(d2_71__N_490[66]), .S1(d2_71__N_490[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1082_33.INIT0 = 16'h74b8;
    defparam add_1082_33.INIT1 = 16'h74b8;
    defparam add_1082_33.INJECT1_0 = "NO";
    defparam add_1082_33.INJECT1_1 = "NO";
    CCU2D add_1097_27 (.A0(d5[60]), .B0(n5667), .C0(n5668[24]), .D0(d4[60]), 
          .A1(d5[61]), .B1(n5667), .C1(n5668[25]), .D1(d4[61]), .CIN(n11603), 
          .COUT(n11604), .S0(d5_71__N_706[60]), .S1(d5_71__N_706[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1097_27.INIT0 = 16'h74b8;
    defparam add_1097_27.INIT1 = 16'h74b8;
    defparam add_1097_27.INJECT1_0 = "NO";
    defparam add_1097_27.INJECT1_1 = "NO";
    CCU2D add_1097_31 (.A0(d5[64]), .B0(n5667), .C0(n5668[28]), .D0(d4[64]), 
          .A1(d5[65]), .B1(n5667), .C1(n5668[29]), .D1(d4[65]), .CIN(n11605), 
          .COUT(n11606), .S0(d5_71__N_706[64]), .S1(d5_71__N_706[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1097_31.INIT0 = 16'h74b8;
    defparam add_1097_31.INIT1 = 16'h74b8;
    defparam add_1097_31.INJECT1_0 = "NO";
    defparam add_1097_31.INJECT1_1 = "NO";
    CCU2D add_1082_31 (.A0(d2[64]), .B0(n5211), .C0(n5212[28]), .D0(d1[64]), 
          .A1(d2[65]), .B1(n5211), .C1(n5212[29]), .D1(d1[65]), .CIN(n11728), 
          .COUT(n11729), .S0(d2_71__N_490[64]), .S1(d2_71__N_490[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1082_31.INIT0 = 16'h74b8;
    defparam add_1082_31.INIT1 = 16'h74b8;
    defparam add_1082_31.INJECT1_0 = "NO";
    defparam add_1082_31.INJECT1_1 = "NO";
    CCU2D add_1082_29 (.A0(d2[62]), .B0(n5211), .C0(n5212[26]), .D0(d1[62]), 
          .A1(d2[63]), .B1(n5211), .C1(n5212[27]), .D1(d1[63]), .CIN(n11727), 
          .COUT(n11728), .S0(d2_71__N_490[62]), .S1(d2_71__N_490[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1082_29.INIT0 = 16'h74b8;
    defparam add_1082_29.INIT1 = 16'h74b8;
    defparam add_1082_29.INJECT1_0 = "NO";
    defparam add_1082_29.INJECT1_1 = "NO";
    CCU2D add_1082_27 (.A0(d2[60]), .B0(n5211), .C0(n5212[24]), .D0(d1[60]), 
          .A1(d2[61]), .B1(n5211), .C1(n5212[25]), .D1(d1[61]), .CIN(n11726), 
          .COUT(n11727), .S0(d2_71__N_490[60]), .S1(d2_71__N_490[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1082_27.INIT0 = 16'h74b8;
    defparam add_1082_27.INIT1 = 16'h74b8;
    defparam add_1082_27.INJECT1_0 = "NO";
    defparam add_1082_27.INJECT1_1 = "NO";
    CCU2D add_1082_25 (.A0(d2[58]), .B0(n5211), .C0(n5212[22]), .D0(d1[58]), 
          .A1(d2[59]), .B1(n5211), .C1(n5212[23]), .D1(d1[59]), .CIN(n11725), 
          .COUT(n11726), .S0(d2_71__N_490[58]), .S1(d2_71__N_490[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1082_25.INIT0 = 16'h74b8;
    defparam add_1082_25.INIT1 = 16'h74b8;
    defparam add_1082_25.INJECT1_0 = "NO";
    defparam add_1082_25.INJECT1_1 = "NO";
    CCU2D add_1082_23 (.A0(d2[56]), .B0(n5211), .C0(n5212[20]), .D0(d1[56]), 
          .A1(d2[57]), .B1(n5211), .C1(n5212[21]), .D1(d1[57]), .CIN(n11724), 
          .COUT(n11725), .S0(d2_71__N_490[56]), .S1(d2_71__N_490[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1082_23.INIT0 = 16'h74b8;
    defparam add_1082_23.INIT1 = 16'h74b8;
    defparam add_1082_23.INJECT1_0 = "NO";
    defparam add_1082_23.INJECT1_1 = "NO";
    CCU2D add_1097_23 (.A0(d5[56]), .B0(n5667), .C0(n5668[20]), .D0(d4[56]), 
          .A1(d5[57]), .B1(n5667), .C1(n5668[21]), .D1(d4[57]), .CIN(n11601), 
          .COUT(n11602), .S0(d5_71__N_706[56]), .S1(d5_71__N_706[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1097_23.INIT0 = 16'h74b8;
    defparam add_1097_23.INIT1 = 16'h74b8;
    defparam add_1097_23.INJECT1_0 = "NO";
    defparam add_1097_23.INJECT1_1 = "NO";
    CCU2D add_1111_35 (.A0(d_tmp[69]), .B0(d_d_tmp[69]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[70]), .B1(d_d_tmp[70]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11329), .COUT(n11330), .S0(n6124[33]), 
          .S1(n6124[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1111_35.INIT0 = 16'h5999;
    defparam add_1111_35.INIT1 = 16'h5999;
    defparam add_1111_35.INJECT1_0 = "NO";
    defparam add_1111_35.INJECT1_1 = "NO";
    CCU2D add_1111_33 (.A0(d_tmp[67]), .B0(d_d_tmp[67]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[68]), .B1(d_d_tmp[68]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11328), .COUT(n11329), .S0(n6124[31]), 
          .S1(n6124[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1111_33.INIT0 = 16'h5999;
    defparam add_1111_33.INIT1 = 16'h5999;
    defparam add_1111_33.INJECT1_0 = "NO";
    defparam add_1111_33.INJECT1_1 = "NO";
    CCU2D add_1111_31 (.A0(d_tmp[65]), .B0(d_d_tmp[65]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[66]), .B1(d_d_tmp[66]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11327), .COUT(n11328), .S0(n6124[29]), 
          .S1(n6124[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1111_31.INIT0 = 16'h5999;
    defparam add_1111_31.INIT1 = 16'h5999;
    defparam add_1111_31.INJECT1_0 = "NO";
    defparam add_1111_31.INJECT1_1 = "NO";
    CCU2D add_1111_29 (.A0(d_tmp[63]), .B0(d_d_tmp[63]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[64]), .B1(d_d_tmp[64]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11326), .COUT(n11327), .S0(n6124[27]), 
          .S1(n6124[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1111_29.INIT0 = 16'h5999;
    defparam add_1111_29.INIT1 = 16'h5999;
    defparam add_1111_29.INJECT1_0 = "NO";
    defparam add_1111_29.INJECT1_1 = "NO";
    CCU2D add_1111_27 (.A0(d_tmp[61]), .B0(d_d_tmp[61]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[62]), .B1(d_d_tmp[62]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11325), .COUT(n11326), .S0(n6124[25]), 
          .S1(n6124[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1111_27.INIT0 = 16'h5999;
    defparam add_1111_27.INIT1 = 16'h5999;
    defparam add_1111_27.INJECT1_0 = "NO";
    defparam add_1111_27.INJECT1_1 = "NO";
    CCU2D add_1111_25 (.A0(d_tmp[59]), .B0(d_d_tmp[59]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[60]), .B1(d_d_tmp[60]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11324), .COUT(n11325), .S0(n6124[23]), 
          .S1(n6124[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1111_25.INIT0 = 16'h5999;
    defparam add_1111_25.INIT1 = 16'h5999;
    defparam add_1111_25.INJECT1_0 = "NO";
    defparam add_1111_25.INJECT1_1 = "NO";
    CCU2D add_1111_23 (.A0(d_tmp[57]), .B0(d_d_tmp[57]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[58]), .B1(d_d_tmp[58]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11323), .COUT(n11324), .S0(n6124[21]), 
          .S1(n6124[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1111_23.INIT0 = 16'h5999;
    defparam add_1111_23.INIT1 = 16'h5999;
    defparam add_1111_23.INJECT1_0 = "NO";
    defparam add_1111_23.INJECT1_1 = "NO";
    CCU2D add_1111_21 (.A0(d_tmp[55]), .B0(d_d_tmp[55]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[56]), .B1(d_d_tmp[56]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11322), .COUT(n11323), .S0(n6124[19]), 
          .S1(n6124[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1111_21.INIT0 = 16'h5999;
    defparam add_1111_21.INIT1 = 16'h5999;
    defparam add_1111_21.INJECT1_0 = "NO";
    defparam add_1111_21.INJECT1_1 = "NO";
    CCU2D add_1111_19 (.A0(d_tmp[53]), .B0(d_d_tmp[53]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[54]), .B1(d_d_tmp[54]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11321), .COUT(n11322), .S0(n6124[17]), 
          .S1(n6124[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1111_19.INIT0 = 16'h5999;
    defparam add_1111_19.INIT1 = 16'h5999;
    defparam add_1111_19.INJECT1_0 = "NO";
    defparam add_1111_19.INJECT1_1 = "NO";
    CCU2D add_1086_10 (.A0(d2[44]), .B0(d3[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[45]), .B1(d3[45]), .C1(GND_net), .D1(GND_net), .CIN(n11696), 
          .COUT(n11697), .S0(n5364[8]), .S1(n5364[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1086_10.INIT0 = 16'h5666;
    defparam add_1086_10.INIT1 = 16'h5666;
    defparam add_1086_10.INJECT1_0 = "NO";
    defparam add_1086_10.INJECT1_1 = "NO";
    CCU2D add_1111_17 (.A0(d_tmp[51]), .B0(d_d_tmp[51]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[52]), .B1(d_d_tmp[52]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11320), .COUT(n11321), .S0(n6124[15]), 
          .S1(n6124[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1111_17.INIT0 = 16'h5999;
    defparam add_1111_17.INIT1 = 16'h5999;
    defparam add_1111_17.INJECT1_0 = "NO";
    defparam add_1111_17.INJECT1_1 = "NO";
    CCU2D add_1111_15 (.A0(d_tmp[49]), .B0(d_d_tmp[49]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[50]), .B1(d_d_tmp[50]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11319), .COUT(n11320), .S0(n6124[13]), 
          .S1(n6124[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1111_15.INIT0 = 16'h5999;
    defparam add_1111_15.INIT1 = 16'h5999;
    defparam add_1111_15.INJECT1_0 = "NO";
    defparam add_1111_15.INJECT1_1 = "NO";
    CCU2D add_1111_13 (.A0(d_tmp[47]), .B0(d_d_tmp[47]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[48]), .B1(d_d_tmp[48]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11318), .COUT(n11319), .S0(n6124[11]), 
          .S1(n6124[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1111_13.INIT0 = 16'h5999;
    defparam add_1111_13.INIT1 = 16'h5999;
    defparam add_1111_13.INJECT1_0 = "NO";
    defparam add_1111_13.INJECT1_1 = "NO";
    CCU2D add_1091_22 (.A0(d3[56]), .B0(d4[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[57]), .B1(d4[57]), .C1(GND_net), .D1(GND_net), .CIN(n11661), 
          .COUT(n11662), .S0(n5516[20]), .S1(n5516[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1091_22.INIT0 = 16'h5666;
    defparam add_1091_22.INIT1 = 16'h5666;
    defparam add_1091_22.INJECT1_0 = "NO";
    defparam add_1091_22.INJECT1_1 = "NO";
    CCU2D add_1091_20 (.A0(d3[54]), .B0(d4[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[55]), .B1(d4[55]), .C1(GND_net), .D1(GND_net), .CIN(n11660), 
          .COUT(n11661), .S0(n5516[18]), .S1(n5516[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1091_20.INIT0 = 16'h5666;
    defparam add_1091_20.INIT1 = 16'h5666;
    defparam add_1091_20.INJECT1_0 = "NO";
    defparam add_1091_20.INJECT1_1 = "NO";
    CCU2D add_1086_8 (.A0(d2[42]), .B0(d3[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[43]), .B1(d3[43]), .C1(GND_net), .D1(GND_net), .CIN(n11695), 
          .COUT(n11696), .S0(n5364[6]), .S1(n5364[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1086_8.INIT0 = 16'h5666;
    defparam add_1086_8.INIT1 = 16'h5666;
    defparam add_1086_8.INJECT1_0 = "NO";
    defparam add_1086_8.INJECT1_1 = "NO";
    LUT4 shift_right_31_i66_3_lut (.A(\d10[65] ), .B(\d10[66] ), .C(\CICGain[0] ), 
         .Z(n66)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i66_3_lut.init = 16'hcaca;
    CCU2D add_1097_29 (.A0(d5[62]), .B0(n5667), .C0(n5668[26]), .D0(d4[62]), 
          .A1(d5[63]), .B1(n5667), .C1(n5668[27]), .D1(d4[63]), .CIN(n11604), 
          .COUT(n11605), .S0(d5_71__N_706[62]), .S1(d5_71__N_706[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1097_29.INIT0 = 16'h74b8;
    defparam add_1097_29.INIT1 = 16'h74b8;
    defparam add_1097_29.INJECT1_0 = "NO";
    defparam add_1097_29.INJECT1_1 = "NO";
    CCU2D add_1091_18 (.A0(d3[52]), .B0(d4[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[53]), .B1(d4[53]), .C1(GND_net), .D1(GND_net), .CIN(n11659), 
          .COUT(n11660), .S0(n5516[16]), .S1(n5516[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1091_18.INIT0 = 16'h5666;
    defparam add_1091_18.INIT1 = 16'h5666;
    defparam add_1091_18.INJECT1_0 = "NO";
    defparam add_1091_18.INJECT1_1 = "NO";
    CCU2D add_1086_20 (.A0(d2[54]), .B0(d3[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[55]), .B1(d3[55]), .C1(GND_net), .D1(GND_net), .CIN(n11701), 
          .COUT(n11702), .S0(n5364[18]), .S1(n5364[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1086_20.INIT0 = 16'h5666;
    defparam add_1086_20.INIT1 = 16'h5666;
    defparam add_1086_20.INJECT1_0 = "NO";
    defparam add_1086_20.INJECT1_1 = "NO";
    CCU2D add_1086_6 (.A0(d2[40]), .B0(d3[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[41]), .B1(d3[41]), .C1(GND_net), .D1(GND_net), .CIN(n11694), 
          .COUT(n11695), .S0(n5364[4]), .S1(n5364[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1086_6.INIT0 = 16'h5666;
    defparam add_1086_6.INIT1 = 16'h5666;
    defparam add_1086_6.INJECT1_0 = "NO";
    defparam add_1086_6.INJECT1_1 = "NO";
    CCU2D add_1086_18 (.A0(d2[52]), .B0(d3[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[53]), .B1(d3[53]), .C1(GND_net), .D1(GND_net), .CIN(n11700), 
          .COUT(n11701), .S0(n5364[16]), .S1(n5364[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1086_18.INIT0 = 16'h5666;
    defparam add_1086_18.INIT1 = 16'h5666;
    defparam add_1086_18.INJECT1_0 = "NO";
    defparam add_1086_18.INJECT1_1 = "NO";
    CCU2D add_1086_28 (.A0(d2[62]), .B0(d3[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[63]), .B1(d3[63]), .C1(GND_net), .D1(GND_net), .CIN(n11705), 
          .COUT(n11706), .S0(n5364[26]), .S1(n5364[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1086_28.INIT0 = 16'h5666;
    defparam add_1086_28.INIT1 = 16'h5666;
    defparam add_1086_28.INJECT1_0 = "NO";
    defparam add_1086_28.INJECT1_1 = "NO";
    CCU2D add_1086_16 (.A0(d2[50]), .B0(d3[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[51]), .B1(d3[51]), .C1(GND_net), .D1(GND_net), .CIN(n11699), 
          .COUT(n11700), .S0(n5364[14]), .S1(n5364[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1086_16.INIT0 = 16'h5666;
    defparam add_1086_16.INIT1 = 16'h5666;
    defparam add_1086_16.INJECT1_0 = "NO";
    defparam add_1086_16.INJECT1_1 = "NO";
    CCU2D add_1086_4 (.A0(d2[38]), .B0(d3[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[39]), .B1(d3[39]), .C1(GND_net), .D1(GND_net), .CIN(n11693), 
          .COUT(n11694), .S0(n5364[2]), .S1(n5364[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1086_4.INIT0 = 16'h5666;
    defparam add_1086_4.INIT1 = 16'h5666;
    defparam add_1086_4.INJECT1_0 = "NO";
    defparam add_1086_4.INJECT1_1 = "NO";
    CCU2D add_1086_14 (.A0(d2[48]), .B0(d3[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[49]), .B1(d3[49]), .C1(GND_net), .D1(GND_net), .CIN(n11698), 
          .COUT(n11699), .S0(n5364[12]), .S1(n5364[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1086_14.INIT0 = 16'h5666;
    defparam add_1086_14.INIT1 = 16'h5666;
    defparam add_1086_14.INJECT1_0 = "NO";
    defparam add_1086_14.INJECT1_1 = "NO";
    LUT4 i4_4_lut (.A(n7), .B(count[15]), .C(count[11]), .D(count[14]), 
         .Z(n12503)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i4_4_lut.init = 16'hffef;
    LUT4 shift_right_31_i61_3_lut (.A(\d10[60] ), .B(\d10[61] ), .C(\CICGain[0] ), 
         .Z(n61)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i61_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i67_3_lut (.A(\d10[66] ), .B(\d10[67] ), .C(\CICGain[0] ), 
         .Z(n67)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i67_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut (.A(count[13]), .B(count[12]), .Z(n7)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    CCU2D add_1086_26 (.A0(d2[60]), .B0(d3[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[61]), .B1(d3[61]), .C1(GND_net), .D1(GND_net), .CIN(n11704), 
          .COUT(n11705), .S0(n5364[24]), .S1(n5364[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1086_26.INIT0 = 16'h5666;
    defparam add_1086_26.INIT1 = 16'h5666;
    defparam add_1086_26.INJECT1_0 = "NO";
    defparam add_1086_26.INJECT1_1 = "NO";
    CCU2D add_1081_34 (.A0(d1[68]), .B0(d2[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[69]), .B1(d2[69]), .C1(GND_net), .D1(GND_net), .CIN(n11749), 
          .COUT(n11750), .S0(n5212[32]), .S1(n5212[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1081_34.INIT0 = 16'h5666;
    defparam add_1081_34.INIT1 = 16'h5666;
    defparam add_1081_34.INJECT1_0 = "NO";
    defparam add_1081_34.INJECT1_1 = "NO";
    CCU2D add_1081_32 (.A0(d1[66]), .B0(d2[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[67]), .B1(d2[67]), .C1(GND_net), .D1(GND_net), .CIN(n11748), 
          .COUT(n11749), .S0(n5212[30]), .S1(n5212[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1081_32.INIT0 = 16'h5666;
    defparam add_1081_32.INIT1 = 16'h5666;
    defparam add_1081_32.INJECT1_0 = "NO";
    defparam add_1081_32.INJECT1_1 = "NO";
    CCU2D add_1082_21 (.A0(d2[54]), .B0(n5211), .C0(n5212[18]), .D0(d1[54]), 
          .A1(d2[55]), .B1(n5211), .C1(n5212[19]), .D1(d1[55]), .CIN(n11723), 
          .COUT(n11724), .S0(d2_71__N_490[54]), .S1(d2_71__N_490[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1082_21.INIT0 = 16'h74b8;
    defparam add_1082_21.INIT1 = 16'h74b8;
    defparam add_1082_21.INJECT1_0 = "NO";
    defparam add_1082_21.INJECT1_1 = "NO";
    LUT4 shift_right_31_i68_3_lut (.A(\d10[67] ), .B(\d10[68] ), .C(\CICGain[0] ), 
         .Z(n68)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i68_3_lut.init = 16'hcaca;
    CCU2D add_1091_16 (.A0(d3[50]), .B0(d4[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[51]), .B1(d4[51]), .C1(GND_net), .D1(GND_net), .CIN(n11658), 
          .COUT(n11659), .S0(n5516[14]), .S1(n5516[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1091_16.INIT0 = 16'h5666;
    defparam add_1091_16.INIT1 = 16'h5666;
    defparam add_1091_16.INJECT1_0 = "NO";
    defparam add_1091_16.INJECT1_1 = "NO";
    CCU2D add_1082_17 (.A0(d2[50]), .B0(n5211), .C0(n5212[14]), .D0(d1[50]), 
          .A1(d2[51]), .B1(n5211), .C1(n5212[15]), .D1(d1[51]), .CIN(n11721), 
          .COUT(n11722), .S0(d2_71__N_490[50]), .S1(d2_71__N_490[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1082_17.INIT0 = 16'h74b8;
    defparam add_1082_17.INIT1 = 16'h74b8;
    defparam add_1082_17.INJECT1_0 = "NO";
    defparam add_1082_17.INJECT1_1 = "NO";
    CCU2D add_1082_15 (.A0(d2[48]), .B0(n5211), .C0(n5212[12]), .D0(d1[48]), 
          .A1(d2[49]), .B1(n5211), .C1(n5212[13]), .D1(d1[49]), .CIN(n11720), 
          .COUT(n11721), .S0(d2_71__N_490[48]), .S1(d2_71__N_490[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1082_15.INIT0 = 16'h74b8;
    defparam add_1082_15.INIT1 = 16'h74b8;
    defparam add_1082_15.INJECT1_0 = "NO";
    defparam add_1082_15.INJECT1_1 = "NO";
    CCU2D add_1082_19 (.A0(d2[52]), .B0(n5211), .C0(n5212[16]), .D0(d1[52]), 
          .A1(d2[53]), .B1(n5211), .C1(n5212[17]), .D1(d1[53]), .CIN(n11722), 
          .COUT(n11723), .S0(d2_71__N_490[52]), .S1(d2_71__N_490[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1082_19.INIT0 = 16'h74b8;
    defparam add_1082_19.INIT1 = 16'h74b8;
    defparam add_1082_19.INJECT1_0 = "NO";
    defparam add_1082_19.INJECT1_1 = "NO";
    CCU2D add_1081_30 (.A0(d1[64]), .B0(d2[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[65]), .B1(d2[65]), .C1(GND_net), .D1(GND_net), .CIN(n11747), 
          .COUT(n11748), .S0(n5212[28]), .S1(n5212[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1081_30.INIT0 = 16'h5666;
    defparam add_1081_30.INIT1 = 16'h5666;
    defparam add_1081_30.INJECT1_0 = "NO";
    defparam add_1081_30.INJECT1_1 = "NO";
    CCU2D add_1086_12 (.A0(d2[46]), .B0(d3[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[47]), .B1(d3[47]), .C1(GND_net), .D1(GND_net), .CIN(n11697), 
          .COUT(n11698), .S0(n5364[10]), .S1(n5364[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1086_12.INIT0 = 16'h5666;
    defparam add_1086_12.INIT1 = 16'h5666;
    defparam add_1086_12.INJECT1_0 = "NO";
    defparam add_1086_12.INJECT1_1 = "NO";
    CCU2D add_1086_24 (.A0(d2[58]), .B0(d3[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[59]), .B1(d3[59]), .C1(GND_net), .D1(GND_net), .CIN(n11703), 
          .COUT(n11704), .S0(n5364[22]), .S1(n5364[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1086_24.INIT0 = 16'h5666;
    defparam add_1086_24.INIT1 = 16'h5666;
    defparam add_1086_24.INJECT1_0 = "NO";
    defparam add_1086_24.INJECT1_1 = "NO";
    CCU2D add_1081_28 (.A0(d1[62]), .B0(d2[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[63]), .B1(d2[63]), .C1(GND_net), .D1(GND_net), .CIN(n11746), 
          .COUT(n11747), .S0(n5212[26]), .S1(n5212[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1081_28.INIT0 = 16'h5666;
    defparam add_1081_28.INIT1 = 16'h5666;
    defparam add_1081_28.INJECT1_0 = "NO";
    defparam add_1081_28.INJECT1_1 = "NO";
    CCU2D add_1081_26 (.A0(d1[60]), .B0(d2[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[61]), .B1(d2[61]), .C1(GND_net), .D1(GND_net), .CIN(n11745), 
          .COUT(n11746), .S0(n5212[24]), .S1(n5212[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1081_26.INIT0 = 16'h5666;
    defparam add_1081_26.INIT1 = 16'h5666;
    defparam add_1081_26.INJECT1_0 = "NO";
    defparam add_1081_26.INJECT1_1 = "NO";
    LUT4 i4601_2_lut (.A(MixerOutCos[0]), .B(d1[0]), .Z(d1_71__N_418[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4601_2_lut.init = 16'h6666;
    CCU2D add_1091_14 (.A0(d3[48]), .B0(d4[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[49]), .B1(d4[49]), .C1(GND_net), .D1(GND_net), .CIN(n11657), 
          .COUT(n11658), .S0(n5516[12]), .S1(n5516[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1091_14.INIT0 = 16'h5666;
    defparam add_1091_14.INIT1 = 16'h5666;
    defparam add_1091_14.INJECT1_0 = "NO";
    defparam add_1091_14.INJECT1_1 = "NO";
    CCU2D add_1091_12 (.A0(d3[46]), .B0(d4[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[47]), .B1(d4[47]), .C1(GND_net), .D1(GND_net), .CIN(n11656), 
          .COUT(n11657), .S0(n5516[10]), .S1(n5516[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1091_12.INIT0 = 16'h5666;
    defparam add_1091_12.INIT1 = 16'h5666;
    defparam add_1091_12.INJECT1_0 = "NO";
    defparam add_1091_12.INJECT1_1 = "NO";
    CCU2D add_1091_10 (.A0(d3[44]), .B0(d4[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[45]), .B1(d4[45]), .C1(GND_net), .D1(GND_net), .CIN(n11655), 
          .COUT(n11656), .S0(n5516[8]), .S1(n5516[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1091_10.INIT0 = 16'h5666;
    defparam add_1091_10.INIT1 = 16'h5666;
    defparam add_1091_10.INJECT1_0 = "NO";
    defparam add_1091_10.INJECT1_1 = "NO";
    CCU2D add_1091_8 (.A0(d3[42]), .B0(d4[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[43]), .B1(d4[43]), .C1(GND_net), .D1(GND_net), .CIN(n11654), 
          .COUT(n11655), .S0(n5516[6]), .S1(n5516[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1091_8.INIT0 = 16'h5666;
    defparam add_1091_8.INIT1 = 16'h5666;
    defparam add_1091_8.INJECT1_0 = "NO";
    defparam add_1091_8.INJECT1_1 = "NO";
    CCU2D add_1091_6 (.A0(d3[40]), .B0(d4[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[41]), .B1(d4[41]), .C1(GND_net), .D1(GND_net), .CIN(n11653), 
          .COUT(n11654), .S0(n5516[4]), .S1(n5516[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1091_6.INIT0 = 16'h5666;
    defparam add_1091_6.INIT1 = 16'h5666;
    defparam add_1091_6.INJECT1_0 = "NO";
    defparam add_1091_6.INJECT1_1 = "NO";
    CCU2D add_1091_4 (.A0(d3[38]), .B0(d4[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[39]), .B1(d4[39]), .C1(GND_net), .D1(GND_net), .CIN(n11652), 
          .COUT(n11653), .S0(n5516[2]), .S1(n5516[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1091_4.INIT0 = 16'h5666;
    defparam add_1091_4.INIT1 = 16'h5666;
    defparam add_1091_4.INJECT1_0 = "NO";
    defparam add_1091_4.INJECT1_1 = "NO";
    CCU2D add_1091_2 (.A0(d3[36]), .B0(d4[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[37]), .B1(d4[37]), .C1(GND_net), .D1(GND_net), .COUT(n11652), 
          .S1(n5516[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1091_2.INIT0 = 16'h7000;
    defparam add_1091_2.INIT1 = 16'h5666;
    defparam add_1091_2.INJECT1_0 = "NO";
    defparam add_1091_2.INJECT1_1 = "NO";
    LUT4 shift_right_31_i70_3_lut (.A(\d10[69] ), .B(\d10[70] ), .C(\CICGain[0] ), 
         .Z(n70)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i70_3_lut.init = 16'hcaca;
    CCU2D add_1111_11 (.A0(d_tmp[45]), .B0(d_d_tmp[45]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[46]), .B1(d_d_tmp[46]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11317), .COUT(n11318), .S0(n6124[9]), 
          .S1(n6124[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1111_11.INIT0 = 16'h5999;
    defparam add_1111_11.INIT1 = 16'h5999;
    defparam add_1111_11.INJECT1_0 = "NO";
    defparam add_1111_11.INJECT1_1 = "NO";
    CCU2D add_1092_37 (.A0(d4[70]), .B0(n5515), .C0(n5516[34]), .D0(d3[70]), 
          .A1(d4[71]), .B1(n5515), .C1(n5516[35]), .D1(d3[71]), .CIN(n11649), 
          .S0(d4_71__N_634[70]), .S1(d4_71__N_634[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1092_37.INIT0 = 16'h74b8;
    defparam add_1092_37.INIT1 = 16'h74b8;
    defparam add_1092_37.INJECT1_0 = "NO";
    defparam add_1092_37.INJECT1_1 = "NO";
    CCU2D add_1092_35 (.A0(d4[68]), .B0(n5515), .C0(n5516[32]), .D0(d3[68]), 
          .A1(d4[69]), .B1(n5515), .C1(n5516[33]), .D1(d3[69]), .CIN(n11648), 
          .COUT(n11649), .S0(d4_71__N_634[68]), .S1(d4_71__N_634[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1092_35.INIT0 = 16'h74b8;
    defparam add_1092_35.INIT1 = 16'h74b8;
    defparam add_1092_35.INJECT1_0 = "NO";
    defparam add_1092_35.INJECT1_1 = "NO";
    CCU2D add_1092_33 (.A0(d4[66]), .B0(n5515), .C0(n5516[30]), .D0(d3[66]), 
          .A1(d4[67]), .B1(n5515), .C1(n5516[31]), .D1(d3[67]), .CIN(n11647), 
          .COUT(n11648), .S0(d4_71__N_634[66]), .S1(d4_71__N_634[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1092_33.INIT0 = 16'h74b8;
    defparam add_1092_33.INIT1 = 16'h74b8;
    defparam add_1092_33.INJECT1_0 = "NO";
    defparam add_1092_33.INJECT1_1 = "NO";
    CCU2D add_1092_31 (.A0(d4[64]), .B0(n5515), .C0(n5516[28]), .D0(d3[64]), 
          .A1(d4[65]), .B1(n5515), .C1(n5516[29]), .D1(d3[65]), .CIN(n11646), 
          .COUT(n11647), .S0(d4_71__N_634[64]), .S1(d4_71__N_634[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1092_31.INIT0 = 16'h74b8;
    defparam add_1092_31.INIT1 = 16'h74b8;
    defparam add_1092_31.INJECT1_0 = "NO";
    defparam add_1092_31.INJECT1_1 = "NO";
    CCU2D add_1092_29 (.A0(d4[62]), .B0(n5515), .C0(n5516[26]), .D0(d3[62]), 
          .A1(d4[63]), .B1(n5515), .C1(n5516[27]), .D1(d3[63]), .CIN(n11645), 
          .COUT(n11646), .S0(d4_71__N_634[62]), .S1(d4_71__N_634[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1092_29.INIT0 = 16'h74b8;
    defparam add_1092_29.INIT1 = 16'h74b8;
    defparam add_1092_29.INJECT1_0 = "NO";
    defparam add_1092_29.INJECT1_1 = "NO";
    CCU2D add_1092_27 (.A0(d4[60]), .B0(n5515), .C0(n5516[24]), .D0(d3[60]), 
          .A1(d4[61]), .B1(n5515), .C1(n5516[25]), .D1(d3[61]), .CIN(n11644), 
          .COUT(n11645), .S0(d4_71__N_634[60]), .S1(d4_71__N_634[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1092_27.INIT0 = 16'h74b8;
    defparam add_1092_27.INIT1 = 16'h74b8;
    defparam add_1092_27.INJECT1_0 = "NO";
    defparam add_1092_27.INJECT1_1 = "NO";
    CCU2D add_1092_25 (.A0(d4[58]), .B0(n5515), .C0(n5516[22]), .D0(d3[58]), 
          .A1(d4[59]), .B1(n5515), .C1(n5516[23]), .D1(d3[59]), .CIN(n11643), 
          .COUT(n11644), .S0(d4_71__N_634[58]), .S1(d4_71__N_634[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1092_25.INIT0 = 16'h74b8;
    defparam add_1092_25.INIT1 = 16'h74b8;
    defparam add_1092_25.INJECT1_0 = "NO";
    defparam add_1092_25.INJECT1_1 = "NO";
    LUT4 i4637_2_lut (.A(d2[36]), .B(d3[36]), .Z(n5364[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4637_2_lut.init = 16'h6666;
    CCU2D add_1092_23 (.A0(d4[56]), .B0(n5515), .C0(n5516[20]), .D0(d3[56]), 
          .A1(d4[57]), .B1(n5515), .C1(n5516[21]), .D1(d3[57]), .CIN(n11642), 
          .COUT(n11643), .S0(d4_71__N_634[56]), .S1(d4_71__N_634[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1092_23.INIT0 = 16'h74b8;
    defparam add_1092_23.INIT1 = 16'h74b8;
    defparam add_1092_23.INJECT1_0 = "NO";
    defparam add_1092_23.INJECT1_1 = "NO";
    CCU2D add_1092_21 (.A0(d4[54]), .B0(n5515), .C0(n5516[18]), .D0(d3[54]), 
          .A1(d4[55]), .B1(n5515), .C1(n5516[19]), .D1(d3[55]), .CIN(n11641), 
          .COUT(n11642), .S0(d4_71__N_634[54]), .S1(d4_71__N_634[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1092_21.INIT0 = 16'h74b8;
    defparam add_1092_21.INIT1 = 16'h74b8;
    defparam add_1092_21.INJECT1_0 = "NO";
    defparam add_1092_21.INJECT1_1 = "NO";
    CCU2D add_1092_19 (.A0(d4[52]), .B0(n5515), .C0(n5516[16]), .D0(d3[52]), 
          .A1(d4[53]), .B1(n5515), .C1(n5516[17]), .D1(d3[53]), .CIN(n11640), 
          .COUT(n11641), .S0(d4_71__N_634[52]), .S1(d4_71__N_634[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1092_19.INIT0 = 16'h74b8;
    defparam add_1092_19.INIT1 = 16'h74b8;
    defparam add_1092_19.INJECT1_0 = "NO";
    defparam add_1092_19.INJECT1_1 = "NO";
    CCU2D add_1092_17 (.A0(d4[50]), .B0(n5515), .C0(n5516[14]), .D0(d3[50]), 
          .A1(d4[51]), .B1(n5515), .C1(n5516[15]), .D1(d3[51]), .CIN(n11639), 
          .COUT(n11640), .S0(d4_71__N_634[50]), .S1(d4_71__N_634[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1092_17.INIT0 = 16'h74b8;
    defparam add_1092_17.INIT1 = 16'h74b8;
    defparam add_1092_17.INJECT1_0 = "NO";
    defparam add_1092_17.INJECT1_1 = "NO";
    CCU2D add_1092_15 (.A0(d4[48]), .B0(n5515), .C0(n5516[12]), .D0(d3[48]), 
          .A1(d4[49]), .B1(n5515), .C1(n5516[13]), .D1(d3[49]), .CIN(n11638), 
          .COUT(n11639), .S0(d4_71__N_634[48]), .S1(d4_71__N_634[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1092_15.INIT0 = 16'h74b8;
    defparam add_1092_15.INIT1 = 16'h74b8;
    defparam add_1092_15.INJECT1_0 = "NO";
    defparam add_1092_15.INJECT1_1 = "NO";
    CCU2D add_1092_13 (.A0(d4[46]), .B0(n5515), .C0(n5516[10]), .D0(d3[46]), 
          .A1(d4[47]), .B1(n5515), .C1(n5516[11]), .D1(d3[47]), .CIN(n11637), 
          .COUT(n11638), .S0(d4_71__N_634[46]), .S1(d4_71__N_634[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1092_13.INIT0 = 16'h74b8;
    defparam add_1092_13.INIT1 = 16'h74b8;
    defparam add_1092_13.INJECT1_0 = "NO";
    defparam add_1092_13.INJECT1_1 = "NO";
    CCU2D add_1092_11 (.A0(d4[44]), .B0(n5515), .C0(n5516[8]), .D0(d3[44]), 
          .A1(d4[45]), .B1(n5515), .C1(n5516[9]), .D1(d3[45]), .CIN(n11636), 
          .COUT(n11637), .S0(d4_71__N_634[44]), .S1(d4_71__N_634[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1092_11.INIT0 = 16'h74b8;
    defparam add_1092_11.INIT1 = 16'h74b8;
    defparam add_1092_11.INJECT1_0 = "NO";
    defparam add_1092_11.INJECT1_1 = "NO";
    CCU2D add_1092_9 (.A0(d4[42]), .B0(n5515), .C0(n5516[6]), .D0(d3[42]), 
          .A1(d4[43]), .B1(n5515), .C1(n5516[7]), .D1(d3[43]), .CIN(n11635), 
          .COUT(n11636), .S0(d4_71__N_634[42]), .S1(d4_71__N_634[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1092_9.INIT0 = 16'h74b8;
    defparam add_1092_9.INIT1 = 16'h74b8;
    defparam add_1092_9.INJECT1_0 = "NO";
    defparam add_1092_9.INJECT1_1 = "NO";
    CCU2D add_1092_7 (.A0(d4[40]), .B0(n5515), .C0(n5516[4]), .D0(d3[40]), 
          .A1(d4[41]), .B1(n5515), .C1(n5516[5]), .D1(d3[41]), .CIN(n11634), 
          .COUT(n11635), .S0(d4_71__N_634[40]), .S1(d4_71__N_634[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1092_7.INIT0 = 16'h74b8;
    defparam add_1092_7.INIT1 = 16'h74b8;
    defparam add_1092_7.INJECT1_0 = "NO";
    defparam add_1092_7.INJECT1_1 = "NO";
    CCU2D add_1092_5 (.A0(d4[38]), .B0(n5515), .C0(n5516[2]), .D0(d3[38]), 
          .A1(d4[39]), .B1(n5515), .C1(n5516[3]), .D1(d3[39]), .CIN(n11633), 
          .COUT(n11634), .S0(d4_71__N_634[38]), .S1(d4_71__N_634[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1092_5.INIT0 = 16'h74b8;
    defparam add_1092_5.INIT1 = 16'h74b8;
    defparam add_1092_5.INJECT1_0 = "NO";
    defparam add_1092_5.INJECT1_1 = "NO";
    CCU2D add_1092_3 (.A0(d4[36]), .B0(n5515), .C0(n5516[0]), .D0(d3[36]), 
          .A1(d4[37]), .B1(n5515), .C1(n5516[1]), .D1(d3[37]), .CIN(n11632), 
          .COUT(n11633), .S0(d4_71__N_634[36]), .S1(d4_71__N_634[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1092_3.INIT0 = 16'h74b8;
    defparam add_1092_3.INIT1 = 16'h74b8;
    defparam add_1092_3.INJECT1_0 = "NO";
    defparam add_1092_3.INJECT1_1 = "NO";
    CCU2D add_1092_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5515), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11632));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1092_1.INIT0 = 16'hF000;
    defparam add_1092_1.INIT1 = 16'h0555;
    defparam add_1092_1.INJECT1_0 = "NO";
    defparam add_1092_1.INJECT1_1 = "NO";
    CCU2D add_1096_36 (.A0(d4[70]), .B0(d5[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[71]), .B1(d5[71]), .C1(GND_net), .D1(GND_net), .CIN(n11627), 
          .S0(n5668[34]), .S1(n5668[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1096_36.INIT0 = 16'h5666;
    defparam add_1096_36.INIT1 = 16'h5666;
    defparam add_1096_36.INJECT1_0 = "NO";
    defparam add_1096_36.INJECT1_1 = "NO";
    CCU2D add_1096_34 (.A0(d4[68]), .B0(d5[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[69]), .B1(d5[69]), .C1(GND_net), .D1(GND_net), .CIN(n11626), 
          .COUT(n11627), .S0(n5668[32]), .S1(n5668[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1096_34.INIT0 = 16'h5666;
    defparam add_1096_34.INIT1 = 16'h5666;
    defparam add_1096_34.INJECT1_0 = "NO";
    defparam add_1096_34.INJECT1_1 = "NO";
    CCU2D add_1096_32 (.A0(d4[66]), .B0(d5[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[67]), .B1(d5[67]), .C1(GND_net), .D1(GND_net), .CIN(n11625), 
          .COUT(n11626), .S0(n5668[30]), .S1(n5668[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1096_32.INIT0 = 16'h5666;
    defparam add_1096_32.INIT1 = 16'h5666;
    defparam add_1096_32.INJECT1_0 = "NO";
    defparam add_1096_32.INJECT1_1 = "NO";
    CCU2D add_1096_30 (.A0(d4[64]), .B0(d5[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[65]), .B1(d5[65]), .C1(GND_net), .D1(GND_net), .CIN(n11624), 
          .COUT(n11625), .S0(n5668[28]), .S1(n5668[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1096_30.INIT0 = 16'h5666;
    defparam add_1096_30.INIT1 = 16'h5666;
    defparam add_1096_30.INJECT1_0 = "NO";
    defparam add_1096_30.INJECT1_1 = "NO";
    CCU2D add_1096_28 (.A0(d4[62]), .B0(d5[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[63]), .B1(d5[63]), .C1(GND_net), .D1(GND_net), .CIN(n11623), 
          .COUT(n11624), .S0(n5668[26]), .S1(n5668[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1096_28.INIT0 = 16'h5666;
    defparam add_1096_28.INIT1 = 16'h5666;
    defparam add_1096_28.INJECT1_0 = "NO";
    defparam add_1096_28.INJECT1_1 = "NO";
    CCU2D add_1096_26 (.A0(d4[60]), .B0(d5[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[61]), .B1(d5[61]), .C1(GND_net), .D1(GND_net), .CIN(n11622), 
          .COUT(n11623), .S0(n5668[24]), .S1(n5668[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1096_26.INIT0 = 16'h5666;
    defparam add_1096_26.INIT1 = 16'h5666;
    defparam add_1096_26.INJECT1_0 = "NO";
    defparam add_1096_26.INJECT1_1 = "NO";
    CCU2D add_1096_24 (.A0(d4[58]), .B0(d5[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[59]), .B1(d5[59]), .C1(GND_net), .D1(GND_net), .CIN(n11621), 
          .COUT(n11622), .S0(n5668[22]), .S1(n5668[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1096_24.INIT0 = 16'h5666;
    defparam add_1096_24.INIT1 = 16'h5666;
    defparam add_1096_24.INJECT1_0 = "NO";
    defparam add_1096_24.INJECT1_1 = "NO";
    CCU2D add_1096_22 (.A0(d4[56]), .B0(d5[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[57]), .B1(d5[57]), .C1(GND_net), .D1(GND_net), .CIN(n11620), 
          .COUT(n11621), .S0(n5668[20]), .S1(n5668[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1096_22.INIT0 = 16'h5666;
    defparam add_1096_22.INIT1 = 16'h5666;
    defparam add_1096_22.INJECT1_0 = "NO";
    defparam add_1096_22.INJECT1_1 = "NO";
    CCU2D add_1096_20 (.A0(d4[54]), .B0(d5[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[55]), .B1(d5[55]), .C1(GND_net), .D1(GND_net), .CIN(n11619), 
          .COUT(n11620), .S0(n5668[18]), .S1(n5668[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1096_20.INIT0 = 16'h5666;
    defparam add_1096_20.INIT1 = 16'h5666;
    defparam add_1096_20.INJECT1_0 = "NO";
    defparam add_1096_20.INJECT1_1 = "NO";
    CCU2D add_1096_18 (.A0(d4[52]), .B0(d5[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[53]), .B1(d5[53]), .C1(GND_net), .D1(GND_net), .CIN(n11618), 
          .COUT(n11619), .S0(n5668[16]), .S1(n5668[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1096_18.INIT0 = 16'h5666;
    defparam add_1096_18.INIT1 = 16'h5666;
    defparam add_1096_18.INJECT1_0 = "NO";
    defparam add_1096_18.INJECT1_1 = "NO";
    CCU2D add_1096_16 (.A0(d4[50]), .B0(d5[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[51]), .B1(d5[51]), .C1(GND_net), .D1(GND_net), .CIN(n11617), 
          .COUT(n11618), .S0(n5668[14]), .S1(n5668[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1096_16.INIT0 = 16'h5666;
    defparam add_1096_16.INIT1 = 16'h5666;
    defparam add_1096_16.INJECT1_0 = "NO";
    defparam add_1096_16.INJECT1_1 = "NO";
    CCU2D add_1096_14 (.A0(d4[48]), .B0(d5[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[49]), .B1(d5[49]), .C1(GND_net), .D1(GND_net), .CIN(n11616), 
          .COUT(n11617), .S0(n5668[12]), .S1(n5668[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1096_14.INIT0 = 16'h5666;
    defparam add_1096_14.INIT1 = 16'h5666;
    defparam add_1096_14.INJECT1_0 = "NO";
    defparam add_1096_14.INJECT1_1 = "NO";
    CCU2D add_1096_12 (.A0(d4[46]), .B0(d5[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[47]), .B1(d5[47]), .C1(GND_net), .D1(GND_net), .CIN(n11615), 
          .COUT(n11616), .S0(n5668[10]), .S1(n5668[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1096_12.INIT0 = 16'h5666;
    defparam add_1096_12.INIT1 = 16'h5666;
    defparam add_1096_12.INJECT1_0 = "NO";
    defparam add_1096_12.INJECT1_1 = "NO";
    CCU2D add_1096_10 (.A0(d4[44]), .B0(d5[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[45]), .B1(d5[45]), .C1(GND_net), .D1(GND_net), .CIN(n11614), 
          .COUT(n11615), .S0(n5668[8]), .S1(n5668[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1096_10.INIT0 = 16'h5666;
    defparam add_1096_10.INIT1 = 16'h5666;
    defparam add_1096_10.INJECT1_0 = "NO";
    defparam add_1096_10.INJECT1_1 = "NO";
    CCU2D add_1096_8 (.A0(d4[42]), .B0(d5[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[43]), .B1(d5[43]), .C1(GND_net), .D1(GND_net), .CIN(n11613), 
          .COUT(n11614), .S0(n5668[6]), .S1(n5668[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1096_8.INIT0 = 16'h5666;
    defparam add_1096_8.INIT1 = 16'h5666;
    defparam add_1096_8.INJECT1_0 = "NO";
    defparam add_1096_8.INJECT1_1 = "NO";
    CCU2D add_1096_6 (.A0(d4[40]), .B0(d5[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[41]), .B1(d5[41]), .C1(GND_net), .D1(GND_net), .CIN(n11612), 
          .COUT(n11613), .S0(n5668[4]), .S1(n5668[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1096_6.INIT0 = 16'h5666;
    defparam add_1096_6.INIT1 = 16'h5666;
    defparam add_1096_6.INJECT1_0 = "NO";
    defparam add_1096_6.INJECT1_1 = "NO";
    CCU2D add_1096_4 (.A0(d4[38]), .B0(d5[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[39]), .B1(d5[39]), .C1(GND_net), .D1(GND_net), .CIN(n11611), 
          .COUT(n11612), .S0(n5668[2]), .S1(n5668[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1096_4.INIT0 = 16'h5666;
    defparam add_1096_4.INIT1 = 16'h5666;
    defparam add_1096_4.INJECT1_0 = "NO";
    defparam add_1096_4.INJECT1_1 = "NO";
    FD1P3AX d_tmp_i0_i1 (.D(d5[1]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i2 (.D(d5[2]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i3 (.D(d5[3]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i4 (.D(d5[4]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i5 (.D(d5[5]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i6 (.D(d5[6]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i7 (.D(d5[7]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i8 (.D(d5[8]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i9 (.D(d5[9]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i10 (.D(d5[10]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i11 (.D(d5[11]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i12 (.D(d5[12]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i13 (.D(d5[13]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i14 (.D(d5[14]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i15 (.D(d5[15]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i16 (.D(d5[16]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i17 (.D(d5[17]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i18 (.D(d5[18]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i19 (.D(d5[19]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i20 (.D(d5[20]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i21 (.D(d5[21]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i22 (.D(d5[22]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i23 (.D(d5[23]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i24 (.D(d5[24]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i25 (.D(d5[25]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i26 (.D(d5[26]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i27 (.D(d5[27]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i28 (.D(d5[28]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i29 (.D(d5[29]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i30 (.D(d5[30]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i31 (.D(d5[31]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i32 (.D(d5[32]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i33 (.D(d5[33]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i34 (.D(d5[34]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i35 (.D(d5[35]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i36 (.D(d5[36]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i37 (.D(d5[37]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i38 (.D(d5[38]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i39 (.D(d5[39]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i40 (.D(d5[40]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i41 (.D(d5[41]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i42 (.D(d5[42]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i43 (.D(d5[43]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i44 (.D(d5[44]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i45 (.D(d5[45]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i46 (.D(d5[46]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i47 (.D(d5[47]), .SP(osc_clk_enable_757), .CK(osc_clk), 
            .Q(d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i48 (.D(d5[48]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i49 (.D(d5[49]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i50 (.D(d5[50]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i51 (.D(d5[51]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i52 (.D(d5[52]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i53 (.D(d5[53]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i54 (.D(d5[54]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i55 (.D(d5[55]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i56 (.D(d5[56]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i57 (.D(d5[57]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i58 (.D(d5[58]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i59 (.D(d5[59]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i60 (.D(d5[60]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i61 (.D(d5[61]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i62 (.D(d5[62]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i63 (.D(d5[63]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i64 (.D(d5[64]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i65 (.D(d5[65]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i66 (.D(d5[66]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i67 (.D(d5[67]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i68 (.D(d5[68]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i69 (.D(d5[69]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i70 (.D(d5[70]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i71 (.D(d5[71]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i1 (.D(d_tmp[1]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i2 (.D(d_tmp[2]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i3 (.D(d_tmp[3]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i4 (.D(d_tmp[4]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i5 (.D(d_tmp[5]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i6 (.D(d_tmp[6]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i7 (.D(d_tmp[7]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i8 (.D(d_tmp[8]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i9 (.D(d_tmp[9]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i10 (.D(d_tmp[10]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i11 (.D(d_tmp[11]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i12 (.D(d_tmp[12]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i13 (.D(d_tmp[13]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i14 (.D(d_tmp[14]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i15 (.D(d_tmp[15]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i16 (.D(d_tmp[16]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i17 (.D(d_tmp[17]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i18 (.D(d_tmp[18]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i19 (.D(d_tmp[19]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i20 (.D(d_tmp[20]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i21 (.D(d_tmp[21]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i22 (.D(d_tmp[22]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i23 (.D(d_tmp[23]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i24 (.D(d_tmp[24]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i25 (.D(d_tmp[25]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i26 (.D(d_tmp[26]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i27 (.D(d_tmp[27]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i28 (.D(d_tmp[28]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i29 (.D(d_tmp[29]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i30 (.D(d_tmp[30]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i31 (.D(d_tmp[31]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i32 (.D(d_tmp[32]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i33 (.D(d_tmp[33]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i34 (.D(d_tmp[34]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i35 (.D(d_tmp[35]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i36 (.D(d_tmp[36]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i37 (.D(d_tmp[37]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i38 (.D(d_tmp[38]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i39 (.D(d_tmp[39]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i40 (.D(d_tmp[40]), .SP(osc_clk_enable_797), .CK(osc_clk), 
            .Q(d_d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i41 (.D(d_tmp[41]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i42 (.D(d_tmp[42]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i43 (.D(d_tmp[43]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i44 (.D(d_tmp[44]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i45 (.D(d_tmp[45]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i46 (.D(d_tmp[46]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i47 (.D(d_tmp[47]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i48 (.D(d_tmp[48]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i49 (.D(d_tmp[49]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i50 (.D(d_tmp[50]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i51 (.D(d_tmp[51]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i52 (.D(d_tmp[52]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i53 (.D(d_tmp[53]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i54 (.D(d_tmp[54]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i55 (.D(d_tmp[55]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i56 (.D(d_tmp[56]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i57 (.D(d_tmp[57]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i58 (.D(d_tmp[58]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i59 (.D(d_tmp[59]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i60 (.D(d_tmp[60]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i61 (.D(d_tmp[61]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i62 (.D(d_tmp[62]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i63 (.D(d_tmp[63]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i64 (.D(d_tmp[64]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i65 (.D(d_tmp[65]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i66 (.D(d_tmp[66]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i67 (.D(d_tmp[67]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i68 (.D(d_tmp[68]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i69 (.D(d_tmp[69]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i70 (.D(d_tmp[70]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i71 (.D(d_tmp[71]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d_d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i71.GSR = "ENABLED";
    FD1S3AX d2_i1 (.D(d2_71__N_490[1]), .CK(osc_clk), .Q(d2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i1.GSR = "ENABLED";
    FD1S3AX d2_i2 (.D(d2_71__N_490[2]), .CK(osc_clk), .Q(d2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i2.GSR = "ENABLED";
    FD1S3AX d2_i3 (.D(d2_71__N_490[3]), .CK(osc_clk), .Q(d2[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i3.GSR = "ENABLED";
    FD1S3AX d2_i4 (.D(d2_71__N_490[4]), .CK(osc_clk), .Q(d2[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i4.GSR = "ENABLED";
    FD1S3AX d2_i5 (.D(d2_71__N_490[5]), .CK(osc_clk), .Q(d2[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i5.GSR = "ENABLED";
    FD1S3AX d2_i6 (.D(d2_71__N_490[6]), .CK(osc_clk), .Q(d2[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i6.GSR = "ENABLED";
    FD1S3AX d2_i7 (.D(d2_71__N_490[7]), .CK(osc_clk), .Q(d2[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i7.GSR = "ENABLED";
    FD1S3AX d2_i8 (.D(d2_71__N_490[8]), .CK(osc_clk), .Q(d2[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i8.GSR = "ENABLED";
    FD1S3AX d2_i9 (.D(d2_71__N_490[9]), .CK(osc_clk), .Q(d2[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i9.GSR = "ENABLED";
    FD1S3AX d2_i10 (.D(d2_71__N_490[10]), .CK(osc_clk), .Q(d2[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i10.GSR = "ENABLED";
    FD1S3AX d2_i11 (.D(d2_71__N_490[11]), .CK(osc_clk), .Q(d2[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i11.GSR = "ENABLED";
    FD1S3AX d2_i12 (.D(d2_71__N_490[12]), .CK(osc_clk), .Q(d2[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i12.GSR = "ENABLED";
    FD1S3AX d2_i13 (.D(d2_71__N_490[13]), .CK(osc_clk), .Q(d2[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i13.GSR = "ENABLED";
    FD1S3AX d2_i14 (.D(d2_71__N_490[14]), .CK(osc_clk), .Q(d2[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i14.GSR = "ENABLED";
    FD1S3AX d2_i15 (.D(d2_71__N_490[15]), .CK(osc_clk), .Q(d2[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i15.GSR = "ENABLED";
    FD1S3AX d2_i16 (.D(d2_71__N_490[16]), .CK(osc_clk), .Q(d2[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i16.GSR = "ENABLED";
    FD1S3AX d2_i17 (.D(d2_71__N_490[17]), .CK(osc_clk), .Q(d2[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i17.GSR = "ENABLED";
    FD1S3AX d2_i18 (.D(d2_71__N_490[18]), .CK(osc_clk), .Q(d2[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i18.GSR = "ENABLED";
    FD1S3AX d2_i19 (.D(d2_71__N_490[19]), .CK(osc_clk), .Q(d2[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i19.GSR = "ENABLED";
    FD1S3AX d2_i20 (.D(d2_71__N_490[20]), .CK(osc_clk), .Q(d2[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i20.GSR = "ENABLED";
    FD1S3AX d2_i21 (.D(d2_71__N_490[21]), .CK(osc_clk), .Q(d2[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i21.GSR = "ENABLED";
    FD1S3AX d2_i22 (.D(d2_71__N_490[22]), .CK(osc_clk), .Q(d2[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i22.GSR = "ENABLED";
    FD1S3AX d2_i23 (.D(d2_71__N_490[23]), .CK(osc_clk), .Q(d2[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i23.GSR = "ENABLED";
    FD1S3AX d2_i24 (.D(d2_71__N_490[24]), .CK(osc_clk), .Q(d2[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i24.GSR = "ENABLED";
    FD1S3AX d2_i25 (.D(d2_71__N_490[25]), .CK(osc_clk), .Q(d2[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i25.GSR = "ENABLED";
    FD1S3AX d2_i26 (.D(d2_71__N_490[26]), .CK(osc_clk), .Q(d2[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i26.GSR = "ENABLED";
    FD1S3AX d2_i27 (.D(d2_71__N_490[27]), .CK(osc_clk), .Q(d2[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i27.GSR = "ENABLED";
    FD1S3AX d2_i28 (.D(d2_71__N_490[28]), .CK(osc_clk), .Q(d2[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i28.GSR = "ENABLED";
    FD1S3AX d2_i29 (.D(d2_71__N_490[29]), .CK(osc_clk), .Q(d2[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i29.GSR = "ENABLED";
    FD1S3AX d2_i30 (.D(d2_71__N_490[30]), .CK(osc_clk), .Q(d2[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i30.GSR = "ENABLED";
    FD1S3AX d2_i31 (.D(d2_71__N_490[31]), .CK(osc_clk), .Q(d2[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i31.GSR = "ENABLED";
    FD1S3AX d2_i32 (.D(d2_71__N_490[32]), .CK(osc_clk), .Q(d2[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i32.GSR = "ENABLED";
    FD1S3AX d2_i33 (.D(d2_71__N_490[33]), .CK(osc_clk), .Q(d2[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i33.GSR = "ENABLED";
    FD1S3AX d2_i34 (.D(d2_71__N_490[34]), .CK(osc_clk), .Q(d2[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i34.GSR = "ENABLED";
    FD1S3AX d2_i35 (.D(d2_71__N_490[35]), .CK(osc_clk), .Q(d2[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i35.GSR = "ENABLED";
    FD1S3AX d2_i36 (.D(d2_71__N_490[36]), .CK(osc_clk), .Q(d2[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i36.GSR = "ENABLED";
    FD1S3AX d2_i37 (.D(d2_71__N_490[37]), .CK(osc_clk), .Q(d2[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i37.GSR = "ENABLED";
    FD1S3AX d2_i38 (.D(d2_71__N_490[38]), .CK(osc_clk), .Q(d2[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i38.GSR = "ENABLED";
    FD1S3AX d2_i39 (.D(d2_71__N_490[39]), .CK(osc_clk), .Q(d2[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i39.GSR = "ENABLED";
    FD1S3AX d2_i40 (.D(d2_71__N_490[40]), .CK(osc_clk), .Q(d2[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i40.GSR = "ENABLED";
    FD1S3AX d2_i41 (.D(d2_71__N_490[41]), .CK(osc_clk), .Q(d2[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i41.GSR = "ENABLED";
    FD1S3AX d2_i42 (.D(d2_71__N_490[42]), .CK(osc_clk), .Q(d2[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i42.GSR = "ENABLED";
    FD1S3AX d2_i43 (.D(d2_71__N_490[43]), .CK(osc_clk), .Q(d2[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i43.GSR = "ENABLED";
    FD1S3AX d2_i44 (.D(d2_71__N_490[44]), .CK(osc_clk), .Q(d2[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i44.GSR = "ENABLED";
    FD1S3AX d2_i45 (.D(d2_71__N_490[45]), .CK(osc_clk), .Q(d2[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i45.GSR = "ENABLED";
    FD1S3AX d2_i46 (.D(d2_71__N_490[46]), .CK(osc_clk), .Q(d2[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i46.GSR = "ENABLED";
    FD1S3AX d2_i47 (.D(d2_71__N_490[47]), .CK(osc_clk), .Q(d2[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i47.GSR = "ENABLED";
    FD1S3AX d2_i48 (.D(d2_71__N_490[48]), .CK(osc_clk), .Q(d2[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i48.GSR = "ENABLED";
    FD1S3AX d2_i49 (.D(d2_71__N_490[49]), .CK(osc_clk), .Q(d2[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i49.GSR = "ENABLED";
    FD1S3AX d2_i50 (.D(d2_71__N_490[50]), .CK(osc_clk), .Q(d2[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i50.GSR = "ENABLED";
    FD1S3AX d2_i51 (.D(d2_71__N_490[51]), .CK(osc_clk), .Q(d2[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i51.GSR = "ENABLED";
    FD1S3AX d2_i52 (.D(d2_71__N_490[52]), .CK(osc_clk), .Q(d2[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i52.GSR = "ENABLED";
    FD1S3AX d2_i53 (.D(d2_71__N_490[53]), .CK(osc_clk), .Q(d2[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i53.GSR = "ENABLED";
    FD1S3AX d2_i54 (.D(d2_71__N_490[54]), .CK(osc_clk), .Q(d2[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i54.GSR = "ENABLED";
    FD1S3AX d2_i55 (.D(d2_71__N_490[55]), .CK(osc_clk), .Q(d2[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i55.GSR = "ENABLED";
    FD1S3AX d2_i56 (.D(d2_71__N_490[56]), .CK(osc_clk), .Q(d2[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i56.GSR = "ENABLED";
    FD1S3AX d2_i57 (.D(d2_71__N_490[57]), .CK(osc_clk), .Q(d2[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i57.GSR = "ENABLED";
    FD1S3AX d2_i58 (.D(d2_71__N_490[58]), .CK(osc_clk), .Q(d2[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i58.GSR = "ENABLED";
    FD1S3AX d2_i59 (.D(d2_71__N_490[59]), .CK(osc_clk), .Q(d2[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i59.GSR = "ENABLED";
    FD1S3AX d2_i60 (.D(d2_71__N_490[60]), .CK(osc_clk), .Q(d2[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i60.GSR = "ENABLED";
    FD1S3AX d2_i61 (.D(d2_71__N_490[61]), .CK(osc_clk), .Q(d2[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i61.GSR = "ENABLED";
    FD1S3AX d2_i62 (.D(d2_71__N_490[62]), .CK(osc_clk), .Q(d2[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i62.GSR = "ENABLED";
    FD1S3AX d2_i63 (.D(d2_71__N_490[63]), .CK(osc_clk), .Q(d2[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i63.GSR = "ENABLED";
    FD1S3AX d2_i64 (.D(d2_71__N_490[64]), .CK(osc_clk), .Q(d2[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i64.GSR = "ENABLED";
    FD1S3AX d2_i65 (.D(d2_71__N_490[65]), .CK(osc_clk), .Q(d2[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i65.GSR = "ENABLED";
    FD1S3AX d2_i66 (.D(d2_71__N_490[66]), .CK(osc_clk), .Q(d2[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i66.GSR = "ENABLED";
    FD1S3AX d2_i67 (.D(d2_71__N_490[67]), .CK(osc_clk), .Q(d2[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i67.GSR = "ENABLED";
    FD1S3AX d2_i68 (.D(d2_71__N_490[68]), .CK(osc_clk), .Q(d2[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i68.GSR = "ENABLED";
    FD1S3AX d2_i69 (.D(d2_71__N_490[69]), .CK(osc_clk), .Q(d2[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i69.GSR = "ENABLED";
    FD1S3AX d2_i70 (.D(d2_71__N_490[70]), .CK(osc_clk), .Q(d2[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i70.GSR = "ENABLED";
    FD1S3AX d2_i71 (.D(d2_71__N_490[71]), .CK(osc_clk), .Q(d2[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i71.GSR = "ENABLED";
    FD1S3AX d3_i1 (.D(d3_71__N_562[1]), .CK(osc_clk), .Q(d3[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i1.GSR = "ENABLED";
    FD1S3AX d3_i2 (.D(d3_71__N_562[2]), .CK(osc_clk), .Q(d3[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i2.GSR = "ENABLED";
    FD1S3AX d3_i3 (.D(d3_71__N_562[3]), .CK(osc_clk), .Q(d3[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i3.GSR = "ENABLED";
    FD1S3AX d3_i4 (.D(d3_71__N_562[4]), .CK(osc_clk), .Q(d3[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i4.GSR = "ENABLED";
    FD1S3AX d3_i5 (.D(d3_71__N_562[5]), .CK(osc_clk), .Q(d3[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i5.GSR = "ENABLED";
    FD1S3AX d3_i6 (.D(d3_71__N_562[6]), .CK(osc_clk), .Q(d3[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i6.GSR = "ENABLED";
    FD1S3AX d3_i7 (.D(d3_71__N_562[7]), .CK(osc_clk), .Q(d3[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i7.GSR = "ENABLED";
    FD1S3AX d3_i8 (.D(d3_71__N_562[8]), .CK(osc_clk), .Q(d3[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i8.GSR = "ENABLED";
    FD1S3AX d3_i9 (.D(d3_71__N_562[9]), .CK(osc_clk), .Q(d3[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i9.GSR = "ENABLED";
    FD1S3AX d3_i10 (.D(d3_71__N_562[10]), .CK(osc_clk), .Q(d3[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i10.GSR = "ENABLED";
    FD1S3AX d3_i11 (.D(d3_71__N_562[11]), .CK(osc_clk), .Q(d3[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i11.GSR = "ENABLED";
    FD1S3AX d3_i12 (.D(d3_71__N_562[12]), .CK(osc_clk), .Q(d3[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i12.GSR = "ENABLED";
    FD1S3AX d3_i13 (.D(d3_71__N_562[13]), .CK(osc_clk), .Q(d3[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i13.GSR = "ENABLED";
    FD1S3AX d3_i14 (.D(d3_71__N_562[14]), .CK(osc_clk), .Q(d3[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i14.GSR = "ENABLED";
    FD1S3AX d3_i15 (.D(d3_71__N_562[15]), .CK(osc_clk), .Q(d3[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i15.GSR = "ENABLED";
    FD1S3AX d3_i16 (.D(d3_71__N_562[16]), .CK(osc_clk), .Q(d3[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i16.GSR = "ENABLED";
    FD1S3AX d3_i17 (.D(d3_71__N_562[17]), .CK(osc_clk), .Q(d3[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i17.GSR = "ENABLED";
    FD1S3AX d3_i18 (.D(d3_71__N_562[18]), .CK(osc_clk), .Q(d3[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i18.GSR = "ENABLED";
    FD1S3AX d3_i19 (.D(d3_71__N_562[19]), .CK(osc_clk), .Q(d3[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i19.GSR = "ENABLED";
    FD1S3AX d3_i20 (.D(d3_71__N_562[20]), .CK(osc_clk), .Q(d3[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i20.GSR = "ENABLED";
    FD1S3AX d3_i21 (.D(d3_71__N_562[21]), .CK(osc_clk), .Q(d3[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i21.GSR = "ENABLED";
    FD1S3AX d3_i22 (.D(d3_71__N_562[22]), .CK(osc_clk), .Q(d3[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i22.GSR = "ENABLED";
    FD1S3AX d3_i23 (.D(d3_71__N_562[23]), .CK(osc_clk), .Q(d3[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i23.GSR = "ENABLED";
    FD1S3AX d3_i24 (.D(d3_71__N_562[24]), .CK(osc_clk), .Q(d3[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i24.GSR = "ENABLED";
    FD1S3AX d3_i25 (.D(d3_71__N_562[25]), .CK(osc_clk), .Q(d3[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i25.GSR = "ENABLED";
    FD1S3AX d3_i26 (.D(d3_71__N_562[26]), .CK(osc_clk), .Q(d3[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i26.GSR = "ENABLED";
    FD1S3AX d3_i27 (.D(d3_71__N_562[27]), .CK(osc_clk), .Q(d3[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i27.GSR = "ENABLED";
    FD1S3AX d3_i28 (.D(d3_71__N_562[28]), .CK(osc_clk), .Q(d3[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i28.GSR = "ENABLED";
    FD1S3AX d3_i29 (.D(d3_71__N_562[29]), .CK(osc_clk), .Q(d3[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i29.GSR = "ENABLED";
    FD1S3AX d3_i30 (.D(d3_71__N_562[30]), .CK(osc_clk), .Q(d3[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i30.GSR = "ENABLED";
    FD1S3AX d3_i31 (.D(d3_71__N_562[31]), .CK(osc_clk), .Q(d3[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i31.GSR = "ENABLED";
    FD1S3AX d3_i32 (.D(d3_71__N_562[32]), .CK(osc_clk), .Q(d3[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i32.GSR = "ENABLED";
    FD1S3AX d3_i33 (.D(d3_71__N_562[33]), .CK(osc_clk), .Q(d3[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i33.GSR = "ENABLED";
    FD1S3AX d3_i34 (.D(d3_71__N_562[34]), .CK(osc_clk), .Q(d3[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i34.GSR = "ENABLED";
    FD1S3AX d3_i35 (.D(d3_71__N_562[35]), .CK(osc_clk), .Q(d3[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i35.GSR = "ENABLED";
    FD1S3AX d3_i36 (.D(d3_71__N_562[36]), .CK(osc_clk), .Q(d3[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i36.GSR = "ENABLED";
    FD1S3AX d3_i37 (.D(d3_71__N_562[37]), .CK(osc_clk), .Q(d3[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i37.GSR = "ENABLED";
    FD1S3AX d3_i38 (.D(d3_71__N_562[38]), .CK(osc_clk), .Q(d3[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i38.GSR = "ENABLED";
    FD1S3AX d3_i39 (.D(d3_71__N_562[39]), .CK(osc_clk), .Q(d3[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i39.GSR = "ENABLED";
    FD1S3AX d3_i40 (.D(d3_71__N_562[40]), .CK(osc_clk), .Q(d3[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i40.GSR = "ENABLED";
    FD1S3AX d3_i41 (.D(d3_71__N_562[41]), .CK(osc_clk), .Q(d3[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i41.GSR = "ENABLED";
    FD1S3AX d3_i42 (.D(d3_71__N_562[42]), .CK(osc_clk), .Q(d3[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i42.GSR = "ENABLED";
    FD1S3AX d3_i43 (.D(d3_71__N_562[43]), .CK(osc_clk), .Q(d3[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i43.GSR = "ENABLED";
    FD1S3AX d3_i44 (.D(d3_71__N_562[44]), .CK(osc_clk), .Q(d3[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i44.GSR = "ENABLED";
    FD1S3AX d3_i45 (.D(d3_71__N_562[45]), .CK(osc_clk), .Q(d3[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i45.GSR = "ENABLED";
    FD1S3AX d3_i46 (.D(d3_71__N_562[46]), .CK(osc_clk), .Q(d3[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i46.GSR = "ENABLED";
    FD1S3AX d3_i47 (.D(d3_71__N_562[47]), .CK(osc_clk), .Q(d3[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i47.GSR = "ENABLED";
    FD1S3AX d3_i48 (.D(d3_71__N_562[48]), .CK(osc_clk), .Q(d3[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i48.GSR = "ENABLED";
    FD1S3AX d3_i49 (.D(d3_71__N_562[49]), .CK(osc_clk), .Q(d3[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i49.GSR = "ENABLED";
    FD1S3AX d3_i50 (.D(d3_71__N_562[50]), .CK(osc_clk), .Q(d3[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i50.GSR = "ENABLED";
    FD1S3AX d3_i51 (.D(d3_71__N_562[51]), .CK(osc_clk), .Q(d3[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i51.GSR = "ENABLED";
    FD1S3AX d3_i52 (.D(d3_71__N_562[52]), .CK(osc_clk), .Q(d3[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i52.GSR = "ENABLED";
    FD1S3AX d3_i53 (.D(d3_71__N_562[53]), .CK(osc_clk), .Q(d3[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i53.GSR = "ENABLED";
    FD1S3AX d3_i54 (.D(d3_71__N_562[54]), .CK(osc_clk), .Q(d3[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i54.GSR = "ENABLED";
    FD1S3AX d3_i55 (.D(d3_71__N_562[55]), .CK(osc_clk), .Q(d3[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i55.GSR = "ENABLED";
    FD1S3AX d3_i56 (.D(d3_71__N_562[56]), .CK(osc_clk), .Q(d3[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i56.GSR = "ENABLED";
    FD1S3AX d3_i57 (.D(d3_71__N_562[57]), .CK(osc_clk), .Q(d3[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i57.GSR = "ENABLED";
    FD1S3AX d3_i58 (.D(d3_71__N_562[58]), .CK(osc_clk), .Q(d3[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i58.GSR = "ENABLED";
    FD1S3AX d3_i59 (.D(d3_71__N_562[59]), .CK(osc_clk), .Q(d3[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i59.GSR = "ENABLED";
    FD1S3AX d3_i60 (.D(d3_71__N_562[60]), .CK(osc_clk), .Q(d3[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i60.GSR = "ENABLED";
    FD1S3AX d3_i61 (.D(d3_71__N_562[61]), .CK(osc_clk), .Q(d3[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i61.GSR = "ENABLED";
    FD1S3AX d3_i62 (.D(d3_71__N_562[62]), .CK(osc_clk), .Q(d3[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i62.GSR = "ENABLED";
    FD1S3AX d3_i63 (.D(d3_71__N_562[63]), .CK(osc_clk), .Q(d3[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i63.GSR = "ENABLED";
    FD1S3AX d3_i64 (.D(d3_71__N_562[64]), .CK(osc_clk), .Q(d3[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i64.GSR = "ENABLED";
    FD1S3AX d3_i65 (.D(d3_71__N_562[65]), .CK(osc_clk), .Q(d3[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i65.GSR = "ENABLED";
    FD1S3AX d3_i66 (.D(d3_71__N_562[66]), .CK(osc_clk), .Q(d3[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i66.GSR = "ENABLED";
    FD1S3AX d3_i67 (.D(d3_71__N_562[67]), .CK(osc_clk), .Q(d3[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i67.GSR = "ENABLED";
    FD1S3AX d3_i68 (.D(d3_71__N_562[68]), .CK(osc_clk), .Q(d3[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i68.GSR = "ENABLED";
    FD1S3AX d3_i69 (.D(d3_71__N_562[69]), .CK(osc_clk), .Q(d3[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i69.GSR = "ENABLED";
    FD1S3AX d3_i70 (.D(d3_71__N_562[70]), .CK(osc_clk), .Q(d3[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i70.GSR = "ENABLED";
    FD1S3AX d3_i71 (.D(d3_71__N_562[71]), .CK(osc_clk), .Q(d3[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i71.GSR = "ENABLED";
    FD1S3AX d4_i1 (.D(d4_71__N_634[1]), .CK(osc_clk), .Q(d4[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i1.GSR = "ENABLED";
    FD1S3AX d4_i2 (.D(d4_71__N_634[2]), .CK(osc_clk), .Q(d4[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i2.GSR = "ENABLED";
    FD1S3AX d4_i3 (.D(d4_71__N_634[3]), .CK(osc_clk), .Q(d4[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i3.GSR = "ENABLED";
    FD1S3AX d4_i4 (.D(d4_71__N_634[4]), .CK(osc_clk), .Q(d4[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i4.GSR = "ENABLED";
    FD1S3AX d4_i5 (.D(d4_71__N_634[5]), .CK(osc_clk), .Q(d4[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i5.GSR = "ENABLED";
    FD1S3AX d4_i6 (.D(d4_71__N_634[6]), .CK(osc_clk), .Q(d4[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i6.GSR = "ENABLED";
    FD1S3AX d4_i7 (.D(d4_71__N_634[7]), .CK(osc_clk), .Q(d4[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i7.GSR = "ENABLED";
    FD1S3AX d4_i8 (.D(d4_71__N_634[8]), .CK(osc_clk), .Q(d4[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i8.GSR = "ENABLED";
    FD1S3AX d4_i9 (.D(d4_71__N_634[9]), .CK(osc_clk), .Q(d4[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i9.GSR = "ENABLED";
    FD1S3AX d4_i10 (.D(d4_71__N_634[10]), .CK(osc_clk), .Q(d4[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i10.GSR = "ENABLED";
    FD1S3AX d4_i11 (.D(d4_71__N_634[11]), .CK(osc_clk), .Q(d4[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i11.GSR = "ENABLED";
    FD1S3AX d4_i12 (.D(d4_71__N_634[12]), .CK(osc_clk), .Q(d4[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i12.GSR = "ENABLED";
    FD1S3AX d4_i13 (.D(d4_71__N_634[13]), .CK(osc_clk), .Q(d4[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i13.GSR = "ENABLED";
    FD1S3AX d4_i14 (.D(d4_71__N_634[14]), .CK(osc_clk), .Q(d4[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i14.GSR = "ENABLED";
    FD1S3AX d4_i15 (.D(d4_71__N_634[15]), .CK(osc_clk), .Q(d4[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i15.GSR = "ENABLED";
    FD1S3AX d4_i16 (.D(d4_71__N_634[16]), .CK(osc_clk), .Q(d4[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i16.GSR = "ENABLED";
    FD1S3AX d4_i17 (.D(d4_71__N_634[17]), .CK(osc_clk), .Q(d4[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i17.GSR = "ENABLED";
    FD1S3AX d4_i18 (.D(d4_71__N_634[18]), .CK(osc_clk), .Q(d4[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i18.GSR = "ENABLED";
    FD1S3AX d4_i19 (.D(d4_71__N_634[19]), .CK(osc_clk), .Q(d4[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i19.GSR = "ENABLED";
    FD1S3AX d4_i20 (.D(d4_71__N_634[20]), .CK(osc_clk), .Q(d4[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i20.GSR = "ENABLED";
    FD1S3AX d4_i21 (.D(d4_71__N_634[21]), .CK(osc_clk), .Q(d4[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i21.GSR = "ENABLED";
    FD1S3AX d4_i22 (.D(d4_71__N_634[22]), .CK(osc_clk), .Q(d4[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i22.GSR = "ENABLED";
    FD1S3AX d4_i23 (.D(d4_71__N_634[23]), .CK(osc_clk), .Q(d4[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i23.GSR = "ENABLED";
    FD1S3AX d4_i24 (.D(d4_71__N_634[24]), .CK(osc_clk), .Q(d4[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i24.GSR = "ENABLED";
    FD1S3AX d4_i25 (.D(d4_71__N_634[25]), .CK(osc_clk), .Q(d4[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i25.GSR = "ENABLED";
    FD1S3AX d4_i26 (.D(d4_71__N_634[26]), .CK(osc_clk), .Q(d4[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i26.GSR = "ENABLED";
    FD1S3AX d4_i27 (.D(d4_71__N_634[27]), .CK(osc_clk), .Q(d4[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i27.GSR = "ENABLED";
    FD1S3AX d4_i28 (.D(d4_71__N_634[28]), .CK(osc_clk), .Q(d4[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i28.GSR = "ENABLED";
    FD1S3AX d4_i29 (.D(d4_71__N_634[29]), .CK(osc_clk), .Q(d4[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i29.GSR = "ENABLED";
    FD1S3AX d4_i30 (.D(d4_71__N_634[30]), .CK(osc_clk), .Q(d4[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i30.GSR = "ENABLED";
    FD1S3AX d4_i31 (.D(d4_71__N_634[31]), .CK(osc_clk), .Q(d4[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i31.GSR = "ENABLED";
    FD1S3AX d4_i32 (.D(d4_71__N_634[32]), .CK(osc_clk), .Q(d4[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i32.GSR = "ENABLED";
    FD1S3AX d4_i33 (.D(d4_71__N_634[33]), .CK(osc_clk), .Q(d4[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i33.GSR = "ENABLED";
    FD1S3AX d4_i34 (.D(d4_71__N_634[34]), .CK(osc_clk), .Q(d4[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i34.GSR = "ENABLED";
    FD1S3AX d4_i35 (.D(d4_71__N_634[35]), .CK(osc_clk), .Q(d4[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i35.GSR = "ENABLED";
    FD1S3AX d4_i36 (.D(d4_71__N_634[36]), .CK(osc_clk), .Q(d4[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i36.GSR = "ENABLED";
    FD1S3AX d4_i37 (.D(d4_71__N_634[37]), .CK(osc_clk), .Q(d4[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i37.GSR = "ENABLED";
    FD1S3AX d4_i38 (.D(d4_71__N_634[38]), .CK(osc_clk), .Q(d4[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i38.GSR = "ENABLED";
    FD1S3AX d4_i39 (.D(d4_71__N_634[39]), .CK(osc_clk), .Q(d4[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i39.GSR = "ENABLED";
    FD1S3AX d4_i40 (.D(d4_71__N_634[40]), .CK(osc_clk), .Q(d4[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i40.GSR = "ENABLED";
    FD1S3AX d4_i41 (.D(d4_71__N_634[41]), .CK(osc_clk), .Q(d4[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i41.GSR = "ENABLED";
    FD1S3AX d4_i42 (.D(d4_71__N_634[42]), .CK(osc_clk), .Q(d4[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i42.GSR = "ENABLED";
    FD1S3AX d4_i43 (.D(d4_71__N_634[43]), .CK(osc_clk), .Q(d4[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i43.GSR = "ENABLED";
    FD1S3AX d4_i44 (.D(d4_71__N_634[44]), .CK(osc_clk), .Q(d4[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i44.GSR = "ENABLED";
    FD1S3AX d4_i45 (.D(d4_71__N_634[45]), .CK(osc_clk), .Q(d4[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i45.GSR = "ENABLED";
    FD1S3AX d4_i46 (.D(d4_71__N_634[46]), .CK(osc_clk), .Q(d4[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i46.GSR = "ENABLED";
    FD1S3AX d4_i47 (.D(d4_71__N_634[47]), .CK(osc_clk), .Q(d4[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i47.GSR = "ENABLED";
    FD1S3AX d4_i48 (.D(d4_71__N_634[48]), .CK(osc_clk), .Q(d4[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i48.GSR = "ENABLED";
    FD1S3AX d4_i49 (.D(d4_71__N_634[49]), .CK(osc_clk), .Q(d4[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i49.GSR = "ENABLED";
    FD1S3AX d4_i50 (.D(d4_71__N_634[50]), .CK(osc_clk), .Q(d4[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i50.GSR = "ENABLED";
    FD1S3AX d4_i51 (.D(d4_71__N_634[51]), .CK(osc_clk), .Q(d4[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i51.GSR = "ENABLED";
    FD1S3AX d4_i52 (.D(d4_71__N_634[52]), .CK(osc_clk), .Q(d4[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i52.GSR = "ENABLED";
    FD1S3AX d4_i53 (.D(d4_71__N_634[53]), .CK(osc_clk), .Q(d4[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i53.GSR = "ENABLED";
    FD1S3AX d4_i54 (.D(d4_71__N_634[54]), .CK(osc_clk), .Q(d4[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i54.GSR = "ENABLED";
    FD1S3AX d4_i55 (.D(d4_71__N_634[55]), .CK(osc_clk), .Q(d4[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i55.GSR = "ENABLED";
    FD1S3AX d4_i56 (.D(d4_71__N_634[56]), .CK(osc_clk), .Q(d4[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i56.GSR = "ENABLED";
    FD1S3AX d4_i57 (.D(d4_71__N_634[57]), .CK(osc_clk), .Q(d4[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i57.GSR = "ENABLED";
    FD1S3AX d4_i58 (.D(d4_71__N_634[58]), .CK(osc_clk), .Q(d4[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i58.GSR = "ENABLED";
    FD1S3AX d4_i59 (.D(d4_71__N_634[59]), .CK(osc_clk), .Q(d4[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i59.GSR = "ENABLED";
    FD1S3AX d4_i60 (.D(d4_71__N_634[60]), .CK(osc_clk), .Q(d4[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i60.GSR = "ENABLED";
    FD1S3AX d4_i61 (.D(d4_71__N_634[61]), .CK(osc_clk), .Q(d4[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i61.GSR = "ENABLED";
    FD1S3AX d4_i62 (.D(d4_71__N_634[62]), .CK(osc_clk), .Q(d4[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i62.GSR = "ENABLED";
    FD1S3AX d4_i63 (.D(d4_71__N_634[63]), .CK(osc_clk), .Q(d4[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i63.GSR = "ENABLED";
    FD1S3AX d4_i64 (.D(d4_71__N_634[64]), .CK(osc_clk), .Q(d4[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i64.GSR = "ENABLED";
    FD1S3AX d4_i65 (.D(d4_71__N_634[65]), .CK(osc_clk), .Q(d4[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i65.GSR = "ENABLED";
    FD1S3AX d4_i66 (.D(d4_71__N_634[66]), .CK(osc_clk), .Q(d4[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i66.GSR = "ENABLED";
    FD1S3AX d4_i67 (.D(d4_71__N_634[67]), .CK(osc_clk), .Q(d4[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i67.GSR = "ENABLED";
    FD1S3AX d4_i68 (.D(d4_71__N_634[68]), .CK(osc_clk), .Q(d4[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i68.GSR = "ENABLED";
    FD1S3AX d4_i69 (.D(d4_71__N_634[69]), .CK(osc_clk), .Q(d4[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i69.GSR = "ENABLED";
    FD1S3AX d4_i70 (.D(d4_71__N_634[70]), .CK(osc_clk), .Q(d4[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i70.GSR = "ENABLED";
    FD1S3AX d4_i71 (.D(d4_71__N_634[71]), .CK(osc_clk), .Q(d4[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i71.GSR = "ENABLED";
    FD1S3AX d5_i1 (.D(d5_71__N_706[1]), .CK(osc_clk), .Q(d5[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i1.GSR = "ENABLED";
    FD1S3AX d5_i2 (.D(d5_71__N_706[2]), .CK(osc_clk), .Q(d5[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i2.GSR = "ENABLED";
    FD1S3AX d5_i3 (.D(d5_71__N_706[3]), .CK(osc_clk), .Q(d5[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i3.GSR = "ENABLED";
    FD1S3AX d5_i4 (.D(d5_71__N_706[4]), .CK(osc_clk), .Q(d5[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i4.GSR = "ENABLED";
    FD1S3AX d5_i5 (.D(d5_71__N_706[5]), .CK(osc_clk), .Q(d5[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i5.GSR = "ENABLED";
    FD1S3AX d5_i6 (.D(d5_71__N_706[6]), .CK(osc_clk), .Q(d5[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i6.GSR = "ENABLED";
    FD1S3AX d5_i7 (.D(d5_71__N_706[7]), .CK(osc_clk), .Q(d5[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i7.GSR = "ENABLED";
    FD1S3AX d5_i8 (.D(d5_71__N_706[8]), .CK(osc_clk), .Q(d5[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i8.GSR = "ENABLED";
    FD1S3AX d5_i9 (.D(d5_71__N_706[9]), .CK(osc_clk), .Q(d5[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i9.GSR = "ENABLED";
    FD1S3AX d5_i10 (.D(d5_71__N_706[10]), .CK(osc_clk), .Q(d5[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i10.GSR = "ENABLED";
    FD1S3AX d5_i11 (.D(d5_71__N_706[11]), .CK(osc_clk), .Q(d5[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i11.GSR = "ENABLED";
    FD1S3AX d5_i12 (.D(d5_71__N_706[12]), .CK(osc_clk), .Q(d5[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i12.GSR = "ENABLED";
    FD1S3AX d5_i13 (.D(d5_71__N_706[13]), .CK(osc_clk), .Q(d5[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i13.GSR = "ENABLED";
    FD1S3AX d5_i14 (.D(d5_71__N_706[14]), .CK(osc_clk), .Q(d5[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i14.GSR = "ENABLED";
    FD1S3AX d5_i15 (.D(d5_71__N_706[15]), .CK(osc_clk), .Q(d5[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i15.GSR = "ENABLED";
    FD1S3AX d5_i16 (.D(d5_71__N_706[16]), .CK(osc_clk), .Q(d5[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i16.GSR = "ENABLED";
    FD1S3AX d5_i17 (.D(d5_71__N_706[17]), .CK(osc_clk), .Q(d5[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i17.GSR = "ENABLED";
    FD1S3AX d5_i18 (.D(d5_71__N_706[18]), .CK(osc_clk), .Q(d5[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i18.GSR = "ENABLED";
    FD1S3AX d5_i19 (.D(d5_71__N_706[19]), .CK(osc_clk), .Q(d5[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i19.GSR = "ENABLED";
    FD1S3AX d5_i20 (.D(d5_71__N_706[20]), .CK(osc_clk), .Q(d5[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i20.GSR = "ENABLED";
    FD1S3AX d5_i21 (.D(d5_71__N_706[21]), .CK(osc_clk), .Q(d5[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i21.GSR = "ENABLED";
    FD1S3AX d5_i22 (.D(d5_71__N_706[22]), .CK(osc_clk), .Q(d5[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i22.GSR = "ENABLED";
    FD1S3AX d5_i23 (.D(d5_71__N_706[23]), .CK(osc_clk), .Q(d5[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i23.GSR = "ENABLED";
    FD1S3AX d5_i24 (.D(d5_71__N_706[24]), .CK(osc_clk), .Q(d5[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i24.GSR = "ENABLED";
    FD1S3AX d5_i25 (.D(d5_71__N_706[25]), .CK(osc_clk), .Q(d5[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i25.GSR = "ENABLED";
    FD1S3AX d5_i26 (.D(d5_71__N_706[26]), .CK(osc_clk), .Q(d5[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i26.GSR = "ENABLED";
    FD1S3AX d5_i27 (.D(d5_71__N_706[27]), .CK(osc_clk), .Q(d5[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i27.GSR = "ENABLED";
    FD1S3AX d5_i28 (.D(d5_71__N_706[28]), .CK(osc_clk), .Q(d5[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i28.GSR = "ENABLED";
    FD1S3AX d5_i29 (.D(d5_71__N_706[29]), .CK(osc_clk), .Q(d5[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i29.GSR = "ENABLED";
    FD1S3AX d5_i30 (.D(d5_71__N_706[30]), .CK(osc_clk), .Q(d5[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i30.GSR = "ENABLED";
    FD1S3AX d5_i31 (.D(d5_71__N_706[31]), .CK(osc_clk), .Q(d5[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i31.GSR = "ENABLED";
    FD1S3AX d5_i32 (.D(d5_71__N_706[32]), .CK(osc_clk), .Q(d5[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i32.GSR = "ENABLED";
    FD1S3AX d5_i33 (.D(d5_71__N_706[33]), .CK(osc_clk), .Q(d5[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i33.GSR = "ENABLED";
    FD1S3AX d5_i34 (.D(d5_71__N_706[34]), .CK(osc_clk), .Q(d5[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i34.GSR = "ENABLED";
    FD1S3AX d5_i35 (.D(d5_71__N_706[35]), .CK(osc_clk), .Q(d5[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i35.GSR = "ENABLED";
    FD1S3AX d5_i36 (.D(d5_71__N_706[36]), .CK(osc_clk), .Q(d5[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i36.GSR = "ENABLED";
    FD1S3AX d5_i37 (.D(d5_71__N_706[37]), .CK(osc_clk), .Q(d5[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i37.GSR = "ENABLED";
    FD1S3AX d5_i38 (.D(d5_71__N_706[38]), .CK(osc_clk), .Q(d5[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i38.GSR = "ENABLED";
    FD1S3AX d5_i39 (.D(d5_71__N_706[39]), .CK(osc_clk), .Q(d5[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i39.GSR = "ENABLED";
    FD1S3AX d5_i40 (.D(d5_71__N_706[40]), .CK(osc_clk), .Q(d5[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i40.GSR = "ENABLED";
    FD1S3AX d5_i41 (.D(d5_71__N_706[41]), .CK(osc_clk), .Q(d5[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i41.GSR = "ENABLED";
    FD1S3AX d5_i42 (.D(d5_71__N_706[42]), .CK(osc_clk), .Q(d5[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i42.GSR = "ENABLED";
    FD1S3AX d5_i43 (.D(d5_71__N_706[43]), .CK(osc_clk), .Q(d5[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i43.GSR = "ENABLED";
    FD1S3AX d5_i44 (.D(d5_71__N_706[44]), .CK(osc_clk), .Q(d5[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i44.GSR = "ENABLED";
    FD1S3AX d5_i45 (.D(d5_71__N_706[45]), .CK(osc_clk), .Q(d5[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i45.GSR = "ENABLED";
    FD1S3AX d5_i46 (.D(d5_71__N_706[46]), .CK(osc_clk), .Q(d5[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i46.GSR = "ENABLED";
    FD1S3AX d5_i47 (.D(d5_71__N_706[47]), .CK(osc_clk), .Q(d5[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i47.GSR = "ENABLED";
    FD1S3AX d5_i48 (.D(d5_71__N_706[48]), .CK(osc_clk), .Q(d5[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i48.GSR = "ENABLED";
    FD1S3AX d5_i49 (.D(d5_71__N_706[49]), .CK(osc_clk), .Q(d5[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i49.GSR = "ENABLED";
    FD1S3AX d5_i50 (.D(d5_71__N_706[50]), .CK(osc_clk), .Q(d5[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i50.GSR = "ENABLED";
    FD1S3AX d5_i51 (.D(d5_71__N_706[51]), .CK(osc_clk), .Q(d5[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i51.GSR = "ENABLED";
    FD1S3AX d5_i52 (.D(d5_71__N_706[52]), .CK(osc_clk), .Q(d5[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i52.GSR = "ENABLED";
    FD1S3AX d5_i53 (.D(d5_71__N_706[53]), .CK(osc_clk), .Q(d5[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i53.GSR = "ENABLED";
    FD1S3AX d5_i54 (.D(d5_71__N_706[54]), .CK(osc_clk), .Q(d5[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i54.GSR = "ENABLED";
    FD1S3AX d5_i55 (.D(d5_71__N_706[55]), .CK(osc_clk), .Q(d5[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i55.GSR = "ENABLED";
    FD1S3AX d5_i56 (.D(d5_71__N_706[56]), .CK(osc_clk), .Q(d5[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i56.GSR = "ENABLED";
    FD1S3AX d5_i57 (.D(d5_71__N_706[57]), .CK(osc_clk), .Q(d5[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i57.GSR = "ENABLED";
    FD1S3AX d5_i58 (.D(d5_71__N_706[58]), .CK(osc_clk), .Q(d5[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i58.GSR = "ENABLED";
    FD1S3AX d5_i59 (.D(d5_71__N_706[59]), .CK(osc_clk), .Q(d5[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i59.GSR = "ENABLED";
    FD1S3AX d5_i60 (.D(d5_71__N_706[60]), .CK(osc_clk), .Q(d5[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i60.GSR = "ENABLED";
    FD1S3AX d5_i61 (.D(d5_71__N_706[61]), .CK(osc_clk), .Q(d5[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i61.GSR = "ENABLED";
    FD1S3AX d5_i62 (.D(d5_71__N_706[62]), .CK(osc_clk), .Q(d5[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i62.GSR = "ENABLED";
    FD1S3AX d5_i63 (.D(d5_71__N_706[63]), .CK(osc_clk), .Q(d5[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i63.GSR = "ENABLED";
    FD1S3AX d5_i64 (.D(d5_71__N_706[64]), .CK(osc_clk), .Q(d5[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i64.GSR = "ENABLED";
    FD1S3AX d5_i65 (.D(d5_71__N_706[65]), .CK(osc_clk), .Q(d5[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i65.GSR = "ENABLED";
    FD1S3AX d5_i66 (.D(d5_71__N_706[66]), .CK(osc_clk), .Q(d5[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i66.GSR = "ENABLED";
    FD1S3AX d5_i67 (.D(d5_71__N_706[67]), .CK(osc_clk), .Q(d5[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i67.GSR = "ENABLED";
    FD1S3AX d5_i68 (.D(d5_71__N_706[68]), .CK(osc_clk), .Q(d5[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i68.GSR = "ENABLED";
    FD1S3AX d5_i69 (.D(d5_71__N_706[69]), .CK(osc_clk), .Q(d5[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i69.GSR = "ENABLED";
    FD1S3AX d5_i70 (.D(d5_71__N_706[70]), .CK(osc_clk), .Q(d5[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i70.GSR = "ENABLED";
    FD1S3AX d5_i71 (.D(d5_71__N_706[71]), .CK(osc_clk), .Q(d5[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i71.GSR = "ENABLED";
    FD1P3AX d6_i0_i1 (.D(d6_71__N_1459[1]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d6_i0_i2 (.D(d6_71__N_1459[2]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d6_i0_i3 (.D(d6_71__N_1459[3]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d6_i0_i4 (.D(d6_71__N_1459[4]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d6_i0_i5 (.D(d6_71__N_1459[5]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d6_i0_i6 (.D(d6_71__N_1459[6]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d6_i0_i7 (.D(d6_71__N_1459[7]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d6_i0_i8 (.D(d6_71__N_1459[8]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d6_i0_i9 (.D(d6_71__N_1459[9]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d6_i0_i10 (.D(d6_71__N_1459[10]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d6_i0_i11 (.D(d6_71__N_1459[11]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d6_i0_i12 (.D(d6_71__N_1459[12]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d6_i0_i13 (.D(d6_71__N_1459[13]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d6_i0_i14 (.D(d6_71__N_1459[14]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d6_i0_i15 (.D(d6_71__N_1459[15]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d6_i0_i16 (.D(d6_71__N_1459[16]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d6_i0_i17 (.D(d6_71__N_1459[17]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d6_i0_i18 (.D(d6_71__N_1459[18]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d6_i0_i19 (.D(d6_71__N_1459[19]), .SP(osc_clk_enable_847), .CK(osc_clk), 
            .Q(d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d6_i0_i20 (.D(d6_71__N_1459[20]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d6_i0_i21 (.D(d6_71__N_1459[21]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d6_i0_i22 (.D(d6_71__N_1459[22]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d6_i0_i23 (.D(d6_71__N_1459[23]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d6_i0_i24 (.D(d6_71__N_1459[24]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d6_i0_i25 (.D(d6_71__N_1459[25]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d6_i0_i26 (.D(d6_71__N_1459[26]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d6_i0_i27 (.D(d6_71__N_1459[27]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d6_i0_i28 (.D(d6_71__N_1459[28]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d6_i0_i29 (.D(d6_71__N_1459[29]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d6_i0_i30 (.D(d6_71__N_1459[30]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d6_i0_i31 (.D(d6_71__N_1459[31]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d6_i0_i32 (.D(d6_71__N_1459[32]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d6_i0_i33 (.D(d6_71__N_1459[33]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d6_i0_i34 (.D(d6_71__N_1459[34]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d6_i0_i35 (.D(d6_71__N_1459[35]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d6_i0_i36 (.D(d6_71__N_1459[36]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d6_i0_i37 (.D(d6_71__N_1459[37]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d6_i0_i38 (.D(d6_71__N_1459[38]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d6_i0_i39 (.D(d6_71__N_1459[39]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d6_i0_i40 (.D(d6_71__N_1459[40]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d6_i0_i41 (.D(d6_71__N_1459[41]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d6_i0_i42 (.D(d6_71__N_1459[42]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d6_i0_i43 (.D(d6_71__N_1459[43]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d6_i0_i44 (.D(d6_71__N_1459[44]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d6_i0_i45 (.D(d6_71__N_1459[45]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d6_i0_i46 (.D(d6_71__N_1459[46]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d6_i0_i47 (.D(d6_71__N_1459[47]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d6_i0_i48 (.D(d6_71__N_1459[48]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d6_i0_i49 (.D(d6_71__N_1459[49]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d6_i0_i50 (.D(d6_71__N_1459[50]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d6_i0_i51 (.D(d6_71__N_1459[51]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d6_i0_i52 (.D(d6_71__N_1459[52]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d6_i0_i53 (.D(d6_71__N_1459[53]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d6_i0_i54 (.D(d6_71__N_1459[54]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d6_i0_i55 (.D(d6_71__N_1459[55]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d6_i0_i56 (.D(d6_71__N_1459[56]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d6_i0_i57 (.D(d6_71__N_1459[57]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d6_i0_i58 (.D(d6_71__N_1459[58]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d6_i0_i59 (.D(d6_71__N_1459[59]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d6_i0_i60 (.D(d6_71__N_1459[60]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d6_i0_i61 (.D(d6_71__N_1459[61]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d6_i0_i62 (.D(d6_71__N_1459[62]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d6_i0_i63 (.D(d6_71__N_1459[63]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d6_i0_i64 (.D(d6_71__N_1459[64]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d6_i0_i65 (.D(d6_71__N_1459[65]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d6_i0_i66 (.D(d6_71__N_1459[66]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d6_i0_i67 (.D(d6_71__N_1459[67]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d6_i0_i68 (.D(d6_71__N_1459[68]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d6_i0_i69 (.D(d6_71__N_1459[69]), .SP(osc_clk_enable_897), .CK(osc_clk), 
            .Q(d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d6_i0_i70 (.D(d6_71__N_1459[70]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d6_i0_i71 (.D(d6_71__N_1459[71]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i1 (.D(d6[1]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i2 (.D(d6[2]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i3 (.D(d6[3]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i4 (.D(d6[4]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i5 (.D(d6[5]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i6 (.D(d6[6]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i7 (.D(d6[7]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i8 (.D(d6[8]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i9 (.D(d6[9]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i10 (.D(d6[10]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i11 (.D(d6[11]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i12 (.D(d6[12]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i13 (.D(d6[13]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i14 (.D(d6[14]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i15 (.D(d6[15]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i16 (.D(d6[16]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i17 (.D(d6[17]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i18 (.D(d6[18]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i19 (.D(d6[19]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i20 (.D(d6[20]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i21 (.D(d6[21]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i22 (.D(d6[22]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i23 (.D(d6[23]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i24 (.D(d6[24]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i25 (.D(d6[25]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i26 (.D(d6[26]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i27 (.D(d6[27]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i28 (.D(d6[28]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i29 (.D(d6[29]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i30 (.D(d6[30]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i31 (.D(d6[31]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i32 (.D(d6[32]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i33 (.D(d6[33]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i34 (.D(d6[34]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i35 (.D(d6[35]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i36 (.D(d6[36]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i37 (.D(d6[37]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i38 (.D(d6[38]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i39 (.D(d6[39]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i40 (.D(d6[40]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i41 (.D(d6[41]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i42 (.D(d6[42]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i43 (.D(d6[43]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i44 (.D(d6[44]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i45 (.D(d6[45]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i46 (.D(d6[46]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i47 (.D(d6[47]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i48 (.D(d6[48]), .SP(osc_clk_enable_947), .CK(osc_clk), 
            .Q(d_d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i49 (.D(d6[49]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d_d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i50 (.D(d6[50]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d_d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i51 (.D(d6[51]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d_d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i52 (.D(d6[52]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d_d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i53 (.D(d6[53]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d_d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i54 (.D(d6[54]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d_d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i55 (.D(d6[55]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d_d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i56 (.D(d6[56]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d_d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i57 (.D(d6[57]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d_d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i58 (.D(d6[58]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d_d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i59 (.D(d6[59]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d_d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i60 (.D(d6[60]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d_d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i61 (.D(d6[61]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d_d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i62 (.D(d6[62]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d_d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i63 (.D(d6[63]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d_d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i64 (.D(d6[64]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d_d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i65 (.D(d6[65]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d_d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i66 (.D(d6[66]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d_d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i67 (.D(d6[67]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d_d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i68 (.D(d6[68]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d_d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i69 (.D(d6[69]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d_d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i70 (.D(d6[70]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d_d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i71 (.D(d6[71]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d_d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d7_i0_i1 (.D(d7_71__N_1531[1]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d7_i0_i2 (.D(d7_71__N_1531[2]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d7_i0_i3 (.D(d7_71__N_1531[3]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d7_i0_i4 (.D(d7_71__N_1531[4]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d7_i0_i5 (.D(d7_71__N_1531[5]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d7_i0_i6 (.D(d7_71__N_1531[6]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d7_i0_i7 (.D(d7_71__N_1531[7]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d7_i0_i8 (.D(d7_71__N_1531[8]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d7_i0_i9 (.D(d7_71__N_1531[9]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d7_i0_i10 (.D(d7_71__N_1531[10]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d7_i0_i11 (.D(d7_71__N_1531[11]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d7_i0_i12 (.D(d7_71__N_1531[12]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d7_i0_i13 (.D(d7_71__N_1531[13]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d7_i0_i14 (.D(d7_71__N_1531[14]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d7_i0_i15 (.D(d7_71__N_1531[15]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d7_i0_i16 (.D(d7_71__N_1531[16]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d7_i0_i17 (.D(d7_71__N_1531[17]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d7_i0_i18 (.D(d7_71__N_1531[18]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d7_i0_i19 (.D(d7_71__N_1531[19]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d7_i0_i20 (.D(d7_71__N_1531[20]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d7_i0_i21 (.D(d7_71__N_1531[21]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d7_i0_i22 (.D(d7_71__N_1531[22]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d7_i0_i23 (.D(d7_71__N_1531[23]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d7_i0_i24 (.D(d7_71__N_1531[24]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d7_i0_i25 (.D(d7_71__N_1531[25]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d7_i0_i26 (.D(d7_71__N_1531[26]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d7_i0_i27 (.D(d7_71__N_1531[27]), .SP(osc_clk_enable_997), .CK(osc_clk), 
            .Q(d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d7_i0_i28 (.D(d7_71__N_1531[28]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d7_i0_i29 (.D(d7_71__N_1531[29]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d7_i0_i30 (.D(d7_71__N_1531[30]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d7_i0_i31 (.D(d7_71__N_1531[31]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d7_i0_i32 (.D(d7_71__N_1531[32]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d7_i0_i33 (.D(d7_71__N_1531[33]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d7_i0_i34 (.D(d7_71__N_1531[34]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d7_i0_i35 (.D(d7_71__N_1531[35]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d7_i0_i36 (.D(d7_71__N_1531[36]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d7_i0_i37 (.D(d7_71__N_1531[37]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d7_i0_i38 (.D(d7_71__N_1531[38]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d7_i0_i39 (.D(d7_71__N_1531[39]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d7_i0_i40 (.D(d7_71__N_1531[40]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d7_i0_i41 (.D(d7_71__N_1531[41]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d7_i0_i42 (.D(d7_71__N_1531[42]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d7_i0_i43 (.D(d7_71__N_1531[43]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d7_i0_i44 (.D(d7_71__N_1531[44]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d7_i0_i45 (.D(d7_71__N_1531[45]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d7_i0_i46 (.D(d7_71__N_1531[46]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d7_i0_i47 (.D(d7_71__N_1531[47]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d7_i0_i48 (.D(d7_71__N_1531[48]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d7_i0_i49 (.D(d7_71__N_1531[49]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d7_i0_i50 (.D(d7_71__N_1531[50]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d7_i0_i51 (.D(d7_71__N_1531[51]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d7_i0_i52 (.D(d7_71__N_1531[52]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d7_i0_i53 (.D(d7_71__N_1531[53]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d7_i0_i54 (.D(d7_71__N_1531[54]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d7_i0_i55 (.D(d7_71__N_1531[55]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d7_i0_i56 (.D(d7_71__N_1531[56]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d7_i0_i57 (.D(d7_71__N_1531[57]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d7_i0_i58 (.D(d7_71__N_1531[58]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d7_i0_i59 (.D(d7_71__N_1531[59]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d7_i0_i60 (.D(d7_71__N_1531[60]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d7_i0_i61 (.D(d7_71__N_1531[61]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d7_i0_i62 (.D(d7_71__N_1531[62]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d7_i0_i63 (.D(d7_71__N_1531[63]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d7_i0_i64 (.D(d7_71__N_1531[64]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d7_i0_i65 (.D(d7_71__N_1531[65]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d7_i0_i66 (.D(d7_71__N_1531[66]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d7_i0_i67 (.D(d7_71__N_1531[67]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d7_i0_i68 (.D(d7_71__N_1531[68]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d7_i0_i69 (.D(d7_71__N_1531[69]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d7_i0_i70 (.D(d7_71__N_1531[70]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d7_i0_i71 (.D(d7_71__N_1531[71]), .SP(osc_clk_enable_1047), 
            .CK(osc_clk), .Q(d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i1 (.D(d7[1]), .SP(osc_clk_enable_1047), .CK(osc_clk), 
            .Q(d_d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i2 (.D(d7[2]), .SP(osc_clk_enable_1047), .CK(osc_clk), 
            .Q(d_d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i3 (.D(d7[3]), .SP(osc_clk_enable_1047), .CK(osc_clk), 
            .Q(d_d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i4 (.D(d7[4]), .SP(osc_clk_enable_1047), .CK(osc_clk), 
            .Q(d_d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i5 (.D(d7[5]), .SP(osc_clk_enable_1047), .CK(osc_clk), 
            .Q(d_d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i6 (.D(d7[6]), .SP(osc_clk_enable_1047), .CK(osc_clk), 
            .Q(d_d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i7 (.D(d7[7]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i8 (.D(d7[8]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i9 (.D(d7[9]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i10 (.D(d7[10]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i11 (.D(d7[11]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i12 (.D(d7[12]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i13 (.D(d7[13]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i14 (.D(d7[14]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i15 (.D(d7[15]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i16 (.D(d7[16]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i17 (.D(d7[17]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i18 (.D(d7[18]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i19 (.D(d7[19]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i20 (.D(d7[20]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i21 (.D(d7[21]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i22 (.D(d7[22]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i23 (.D(d7[23]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i24 (.D(d7[24]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i25 (.D(d7[25]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i26 (.D(d7[26]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i27 (.D(d7[27]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i28 (.D(d7[28]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i29 (.D(d7[29]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i30 (.D(d7[30]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i31 (.D(d7[31]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i32 (.D(d7[32]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i33 (.D(d7[33]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i34 (.D(d7[34]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i35 (.D(d7[35]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i36 (.D(d7[36]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i37 (.D(d7[37]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i38 (.D(d7[38]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i39 (.D(d7[39]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i40 (.D(d7[40]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i41 (.D(d7[41]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i42 (.D(d7[42]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i43 (.D(d7[43]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i44 (.D(d7[44]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i45 (.D(d7[45]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i46 (.D(d7[46]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i47 (.D(d7[47]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i48 (.D(d7[48]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i49 (.D(d7[49]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i50 (.D(d7[50]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i51 (.D(d7[51]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i52 (.D(d7[52]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i53 (.D(d7[53]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i54 (.D(d7[54]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i55 (.D(d7[55]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i56 (.D(d7[56]), .SP(osc_clk_enable_1097), .CK(osc_clk), 
            .Q(d_d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i57 (.D(d7[57]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d_d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i58 (.D(d7[58]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d_d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i59 (.D(d7[59]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d_d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i60 (.D(d7[60]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d_d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i61 (.D(d7[61]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d_d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i62 (.D(d7[62]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d_d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i63 (.D(d7[63]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d_d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i64 (.D(d7[64]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d_d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i65 (.D(d7[65]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d_d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i66 (.D(d7[66]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d_d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i67 (.D(d7[67]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d_d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i68 (.D(d7[68]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d_d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i69 (.D(d7[69]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d_d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i70 (.D(d7[70]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d_d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i71 (.D(d7[71]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d_d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d8_i0_i1 (.D(d8_71__N_1603[1]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d8_i0_i2 (.D(d8_71__N_1603[2]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d8_i0_i3 (.D(d8_71__N_1603[3]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d8_i0_i4 (.D(d8_71__N_1603[4]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d8_i0_i5 (.D(d8_71__N_1603[5]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d8_i0_i6 (.D(d8_71__N_1603[6]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d8_i0_i7 (.D(d8_71__N_1603[7]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d8_i0_i8 (.D(d8_71__N_1603[8]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d8_i0_i9 (.D(d8_71__N_1603[9]), .SP(osc_clk_enable_1147), .CK(osc_clk), 
            .Q(d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d8_i0_i10 (.D(d8_71__N_1603[10]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d8_i0_i11 (.D(d8_71__N_1603[11]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d8_i0_i12 (.D(d8_71__N_1603[12]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d8_i0_i13 (.D(d8_71__N_1603[13]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d8_i0_i14 (.D(d8_71__N_1603[14]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d8_i0_i15 (.D(d8_71__N_1603[15]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d8_i0_i16 (.D(d8_71__N_1603[16]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d8_i0_i17 (.D(d8_71__N_1603[17]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d8_i0_i18 (.D(d8_71__N_1603[18]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d8_i0_i19 (.D(d8_71__N_1603[19]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d8_i0_i20 (.D(d8_71__N_1603[20]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d8_i0_i21 (.D(d8_71__N_1603[21]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d8_i0_i22 (.D(d8_71__N_1603[22]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d8_i0_i23 (.D(d8_71__N_1603[23]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d8_i0_i24 (.D(d8_71__N_1603[24]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d8_i0_i25 (.D(d8_71__N_1603[25]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d8_i0_i26 (.D(d8_71__N_1603[26]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d8_i0_i27 (.D(d8_71__N_1603[27]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d8_i0_i28 (.D(d8_71__N_1603[28]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d8_i0_i29 (.D(d8_71__N_1603[29]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d8_i0_i30 (.D(d8_71__N_1603[30]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d8_i0_i31 (.D(d8_71__N_1603[31]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d8_i0_i32 (.D(d8_71__N_1603[32]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d8_i0_i33 (.D(d8_71__N_1603[33]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d8_i0_i34 (.D(d8_71__N_1603[34]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d8_i0_i35 (.D(d8_71__N_1603[35]), .SP(osc_clk_enable_1147), 
            .CK(osc_clk), .Q(d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d8_i0_i36 (.D(d8_71__N_1603[36]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d8_i0_i37 (.D(d8_71__N_1603[37]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d8_i0_i38 (.D(d8_71__N_1603[38]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d8_i0_i39 (.D(d8_71__N_1603[39]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d8_i0_i40 (.D(d8_71__N_1603[40]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d8_i0_i41 (.D(d8_71__N_1603[41]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d8_i0_i42 (.D(d8_71__N_1603[42]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d8_i0_i43 (.D(d8_71__N_1603[43]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d8_i0_i44 (.D(d8_71__N_1603[44]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d8_i0_i45 (.D(d8_71__N_1603[45]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d8_i0_i46 (.D(d8_71__N_1603[46]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d8_i0_i47 (.D(d8_71__N_1603[47]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d8_i0_i48 (.D(d8_71__N_1603[48]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d8_i0_i49 (.D(d8_71__N_1603[49]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d8_i0_i50 (.D(d8_71__N_1603[50]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d8_i0_i51 (.D(d8_71__N_1603[51]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d8_i0_i52 (.D(d8_71__N_1603[52]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d8_i0_i53 (.D(d8_71__N_1603[53]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d8_i0_i54 (.D(d8_71__N_1603[54]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d8_i0_i55 (.D(d8_71__N_1603[55]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d8_i0_i56 (.D(d8_71__N_1603[56]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d8_i0_i57 (.D(d8_71__N_1603[57]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d8_i0_i58 (.D(d8_71__N_1603[58]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d8_i0_i59 (.D(d8_71__N_1603[59]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d8_i0_i60 (.D(d8_71__N_1603[60]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d8_i0_i61 (.D(d8_71__N_1603[61]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d8_i0_i62 (.D(d8_71__N_1603[62]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d8_i0_i63 (.D(d8_71__N_1603[63]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d8_i0_i64 (.D(d8_71__N_1603[64]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d8_i0_i65 (.D(d8_71__N_1603[65]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d8_i0_i66 (.D(d8_71__N_1603[66]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d8_i0_i67 (.D(d8_71__N_1603[67]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d8_i0_i68 (.D(d8_71__N_1603[68]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d8_i0_i69 (.D(d8_71__N_1603[69]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d8_i0_i70 (.D(d8_71__N_1603[70]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d8_i0_i71 (.D(d8_71__N_1603[71]), .SP(osc_clk_enable_1197), 
            .CK(osc_clk), .Q(d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i1 (.D(d8[1]), .SP(osc_clk_enable_1197), .CK(osc_clk), 
            .Q(d_d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i2 (.D(d8[2]), .SP(osc_clk_enable_1197), .CK(osc_clk), 
            .Q(d_d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i3 (.D(d8[3]), .SP(osc_clk_enable_1197), .CK(osc_clk), 
            .Q(d_d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i4 (.D(d8[4]), .SP(osc_clk_enable_1197), .CK(osc_clk), 
            .Q(d_d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i5 (.D(d8[5]), .SP(osc_clk_enable_1197), .CK(osc_clk), 
            .Q(d_d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i6 (.D(d8[6]), .SP(osc_clk_enable_1197), .CK(osc_clk), 
            .Q(d_d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i7 (.D(d8[7]), .SP(osc_clk_enable_1197), .CK(osc_clk), 
            .Q(d_d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i8 (.D(d8[8]), .SP(osc_clk_enable_1197), .CK(osc_clk), 
            .Q(d_d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i9 (.D(d8[9]), .SP(osc_clk_enable_1197), .CK(osc_clk), 
            .Q(d_d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i10 (.D(d8[10]), .SP(osc_clk_enable_1197), .CK(osc_clk), 
            .Q(d_d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i11 (.D(d8[11]), .SP(osc_clk_enable_1197), .CK(osc_clk), 
            .Q(d_d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i12 (.D(d8[12]), .SP(osc_clk_enable_1197), .CK(osc_clk), 
            .Q(d_d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i13 (.D(d8[13]), .SP(osc_clk_enable_1197), .CK(osc_clk), 
            .Q(d_d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i14 (.D(d8[14]), .SP(osc_clk_enable_1197), .CK(osc_clk), 
            .Q(d_d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i15 (.D(d8[15]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i16 (.D(d8[16]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i17 (.D(d8[17]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i18 (.D(d8[18]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i19 (.D(d8[19]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i20 (.D(d8[20]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i21 (.D(d8[21]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i22 (.D(d8[22]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i23 (.D(d8[23]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i24 (.D(d8[24]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i25 (.D(d8[25]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i26 (.D(d8[26]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i27 (.D(d8[27]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i28 (.D(d8[28]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i29 (.D(d8[29]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i30 (.D(d8[30]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i31 (.D(d8[31]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i32 (.D(d8[32]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i33 (.D(d8[33]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i34 (.D(d8[34]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i35 (.D(d8[35]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i36 (.D(d8[36]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i37 (.D(d8[37]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i38 (.D(d8[38]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i39 (.D(d8[39]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i40 (.D(d8[40]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i41 (.D(d8[41]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i42 (.D(d8[42]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i43 (.D(d8[43]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i44 (.D(d8[44]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i45 (.D(d8[45]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i46 (.D(d8[46]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i47 (.D(d8[47]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i48 (.D(d8[48]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i49 (.D(d8[49]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i50 (.D(d8[50]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i51 (.D(d8[51]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i52 (.D(d8[52]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i53 (.D(d8[53]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i54 (.D(d8[54]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i55 (.D(d8[55]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i56 (.D(d8[56]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i57 (.D(d8[57]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i58 (.D(d8[58]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i59 (.D(d8[59]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i60 (.D(d8[60]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i61 (.D(d8[61]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i62 (.D(d8[62]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i63 (.D(d8[63]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i64 (.D(d8[64]), .SP(osc_clk_enable_1247), .CK(osc_clk), 
            .Q(d_d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i65 (.D(d8[65]), .SP(osc_clk_enable_1297), .CK(osc_clk), 
            .Q(d_d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i66 (.D(d8[66]), .SP(osc_clk_enable_1297), .CK(osc_clk), 
            .Q(d_d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i67 (.D(d8[67]), .SP(osc_clk_enable_1297), .CK(osc_clk), 
            .Q(d_d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i68 (.D(d8[68]), .SP(osc_clk_enable_1297), .CK(osc_clk), 
            .Q(d_d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i69 (.D(d8[69]), .SP(osc_clk_enable_1297), .CK(osc_clk), 
            .Q(d_d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i70 (.D(d8[70]), .SP(osc_clk_enable_1297), .CK(osc_clk), 
            .Q(d_d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i71 (.D(d8[71]), .SP(osc_clk_enable_1297), .CK(osc_clk), 
            .Q(d_d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d9_i0_i1 (.D(d9_71__N_1675[1]), .SP(osc_clk_enable_1297), .CK(osc_clk), 
            .Q(d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d9_i0_i2 (.D(d9_71__N_1675[2]), .SP(osc_clk_enable_1297), .CK(osc_clk), 
            .Q(d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d9_i0_i3 (.D(d9_71__N_1675[3]), .SP(osc_clk_enable_1297), .CK(osc_clk), 
            .Q(d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d9_i0_i4 (.D(d9_71__N_1675[4]), .SP(osc_clk_enable_1297), .CK(osc_clk), 
            .Q(d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d9_i0_i5 (.D(d9_71__N_1675[5]), .SP(osc_clk_enable_1297), .CK(osc_clk), 
            .Q(d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d9_i0_i6 (.D(d9_71__N_1675[6]), .SP(osc_clk_enable_1297), .CK(osc_clk), 
            .Q(d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d9_i0_i7 (.D(d9_71__N_1675[7]), .SP(osc_clk_enable_1297), .CK(osc_clk), 
            .Q(d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d9_i0_i8 (.D(d9_71__N_1675[8]), .SP(osc_clk_enable_1297), .CK(osc_clk), 
            .Q(d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d9_i0_i9 (.D(d9_71__N_1675[9]), .SP(osc_clk_enable_1297), .CK(osc_clk), 
            .Q(d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d9_i0_i10 (.D(d9_71__N_1675[10]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d9_i0_i11 (.D(d9_71__N_1675[11]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d9_i0_i12 (.D(d9_71__N_1675[12]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d9_i0_i13 (.D(d9_71__N_1675[13]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d9_i0_i14 (.D(d9_71__N_1675[14]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d9_i0_i15 (.D(d9_71__N_1675[15]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d9_i0_i16 (.D(d9_71__N_1675[16]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d9_i0_i17 (.D(d9_71__N_1675[17]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d9_i0_i18 (.D(d9_71__N_1675[18]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d9_i0_i19 (.D(d9_71__N_1675[19]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d9_i0_i20 (.D(d9_71__N_1675[20]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d9_i0_i21 (.D(d9_71__N_1675[21]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d9_i0_i22 (.D(d9_71__N_1675[22]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d9_i0_i23 (.D(d9_71__N_1675[23]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d9_i0_i24 (.D(d9_71__N_1675[24]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d9_i0_i25 (.D(d9_71__N_1675[25]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d9_i0_i26 (.D(d9_71__N_1675[26]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d9_i0_i27 (.D(d9_71__N_1675[27]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d9_i0_i28 (.D(d9_71__N_1675[28]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d9_i0_i29 (.D(d9_71__N_1675[29]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d9_i0_i30 (.D(d9_71__N_1675[30]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d9_i0_i31 (.D(d9_71__N_1675[31]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d9_i0_i32 (.D(d9_71__N_1675[32]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d9_i0_i33 (.D(d9_71__N_1675[33]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d9_i0_i34 (.D(d9_71__N_1675[34]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d9_i0_i35 (.D(d9_71__N_1675[35]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d9_i0_i36 (.D(d9_71__N_1675[36]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d9_i0_i37 (.D(d9_71__N_1675[37]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d9_i0_i38 (.D(d9_71__N_1675[38]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d9_i0_i39 (.D(d9_71__N_1675[39]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d9_i0_i40 (.D(d9_71__N_1675[40]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d9_i0_i41 (.D(d9_71__N_1675[41]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d9_i0_i42 (.D(d9_71__N_1675[42]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d9_i0_i43 (.D(d9_71__N_1675[43]), .SP(osc_clk_enable_1297), 
            .CK(osc_clk), .Q(d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d9_i0_i44 (.D(d9_71__N_1675[44]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d9_i0_i45 (.D(d9_71__N_1675[45]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d9_i0_i46 (.D(d9_71__N_1675[46]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d9_i0_i47 (.D(d9_71__N_1675[47]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d9_i0_i48 (.D(d9_71__N_1675[48]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d9_i0_i49 (.D(d9_71__N_1675[49]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d9_i0_i50 (.D(d9_71__N_1675[50]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d9_i0_i51 (.D(d9_71__N_1675[51]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d9_i0_i52 (.D(d9_71__N_1675[52]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d9_i0_i53 (.D(d9_71__N_1675[53]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d9_i0_i54 (.D(d9_71__N_1675[54]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d9_i0_i55 (.D(d9_71__N_1675[55]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d9_i0_i56 (.D(d9_71__N_1675[56]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d9_i0_i57 (.D(d9_71__N_1675[57]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d9_i0_i58 (.D(d9_71__N_1675[58]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d9_i0_i59 (.D(d9_71__N_1675[59]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d9_i0_i60 (.D(d9_71__N_1675[60]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d9_i0_i61 (.D(d9_71__N_1675[61]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d9_i0_i62 (.D(d9_71__N_1675[62]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d9_i0_i63 (.D(d9_71__N_1675[63]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d9_i0_i64 (.D(d9_71__N_1675[64]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d9_i0_i65 (.D(d9_71__N_1675[65]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d9_i0_i66 (.D(d9_71__N_1675[66]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d9_i0_i67 (.D(d9_71__N_1675[67]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d9_i0_i68 (.D(d9_71__N_1675[68]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d9_i0_i69 (.D(d9_71__N_1675[69]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d9_i0_i70 (.D(d9_71__N_1675[70]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d9_i0_i71 (.D(d9_71__N_1675[71]), .SP(osc_clk_enable_1347), 
            .CK(osc_clk), .Q(d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i1 (.D(d9[1]), .SP(osc_clk_enable_1347), .CK(osc_clk), 
            .Q(d_d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i2 (.D(d9[2]), .SP(osc_clk_enable_1347), .CK(osc_clk), 
            .Q(d_d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i3 (.D(d9[3]), .SP(osc_clk_enable_1347), .CK(osc_clk), 
            .Q(d_d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i4 (.D(d9[4]), .SP(osc_clk_enable_1347), .CK(osc_clk), 
            .Q(d_d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i5 (.D(d9[5]), .SP(osc_clk_enable_1347), .CK(osc_clk), 
            .Q(d_d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i6 (.D(d9[6]), .SP(osc_clk_enable_1347), .CK(osc_clk), 
            .Q(d_d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i7 (.D(d9[7]), .SP(osc_clk_enable_1347), .CK(osc_clk), 
            .Q(d_d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i8 (.D(d9[8]), .SP(osc_clk_enable_1347), .CK(osc_clk), 
            .Q(d_d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i9 (.D(d9[9]), .SP(osc_clk_enable_1347), .CK(osc_clk), 
            .Q(d_d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i10 (.D(d9[10]), .SP(osc_clk_enable_1347), .CK(osc_clk), 
            .Q(d_d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i11 (.D(d9[11]), .SP(osc_clk_enable_1347), .CK(osc_clk), 
            .Q(d_d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i12 (.D(d9[12]), .SP(osc_clk_enable_1347), .CK(osc_clk), 
            .Q(d_d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i13 (.D(d9[13]), .SP(osc_clk_enable_1347), .CK(osc_clk), 
            .Q(d_d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i14 (.D(d9[14]), .SP(osc_clk_enable_1347), .CK(osc_clk), 
            .Q(d_d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i15 (.D(d9[15]), .SP(osc_clk_enable_1347), .CK(osc_clk), 
            .Q(d_d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i16 (.D(d9[16]), .SP(osc_clk_enable_1347), .CK(osc_clk), 
            .Q(d_d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i17 (.D(d9[17]), .SP(osc_clk_enable_1347), .CK(osc_clk), 
            .Q(d_d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i18 (.D(d9[18]), .SP(osc_clk_enable_1347), .CK(osc_clk), 
            .Q(d_d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i19 (.D(d9[19]), .SP(osc_clk_enable_1347), .CK(osc_clk), 
            .Q(d_d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i20 (.D(d9[20]), .SP(osc_clk_enable_1347), .CK(osc_clk), 
            .Q(d_d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i21 (.D(d9[21]), .SP(osc_clk_enable_1347), .CK(osc_clk), 
            .Q(d_d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i22 (.D(d9[22]), .SP(osc_clk_enable_1347), .CK(osc_clk), 
            .Q(d_d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i23 (.D(d9[23]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i24 (.D(d9[24]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i25 (.D(d9[25]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i26 (.D(d9[26]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i27 (.D(d9[27]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i28 (.D(d9[28]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i29 (.D(d9[29]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i30 (.D(d9[30]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i31 (.D(d9[31]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i32 (.D(d9[32]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i33 (.D(d9[33]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i34 (.D(d9[34]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i35 (.D(d9[35]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i36 (.D(d9[36]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i37 (.D(d9[37]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i38 (.D(d9[38]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i39 (.D(d9[39]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i40 (.D(d9[40]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i41 (.D(d9[41]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i42 (.D(d9[42]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i43 (.D(d9[43]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i44 (.D(d9[44]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i45 (.D(d9[45]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i46 (.D(d9[46]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i47 (.D(d9[47]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i48 (.D(d9[48]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i49 (.D(d9[49]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i50 (.D(d9[50]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i51 (.D(d9[51]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i52 (.D(d9[52]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i53 (.D(d9[53]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i54 (.D(d9[54]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i55 (.D(d9[55]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i56 (.D(d9[56]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i57 (.D(d9[57]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i58 (.D(d9[58]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i59 (.D(d9[59]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i60 (.D(d9[60]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i61 (.D(d9[61]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i62 (.D(d9[62]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i63 (.D(d9[63]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i64 (.D(d9[64]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i65 (.D(d9[65]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i66 (.D(d9[66]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i67 (.D(d9[67]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i68 (.D(d9[68]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i69 (.D(d9[69]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i70 (.D(d9[70]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i71 (.D(d9[71]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d_d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d10__i2 (.D(d10_71__N_1747[57]), .SP(osc_clk_enable_1397), .CK(osc_clk), 
            .Q(d10[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i2.GSR = "ENABLED";
    FD1P3AX d10__i3 (.D(d10_71__N_1747[58]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i3.GSR = "ENABLED";
    FD1P3AX d10__i4 (.D(d10_71__N_1747[59]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[59] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i4.GSR = "ENABLED";
    FD1P3AX d10__i5 (.D(d10_71__N_1747[60]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[60] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i5.GSR = "ENABLED";
    FD1P3AX d10__i6 (.D(d10_71__N_1747[61]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[61] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i6.GSR = "ENABLED";
    FD1P3AX d10__i7 (.D(d10_71__N_1747[62]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[62] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i7.GSR = "ENABLED";
    FD1P3AX d10__i8 (.D(d10_71__N_1747[63]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[63] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i8.GSR = "ENABLED";
    FD1P3AX d10__i9 (.D(d10_71__N_1747[64]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[64] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i9.GSR = "ENABLED";
    FD1P3AX d10__i10 (.D(d10_71__N_1747[65]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[65] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i10.GSR = "ENABLED";
    FD1P3AX d10__i11 (.D(d10_71__N_1747[66]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[66] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i11.GSR = "ENABLED";
    FD1P3AX d10__i12 (.D(d10_71__N_1747[67]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[67] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i12.GSR = "ENABLED";
    FD1P3AX d10__i13 (.D(d10_71__N_1747[68]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[68] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i13.GSR = "ENABLED";
    FD1P3AX d10__i14 (.D(d10_71__N_1747[69]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[69] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i14.GSR = "ENABLED";
    FD1P3AX d10__i15 (.D(d10_71__N_1747[70]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[70] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i15.GSR = "ENABLED";
    FD1P3AX d10__i16 (.D(d10_71__N_1747[71]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[71] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i16.GSR = "ENABLED";
    FD1P3AX d_out_i0_i1 (.D(d_out_11__N_1819[1]), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i1.GSR = "ENABLED";
    FD1P3AX d_out_i0_i2 (.D(\d_out_11__N_1819[2] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i2.GSR = "ENABLED";
    FD1P3AX d_out_i0_i3 (.D(\d_out_11__N_1819[3] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i3.GSR = "ENABLED";
    FD1P3AX d_out_i0_i4 (.D(\d_out_11__N_1819[4] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i4.GSR = "ENABLED";
    FD1P3AX d_out_i0_i5 (.D(\d_out_11__N_1819[5] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i5.GSR = "ENABLED";
    FD1P3AX d_out_i0_i6 (.D(\d_out_11__N_1819[6] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i6.GSR = "ENABLED";
    FD1P3AX d_out_i0_i7 (.D(\d_out_11__N_1819[7] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i7.GSR = "ENABLED";
    FD1P3AX d_out_i0_i8 (.D(\d_out_11__N_1819[8] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i8.GSR = "ENABLED";
    FD1P3AX d_out_i0_i9 (.D(\d_out_11__N_1819[9] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i9.GSR = "ENABLED";
    FD1P3AX d_out_i0_i10 (.D(\d_out_11__N_1819[10] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i10.GSR = "ENABLED";
    FD1P3AX d_out_i0_i11 (.D(\d_out_11__N_1819[11] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i11.GSR = "ENABLED";
    FD1S3AX d1_i1 (.D(d1_71__N_418[1]), .CK(osc_clk), .Q(d1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i1.GSR = "ENABLED";
    FD1S3AX d1_i2 (.D(d1_71__N_418[2]), .CK(osc_clk), .Q(d1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i2.GSR = "ENABLED";
    FD1S3AX d1_i3 (.D(d1_71__N_418[3]), .CK(osc_clk), .Q(d1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i3.GSR = "ENABLED";
    FD1S3AX d1_i4 (.D(d1_71__N_418[4]), .CK(osc_clk), .Q(d1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i4.GSR = "ENABLED";
    FD1S3AX d1_i5 (.D(d1_71__N_418[5]), .CK(osc_clk), .Q(d1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i5.GSR = "ENABLED";
    FD1S3AX d1_i6 (.D(d1_71__N_418[6]), .CK(osc_clk), .Q(d1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i6.GSR = "ENABLED";
    FD1S3AX d1_i7 (.D(d1_71__N_418[7]), .CK(osc_clk), .Q(d1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i7.GSR = "ENABLED";
    FD1S3AX d1_i8 (.D(d1_71__N_418[8]), .CK(osc_clk), .Q(d1[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i8.GSR = "ENABLED";
    FD1S3AX d1_i9 (.D(d1_71__N_418[9]), .CK(osc_clk), .Q(d1[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i9.GSR = "ENABLED";
    FD1S3AX d1_i10 (.D(d1_71__N_418[10]), .CK(osc_clk), .Q(d1[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i10.GSR = "ENABLED";
    FD1S3AX d1_i11 (.D(d1_71__N_418[11]), .CK(osc_clk), .Q(d1[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i11.GSR = "ENABLED";
    FD1S3AX d1_i12 (.D(d1_71__N_418[12]), .CK(osc_clk), .Q(d1[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i12.GSR = "ENABLED";
    FD1S3AX d1_i13 (.D(d1_71__N_418[13]), .CK(osc_clk), .Q(d1[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i13.GSR = "ENABLED";
    FD1S3AX d1_i14 (.D(d1_71__N_418[14]), .CK(osc_clk), .Q(d1[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i14.GSR = "ENABLED";
    FD1S3AX d1_i15 (.D(d1_71__N_418[15]), .CK(osc_clk), .Q(d1[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i15.GSR = "ENABLED";
    FD1S3AX d1_i16 (.D(d1_71__N_418[16]), .CK(osc_clk), .Q(d1[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i16.GSR = "ENABLED";
    FD1S3AX d1_i17 (.D(d1_71__N_418[17]), .CK(osc_clk), .Q(d1[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i17.GSR = "ENABLED";
    FD1S3AX d1_i18 (.D(d1_71__N_418[18]), .CK(osc_clk), .Q(d1[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i18.GSR = "ENABLED";
    FD1S3AX d1_i19 (.D(d1_71__N_418[19]), .CK(osc_clk), .Q(d1[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i19.GSR = "ENABLED";
    FD1S3AX d1_i20 (.D(d1_71__N_418[20]), .CK(osc_clk), .Q(d1[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i20.GSR = "ENABLED";
    FD1S3AX d1_i21 (.D(d1_71__N_418[21]), .CK(osc_clk), .Q(d1[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i21.GSR = "ENABLED";
    FD1S3AX d1_i22 (.D(d1_71__N_418[22]), .CK(osc_clk), .Q(d1[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i22.GSR = "ENABLED";
    FD1S3AX d1_i23 (.D(d1_71__N_418[23]), .CK(osc_clk), .Q(d1[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i23.GSR = "ENABLED";
    FD1S3AX d1_i24 (.D(d1_71__N_418[24]), .CK(osc_clk), .Q(d1[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i24.GSR = "ENABLED";
    FD1S3AX d1_i25 (.D(d1_71__N_418[25]), .CK(osc_clk), .Q(d1[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i25.GSR = "ENABLED";
    FD1S3AX d1_i26 (.D(d1_71__N_418[26]), .CK(osc_clk), .Q(d1[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i26.GSR = "ENABLED";
    FD1S3AX d1_i27 (.D(d1_71__N_418[27]), .CK(osc_clk), .Q(d1[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i27.GSR = "ENABLED";
    FD1S3AX d1_i28 (.D(d1_71__N_418[28]), .CK(osc_clk), .Q(d1[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i28.GSR = "ENABLED";
    FD1S3AX d1_i29 (.D(d1_71__N_418[29]), .CK(osc_clk), .Q(d1[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i29.GSR = "ENABLED";
    FD1S3AX d1_i30 (.D(d1_71__N_418[30]), .CK(osc_clk), .Q(d1[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i30.GSR = "ENABLED";
    FD1S3AX d1_i31 (.D(d1_71__N_418[31]), .CK(osc_clk), .Q(d1[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i31.GSR = "ENABLED";
    FD1S3AX d1_i32 (.D(d1_71__N_418[32]), .CK(osc_clk), .Q(d1[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i32.GSR = "ENABLED";
    FD1S3AX d1_i33 (.D(d1_71__N_418[33]), .CK(osc_clk), .Q(d1[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i33.GSR = "ENABLED";
    FD1S3AX d1_i34 (.D(d1_71__N_418[34]), .CK(osc_clk), .Q(d1[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i34.GSR = "ENABLED";
    FD1S3AX d1_i35 (.D(d1_71__N_418[35]), .CK(osc_clk), .Q(d1[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i35.GSR = "ENABLED";
    FD1S3AX d1_i36 (.D(d1_71__N_418[36]), .CK(osc_clk), .Q(d1[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i36.GSR = "ENABLED";
    FD1S3AX d1_i37 (.D(d1_71__N_418[37]), .CK(osc_clk), .Q(d1[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i37.GSR = "ENABLED";
    FD1S3AX d1_i38 (.D(d1_71__N_418[38]), .CK(osc_clk), .Q(d1[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i38.GSR = "ENABLED";
    FD1S3AX d1_i39 (.D(d1_71__N_418[39]), .CK(osc_clk), .Q(d1[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i39.GSR = "ENABLED";
    FD1S3AX d1_i40 (.D(d1_71__N_418[40]), .CK(osc_clk), .Q(d1[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i40.GSR = "ENABLED";
    FD1S3AX d1_i41 (.D(d1_71__N_418[41]), .CK(osc_clk), .Q(d1[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i41.GSR = "ENABLED";
    FD1S3AX d1_i42 (.D(d1_71__N_418[42]), .CK(osc_clk), .Q(d1[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i42.GSR = "ENABLED";
    FD1S3AX d1_i43 (.D(d1_71__N_418[43]), .CK(osc_clk), .Q(d1[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i43.GSR = "ENABLED";
    FD1S3AX d1_i44 (.D(d1_71__N_418[44]), .CK(osc_clk), .Q(d1[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i44.GSR = "ENABLED";
    FD1S3AX d1_i45 (.D(d1_71__N_418[45]), .CK(osc_clk), .Q(d1[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i45.GSR = "ENABLED";
    FD1S3AX d1_i46 (.D(d1_71__N_418[46]), .CK(osc_clk), .Q(d1[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i46.GSR = "ENABLED";
    FD1S3AX d1_i47 (.D(d1_71__N_418[47]), .CK(osc_clk), .Q(d1[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i47.GSR = "ENABLED";
    FD1S3AX d1_i48 (.D(d1_71__N_418[48]), .CK(osc_clk), .Q(d1[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i48.GSR = "ENABLED";
    FD1S3AX d1_i49 (.D(d1_71__N_418[49]), .CK(osc_clk), .Q(d1[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i49.GSR = "ENABLED";
    FD1S3AX d1_i50 (.D(d1_71__N_418[50]), .CK(osc_clk), .Q(d1[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i50.GSR = "ENABLED";
    FD1S3AX d1_i51 (.D(d1_71__N_418[51]), .CK(osc_clk), .Q(d1[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i51.GSR = "ENABLED";
    FD1S3AX d1_i52 (.D(d1_71__N_418[52]), .CK(osc_clk), .Q(d1[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i52.GSR = "ENABLED";
    FD1S3AX d1_i53 (.D(d1_71__N_418[53]), .CK(osc_clk), .Q(d1[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i53.GSR = "ENABLED";
    FD1S3AX d1_i54 (.D(d1_71__N_418[54]), .CK(osc_clk), .Q(d1[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i54.GSR = "ENABLED";
    FD1S3AX d1_i55 (.D(d1_71__N_418[55]), .CK(osc_clk), .Q(d1[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i55.GSR = "ENABLED";
    FD1S3AX d1_i56 (.D(d1_71__N_418[56]), .CK(osc_clk), .Q(d1[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i56.GSR = "ENABLED";
    FD1S3AX d1_i57 (.D(d1_71__N_418[57]), .CK(osc_clk), .Q(d1[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i57.GSR = "ENABLED";
    FD1S3AX d1_i58 (.D(d1_71__N_418[58]), .CK(osc_clk), .Q(d1[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i58.GSR = "ENABLED";
    FD1S3AX d1_i59 (.D(d1_71__N_418[59]), .CK(osc_clk), .Q(d1[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i59.GSR = "ENABLED";
    FD1S3AX d1_i60 (.D(d1_71__N_418[60]), .CK(osc_clk), .Q(d1[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i60.GSR = "ENABLED";
    FD1S3AX d1_i61 (.D(d1_71__N_418[61]), .CK(osc_clk), .Q(d1[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i61.GSR = "ENABLED";
    FD1S3AX d1_i62 (.D(d1_71__N_418[62]), .CK(osc_clk), .Q(d1[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i62.GSR = "ENABLED";
    FD1S3AX d1_i63 (.D(d1_71__N_418[63]), .CK(osc_clk), .Q(d1[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i63.GSR = "ENABLED";
    FD1S3AX d1_i64 (.D(d1_71__N_418[64]), .CK(osc_clk), .Q(d1[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i64.GSR = "ENABLED";
    FD1S3AX d1_i65 (.D(d1_71__N_418[65]), .CK(osc_clk), .Q(d1[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i65.GSR = "ENABLED";
    FD1S3AX d1_i66 (.D(d1_71__N_418[66]), .CK(osc_clk), .Q(d1[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i66.GSR = "ENABLED";
    FD1S3AX d1_i67 (.D(d1_71__N_418[67]), .CK(osc_clk), .Q(d1[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i67.GSR = "ENABLED";
    FD1S3AX d1_i68 (.D(d1_71__N_418[68]), .CK(osc_clk), .Q(d1[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i68.GSR = "ENABLED";
    FD1S3AX d1_i69 (.D(d1_71__N_418[69]), .CK(osc_clk), .Q(d1[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i69.GSR = "ENABLED";
    FD1S3AX d1_i70 (.D(d1_71__N_418[70]), .CK(osc_clk), .Q(d1[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i70.GSR = "ENABLED";
    FD1S3AX d1_i71 (.D(d1_71__N_418[71]), .CK(osc_clk), .Q(d1[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i71.GSR = "ENABLED";
    CCU2D add_1111_9 (.A0(d_tmp[43]), .B0(d_d_tmp[43]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[44]), .B1(d_d_tmp[44]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11316), .COUT(n11317), .S0(n6124[7]), 
          .S1(n6124[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1111_9.INIT0 = 16'h5999;
    defparam add_1111_9.INIT1 = 16'h5999;
    defparam add_1111_9.INJECT1_0 = "NO";
    defparam add_1111_9.INJECT1_1 = "NO";
    CCU2D add_1111_7 (.A0(d_tmp[41]), .B0(d_d_tmp[41]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[42]), .B1(d_d_tmp[42]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11315), .COUT(n11316), .S0(n6124[5]), 
          .S1(n6124[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1111_7.INIT0 = 16'h5999;
    defparam add_1111_7.INIT1 = 16'h5999;
    defparam add_1111_7.INJECT1_0 = "NO";
    defparam add_1111_7.INJECT1_1 = "NO";
    CCU2D add_1111_5 (.A0(d_tmp[39]), .B0(d_d_tmp[39]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[40]), .B1(d_d_tmp[40]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11314), .COUT(n11315), .S0(n6124[3]), 
          .S1(n6124[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1111_5.INIT0 = 16'h5999;
    defparam add_1111_5.INIT1 = 16'h5999;
    defparam add_1111_5.INJECT1_0 = "NO";
    defparam add_1111_5.INJECT1_1 = "NO";
    CCU2D add_1111_3 (.A0(d_tmp[37]), .B0(d_d_tmp[37]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[38]), .B1(d_d_tmp[38]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11313), .COUT(n11314), .S0(n6124[1]), 
          .S1(n6124[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1111_3.INIT0 = 16'h5999;
    defparam add_1111_3.INIT1 = 16'h5999;
    defparam add_1111_3.INJECT1_0 = "NO";
    defparam add_1111_3.INJECT1_1 = "NO";
    CCU2D add_1111_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[36]), .B1(d_d_tmp[36]), .C1(GND_net), .D1(GND_net), 
          .COUT(n11313), .S1(n6124[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1111_1.INIT0 = 16'hF000;
    defparam add_1111_1.INIT1 = 16'h5999;
    defparam add_1111_1.INJECT1_0 = "NO";
    defparam add_1111_1.INJECT1_1 = "NO";
    CCU2D add_1112_37 (.A0(d_d_tmp[70]), .B0(n6123), .C0(n6124[34]), .D0(d_tmp[70]), 
          .A1(d_d_tmp[71]), .B1(n6123), .C1(n6124[35]), .D1(d_tmp[71]), 
          .CIN(n11311), .S0(d6_71__N_1459[70]), .S1(d6_71__N_1459[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1112_37.INIT0 = 16'hb874;
    defparam add_1112_37.INIT1 = 16'hb874;
    defparam add_1112_37.INJECT1_0 = "NO";
    defparam add_1112_37.INJECT1_1 = "NO";
    CCU2D add_1112_35 (.A0(d_d_tmp[68]), .B0(n6123), .C0(n6124[32]), .D0(d_tmp[68]), 
          .A1(d_d_tmp[69]), .B1(n6123), .C1(n6124[33]), .D1(d_tmp[69]), 
          .CIN(n11310), .COUT(n11311), .S0(d6_71__N_1459[68]), .S1(d6_71__N_1459[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1112_35.INIT0 = 16'hb874;
    defparam add_1112_35.INIT1 = 16'hb874;
    defparam add_1112_35.INJECT1_0 = "NO";
    defparam add_1112_35.INJECT1_1 = "NO";
    CCU2D add_1112_33 (.A0(d_d_tmp[66]), .B0(n6123), .C0(n6124[30]), .D0(d_tmp[66]), 
          .A1(d_d_tmp[67]), .B1(n6123), .C1(n6124[31]), .D1(d_tmp[67]), 
          .CIN(n11309), .COUT(n11310), .S0(d6_71__N_1459[66]), .S1(d6_71__N_1459[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1112_33.INIT0 = 16'hb874;
    defparam add_1112_33.INIT1 = 16'hb874;
    defparam add_1112_33.INJECT1_0 = "NO";
    defparam add_1112_33.INJECT1_1 = "NO";
    CCU2D add_1112_31 (.A0(d_d_tmp[64]), .B0(n6123), .C0(n6124[28]), .D0(d_tmp[64]), 
          .A1(d_d_tmp[65]), .B1(n6123), .C1(n6124[29]), .D1(d_tmp[65]), 
          .CIN(n11308), .COUT(n11309), .S0(d6_71__N_1459[64]), .S1(d6_71__N_1459[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1112_31.INIT0 = 16'hb874;
    defparam add_1112_31.INIT1 = 16'hb874;
    defparam add_1112_31.INJECT1_0 = "NO";
    defparam add_1112_31.INJECT1_1 = "NO";
    CCU2D add_1112_29 (.A0(d_d_tmp[62]), .B0(n6123), .C0(n6124[26]), .D0(d_tmp[62]), 
          .A1(d_d_tmp[63]), .B1(n6123), .C1(n6124[27]), .D1(d_tmp[63]), 
          .CIN(n11307), .COUT(n11308), .S0(d6_71__N_1459[62]), .S1(d6_71__N_1459[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1112_29.INIT0 = 16'hb874;
    defparam add_1112_29.INIT1 = 16'hb874;
    defparam add_1112_29.INJECT1_0 = "NO";
    defparam add_1112_29.INJECT1_1 = "NO";
    CCU2D add_1112_27 (.A0(d_d_tmp[60]), .B0(n6123), .C0(n6124[24]), .D0(d_tmp[60]), 
          .A1(d_d_tmp[61]), .B1(n6123), .C1(n6124[25]), .D1(d_tmp[61]), 
          .CIN(n11306), .COUT(n11307), .S0(d6_71__N_1459[60]), .S1(d6_71__N_1459[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1112_27.INIT0 = 16'hb874;
    defparam add_1112_27.INIT1 = 16'hb874;
    defparam add_1112_27.INJECT1_0 = "NO";
    defparam add_1112_27.INJECT1_1 = "NO";
    CCU2D add_1112_25 (.A0(d_d_tmp[58]), .B0(n6123), .C0(n6124[22]), .D0(d_tmp[58]), 
          .A1(d_d_tmp[59]), .B1(n6123), .C1(n6124[23]), .D1(d_tmp[59]), 
          .CIN(n11305), .COUT(n11306), .S0(d6_71__N_1459[58]), .S1(d6_71__N_1459[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1112_25.INIT0 = 16'hb874;
    defparam add_1112_25.INIT1 = 16'hb874;
    defparam add_1112_25.INJECT1_0 = "NO";
    defparam add_1112_25.INJECT1_1 = "NO";
    CCU2D add_1112_23 (.A0(d_d_tmp[56]), .B0(n6123), .C0(n6124[20]), .D0(d_tmp[56]), 
          .A1(d_d_tmp[57]), .B1(n6123), .C1(n6124[21]), .D1(d_tmp[57]), 
          .CIN(n11304), .COUT(n11305), .S0(d6_71__N_1459[56]), .S1(d6_71__N_1459[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1112_23.INIT0 = 16'hb874;
    defparam add_1112_23.INIT1 = 16'hb874;
    defparam add_1112_23.INJECT1_0 = "NO";
    defparam add_1112_23.INJECT1_1 = "NO";
    CCU2D add_1112_21 (.A0(d_d_tmp[54]), .B0(n6123), .C0(n6124[18]), .D0(d_tmp[54]), 
          .A1(d_d_tmp[55]), .B1(n6123), .C1(n6124[19]), .D1(d_tmp[55]), 
          .CIN(n11303), .COUT(n11304), .S0(d6_71__N_1459[54]), .S1(d6_71__N_1459[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1112_21.INIT0 = 16'hb874;
    defparam add_1112_21.INIT1 = 16'hb874;
    defparam add_1112_21.INJECT1_0 = "NO";
    defparam add_1112_21.INJECT1_1 = "NO";
    CCU2D add_1112_19 (.A0(d_d_tmp[52]), .B0(n6123), .C0(n6124[16]), .D0(d_tmp[52]), 
          .A1(d_d_tmp[53]), .B1(n6123), .C1(n6124[17]), .D1(d_tmp[53]), 
          .CIN(n11302), .COUT(n11303), .S0(d6_71__N_1459[52]), .S1(d6_71__N_1459[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1112_19.INIT0 = 16'hb874;
    defparam add_1112_19.INIT1 = 16'hb874;
    defparam add_1112_19.INJECT1_0 = "NO";
    defparam add_1112_19.INJECT1_1 = "NO";
    CCU2D add_1112_17 (.A0(d_d_tmp[50]), .B0(n6123), .C0(n6124[14]), .D0(d_tmp[50]), 
          .A1(d_d_tmp[51]), .B1(n6123), .C1(n6124[15]), .D1(d_tmp[51]), 
          .CIN(n11301), .COUT(n11302), .S0(d6_71__N_1459[50]), .S1(d6_71__N_1459[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1112_17.INIT0 = 16'hb874;
    defparam add_1112_17.INIT1 = 16'hb874;
    defparam add_1112_17.INJECT1_0 = "NO";
    defparam add_1112_17.INJECT1_1 = "NO";
    CCU2D add_1112_15 (.A0(d_d_tmp[48]), .B0(n6123), .C0(n6124[12]), .D0(d_tmp[48]), 
          .A1(d_d_tmp[49]), .B1(n6123), .C1(n6124[13]), .D1(d_tmp[49]), 
          .CIN(n11300), .COUT(n11301), .S0(d6_71__N_1459[48]), .S1(d6_71__N_1459[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1112_15.INIT0 = 16'hb874;
    defparam add_1112_15.INIT1 = 16'hb874;
    defparam add_1112_15.INJECT1_0 = "NO";
    defparam add_1112_15.INJECT1_1 = "NO";
    CCU2D add_1112_13 (.A0(d_d_tmp[46]), .B0(n6123), .C0(n6124[10]), .D0(d_tmp[46]), 
          .A1(d_d_tmp[47]), .B1(n6123), .C1(n6124[11]), .D1(d_tmp[47]), 
          .CIN(n11299), .COUT(n11300), .S0(d6_71__N_1459[46]), .S1(d6_71__N_1459[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1112_13.INIT0 = 16'hb874;
    defparam add_1112_13.INIT1 = 16'hb874;
    defparam add_1112_13.INJECT1_0 = "NO";
    defparam add_1112_13.INJECT1_1 = "NO";
    CCU2D add_1112_11 (.A0(d_d_tmp[44]), .B0(n6123), .C0(n6124[8]), .D0(d_tmp[44]), 
          .A1(d_d_tmp[45]), .B1(n6123), .C1(n6124[9]), .D1(d_tmp[45]), 
          .CIN(n11298), .COUT(n11299), .S0(d6_71__N_1459[44]), .S1(d6_71__N_1459[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1112_11.INIT0 = 16'hb874;
    defparam add_1112_11.INIT1 = 16'hb874;
    defparam add_1112_11.INJECT1_0 = "NO";
    defparam add_1112_11.INJECT1_1 = "NO";
    CCU2D add_1112_9 (.A0(d_d_tmp[42]), .B0(n6123), .C0(n6124[6]), .D0(d_tmp[42]), 
          .A1(d_d_tmp[43]), .B1(n6123), .C1(n6124[7]), .D1(d_tmp[43]), 
          .CIN(n11297), .COUT(n11298), .S0(d6_71__N_1459[42]), .S1(d6_71__N_1459[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1112_9.INIT0 = 16'hb874;
    defparam add_1112_9.INIT1 = 16'hb874;
    defparam add_1112_9.INJECT1_0 = "NO";
    defparam add_1112_9.INJECT1_1 = "NO";
    CCU2D add_1112_7 (.A0(d_d_tmp[40]), .B0(n6123), .C0(n6124[4]), .D0(d_tmp[40]), 
          .A1(d_d_tmp[41]), .B1(n6123), .C1(n6124[5]), .D1(d_tmp[41]), 
          .CIN(n11296), .COUT(n11297), .S0(d6_71__N_1459[40]), .S1(d6_71__N_1459[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1112_7.INIT0 = 16'hb874;
    defparam add_1112_7.INIT1 = 16'hb874;
    defparam add_1112_7.INJECT1_0 = "NO";
    defparam add_1112_7.INJECT1_1 = "NO";
    CCU2D add_1112_5 (.A0(d_d_tmp[38]), .B0(n6123), .C0(n6124[2]), .D0(d_tmp[38]), 
          .A1(d_d_tmp[39]), .B1(n6123), .C1(n6124[3]), .D1(d_tmp[39]), 
          .CIN(n11295), .COUT(n11296), .S0(d6_71__N_1459[38]), .S1(d6_71__N_1459[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1112_5.INIT0 = 16'hb874;
    defparam add_1112_5.INIT1 = 16'hb874;
    defparam add_1112_5.INJECT1_0 = "NO";
    defparam add_1112_5.INJECT1_1 = "NO";
    CCU2D add_1112_3 (.A0(d_d_tmp[36]), .B0(n6123), .C0(n6124[0]), .D0(d_tmp[36]), 
          .A1(d_d_tmp[37]), .B1(n6123), .C1(n6124[1]), .D1(d_tmp[37]), 
          .CIN(n11294), .COUT(n11295), .S0(d6_71__N_1459[36]), .S1(d6_71__N_1459[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1112_3.INIT0 = 16'hb874;
    defparam add_1112_3.INIT1 = 16'hb874;
    defparam add_1112_3.INJECT1_0 = "NO";
    defparam add_1112_3.INJECT1_1 = "NO";
    CCU2D add_1112_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n6123), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11294));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1112_1.INIT0 = 16'hF000;
    defparam add_1112_1.INIT1 = 16'h0555;
    defparam add_1112_1.INJECT1_0 = "NO";
    defparam add_1112_1.INJECT1_1 = "NO";
    CCU2D add_1116_37 (.A0(d6[71]), .B0(d_d6[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11290), 
          .S0(n6276[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1116_37.INIT0 = 16'h5999;
    defparam add_1116_37.INIT1 = 16'h0000;
    defparam add_1116_37.INJECT1_0 = "NO";
    defparam add_1116_37.INJECT1_1 = "NO";
    CCU2D add_1116_35 (.A0(d6[69]), .B0(d_d6[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[70]), .B1(d_d6[70]), .C1(GND_net), .D1(GND_net), .CIN(n11289), 
          .COUT(n11290), .S0(n6276[33]), .S1(n6276[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1116_35.INIT0 = 16'h5999;
    defparam add_1116_35.INIT1 = 16'h5999;
    defparam add_1116_35.INJECT1_0 = "NO";
    defparam add_1116_35.INJECT1_1 = "NO";
    CCU2D add_1116_33 (.A0(d6[67]), .B0(d_d6[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[68]), .B1(d_d6[68]), .C1(GND_net), .D1(GND_net), .CIN(n11288), 
          .COUT(n11289), .S0(n6276[31]), .S1(n6276[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1116_33.INIT0 = 16'h5999;
    defparam add_1116_33.INIT1 = 16'h5999;
    defparam add_1116_33.INJECT1_0 = "NO";
    defparam add_1116_33.INJECT1_1 = "NO";
    CCU2D add_1116_31 (.A0(d6[65]), .B0(d_d6[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[66]), .B1(d_d6[66]), .C1(GND_net), .D1(GND_net), .CIN(n11287), 
          .COUT(n11288), .S0(n6276[29]), .S1(n6276[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1116_31.INIT0 = 16'h5999;
    defparam add_1116_31.INIT1 = 16'h5999;
    defparam add_1116_31.INJECT1_0 = "NO";
    defparam add_1116_31.INJECT1_1 = "NO";
    CCU2D add_1116_29 (.A0(d6[63]), .B0(d_d6[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[64]), .B1(d_d6[64]), .C1(GND_net), .D1(GND_net), .CIN(n11286), 
          .COUT(n11287), .S0(n6276[27]), .S1(n6276[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1116_29.INIT0 = 16'h5999;
    defparam add_1116_29.INIT1 = 16'h5999;
    defparam add_1116_29.INJECT1_0 = "NO";
    defparam add_1116_29.INJECT1_1 = "NO";
    CCU2D add_1116_27 (.A0(d6[61]), .B0(d_d6[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[62]), .B1(d_d6[62]), .C1(GND_net), .D1(GND_net), .CIN(n11285), 
          .COUT(n11286), .S0(n6276[25]), .S1(n6276[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1116_27.INIT0 = 16'h5999;
    defparam add_1116_27.INIT1 = 16'h5999;
    defparam add_1116_27.INJECT1_0 = "NO";
    defparam add_1116_27.INJECT1_1 = "NO";
    CCU2D add_1116_25 (.A0(d6[59]), .B0(d_d6[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[60]), .B1(d_d6[60]), .C1(GND_net), .D1(GND_net), .CIN(n11284), 
          .COUT(n11285), .S0(n6276[23]), .S1(n6276[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1116_25.INIT0 = 16'h5999;
    defparam add_1116_25.INIT1 = 16'h5999;
    defparam add_1116_25.INJECT1_0 = "NO";
    defparam add_1116_25.INJECT1_1 = "NO";
    CCU2D add_1116_23 (.A0(d6[57]), .B0(d_d6[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[58]), .B1(d_d6[58]), .C1(GND_net), .D1(GND_net), .CIN(n11283), 
          .COUT(n11284), .S0(n6276[21]), .S1(n6276[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1116_23.INIT0 = 16'h5999;
    defparam add_1116_23.INIT1 = 16'h5999;
    defparam add_1116_23.INJECT1_0 = "NO";
    defparam add_1116_23.INJECT1_1 = "NO";
    CCU2D add_1116_21 (.A0(d6[55]), .B0(d_d6[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[56]), .B1(d_d6[56]), .C1(GND_net), .D1(GND_net), .CIN(n11282), 
          .COUT(n11283), .S0(n6276[19]), .S1(n6276[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1116_21.INIT0 = 16'h5999;
    defparam add_1116_21.INIT1 = 16'h5999;
    defparam add_1116_21.INJECT1_0 = "NO";
    defparam add_1116_21.INJECT1_1 = "NO";
    CCU2D add_1116_19 (.A0(d6[53]), .B0(d_d6[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[54]), .B1(d_d6[54]), .C1(GND_net), .D1(GND_net), .CIN(n11281), 
          .COUT(n11282), .S0(n6276[17]), .S1(n6276[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1116_19.INIT0 = 16'h5999;
    defparam add_1116_19.INIT1 = 16'h5999;
    defparam add_1116_19.INJECT1_0 = "NO";
    defparam add_1116_19.INJECT1_1 = "NO";
    CCU2D add_1116_17 (.A0(d6[51]), .B0(d_d6[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[52]), .B1(d_d6[52]), .C1(GND_net), .D1(GND_net), .CIN(n11280), 
          .COUT(n11281), .S0(n6276[15]), .S1(n6276[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1116_17.INIT0 = 16'h5999;
    defparam add_1116_17.INIT1 = 16'h5999;
    defparam add_1116_17.INJECT1_0 = "NO";
    defparam add_1116_17.INJECT1_1 = "NO";
    CCU2D add_1116_15 (.A0(d6[49]), .B0(d_d6[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[50]), .B1(d_d6[50]), .C1(GND_net), .D1(GND_net), .CIN(n11279), 
          .COUT(n11280), .S0(n6276[13]), .S1(n6276[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1116_15.INIT0 = 16'h5999;
    defparam add_1116_15.INIT1 = 16'h5999;
    defparam add_1116_15.INJECT1_0 = "NO";
    defparam add_1116_15.INJECT1_1 = "NO";
    CCU2D add_1116_13 (.A0(d6[47]), .B0(d_d6[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[48]), .B1(d_d6[48]), .C1(GND_net), .D1(GND_net), .CIN(n11278), 
          .COUT(n11279), .S0(n6276[11]), .S1(n6276[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1116_13.INIT0 = 16'h5999;
    defparam add_1116_13.INIT1 = 16'h5999;
    defparam add_1116_13.INJECT1_0 = "NO";
    defparam add_1116_13.INJECT1_1 = "NO";
    CCU2D add_1116_11 (.A0(d6[45]), .B0(d_d6[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[46]), .B1(d_d6[46]), .C1(GND_net), .D1(GND_net), .CIN(n11277), 
          .COUT(n11278), .S0(n6276[9]), .S1(n6276[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1116_11.INIT0 = 16'h5999;
    defparam add_1116_11.INIT1 = 16'h5999;
    defparam add_1116_11.INJECT1_0 = "NO";
    defparam add_1116_11.INJECT1_1 = "NO";
    CCU2D add_1116_9 (.A0(d6[43]), .B0(d_d6[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[44]), .B1(d_d6[44]), .C1(GND_net), .D1(GND_net), .CIN(n11276), 
          .COUT(n11277), .S0(n6276[7]), .S1(n6276[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1116_9.INIT0 = 16'h5999;
    defparam add_1116_9.INIT1 = 16'h5999;
    defparam add_1116_9.INJECT1_0 = "NO";
    defparam add_1116_9.INJECT1_1 = "NO";
    CCU2D add_1116_7 (.A0(d6[41]), .B0(d_d6[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[42]), .B1(d_d6[42]), .C1(GND_net), .D1(GND_net), .CIN(n11275), 
          .COUT(n11276), .S0(n6276[5]), .S1(n6276[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1116_7.INIT0 = 16'h5999;
    defparam add_1116_7.INIT1 = 16'h5999;
    defparam add_1116_7.INJECT1_0 = "NO";
    defparam add_1116_7.INJECT1_1 = "NO";
    CCU2D add_1116_5 (.A0(d6[39]), .B0(d_d6[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[40]), .B1(d_d6[40]), .C1(GND_net), .D1(GND_net), .CIN(n11274), 
          .COUT(n11275), .S0(n6276[3]), .S1(n6276[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1116_5.INIT0 = 16'h5999;
    defparam add_1116_5.INIT1 = 16'h5999;
    defparam add_1116_5.INJECT1_0 = "NO";
    defparam add_1116_5.INJECT1_1 = "NO";
    CCU2D add_1116_3 (.A0(d6[37]), .B0(d_d6[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[38]), .B1(d_d6[38]), .C1(GND_net), .D1(GND_net), .CIN(n11273), 
          .COUT(n11274), .S0(n6276[1]), .S1(n6276[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1116_3.INIT0 = 16'h5999;
    defparam add_1116_3.INIT1 = 16'h5999;
    defparam add_1116_3.INJECT1_0 = "NO";
    defparam add_1116_3.INJECT1_1 = "NO";
    CCU2D add_1116_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d6[36]), .B1(d_d6[36]), .C1(GND_net), .D1(GND_net), .COUT(n11273), 
          .S1(n6276[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1116_1.INIT0 = 16'hF000;
    defparam add_1116_1.INIT1 = 16'h5999;
    defparam add_1116_1.INJECT1_0 = "NO";
    defparam add_1116_1.INJECT1_1 = "NO";
    CCU2D add_1117_37 (.A0(d_d6[70]), .B0(n6275), .C0(n6276[34]), .D0(d6[70]), 
          .A1(d_d6[71]), .B1(n6275), .C1(n6276[35]), .D1(d6[71]), .CIN(n11271), 
          .S0(d7_71__N_1531[70]), .S1(d7_71__N_1531[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1117_37.INIT0 = 16'hb874;
    defparam add_1117_37.INIT1 = 16'hb874;
    defparam add_1117_37.INJECT1_0 = "NO";
    defparam add_1117_37.INJECT1_1 = "NO";
    CCU2D add_1117_35 (.A0(d_d6[68]), .B0(n6275), .C0(n6276[32]), .D0(d6[68]), 
          .A1(d_d6[69]), .B1(n6275), .C1(n6276[33]), .D1(d6[69]), .CIN(n11270), 
          .COUT(n11271), .S0(d7_71__N_1531[68]), .S1(d7_71__N_1531[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1117_35.INIT0 = 16'hb874;
    defparam add_1117_35.INIT1 = 16'hb874;
    defparam add_1117_35.INJECT1_0 = "NO";
    defparam add_1117_35.INJECT1_1 = "NO";
    CCU2D add_1117_33 (.A0(d_d6[66]), .B0(n6275), .C0(n6276[30]), .D0(d6[66]), 
          .A1(d_d6[67]), .B1(n6275), .C1(n6276[31]), .D1(d6[67]), .CIN(n11269), 
          .COUT(n11270), .S0(d7_71__N_1531[66]), .S1(d7_71__N_1531[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1117_33.INIT0 = 16'hb874;
    defparam add_1117_33.INIT1 = 16'hb874;
    defparam add_1117_33.INJECT1_0 = "NO";
    defparam add_1117_33.INJECT1_1 = "NO";
    CCU2D add_1117_31 (.A0(d_d6[64]), .B0(n6275), .C0(n6276[28]), .D0(d6[64]), 
          .A1(d_d6[65]), .B1(n6275), .C1(n6276[29]), .D1(d6[65]), .CIN(n11268), 
          .COUT(n11269), .S0(d7_71__N_1531[64]), .S1(d7_71__N_1531[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1117_31.INIT0 = 16'hb874;
    defparam add_1117_31.INIT1 = 16'hb874;
    defparam add_1117_31.INJECT1_0 = "NO";
    defparam add_1117_31.INJECT1_1 = "NO";
    CCU2D add_1117_29 (.A0(d_d6[62]), .B0(n6275), .C0(n6276[26]), .D0(d6[62]), 
          .A1(d_d6[63]), .B1(n6275), .C1(n6276[27]), .D1(d6[63]), .CIN(n11267), 
          .COUT(n11268), .S0(d7_71__N_1531[62]), .S1(d7_71__N_1531[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1117_29.INIT0 = 16'hb874;
    defparam add_1117_29.INIT1 = 16'hb874;
    defparam add_1117_29.INJECT1_0 = "NO";
    defparam add_1117_29.INJECT1_1 = "NO";
    CCU2D add_1117_27 (.A0(d_d6[60]), .B0(n6275), .C0(n6276[24]), .D0(d6[60]), 
          .A1(d_d6[61]), .B1(n6275), .C1(n6276[25]), .D1(d6[61]), .CIN(n11266), 
          .COUT(n11267), .S0(d7_71__N_1531[60]), .S1(d7_71__N_1531[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1117_27.INIT0 = 16'hb874;
    defparam add_1117_27.INIT1 = 16'hb874;
    defparam add_1117_27.INJECT1_0 = "NO";
    defparam add_1117_27.INJECT1_1 = "NO";
    CCU2D add_1117_25 (.A0(d_d6[58]), .B0(n6275), .C0(n6276[22]), .D0(d6[58]), 
          .A1(d_d6[59]), .B1(n6275), .C1(n6276[23]), .D1(d6[59]), .CIN(n11265), 
          .COUT(n11266), .S0(d7_71__N_1531[58]), .S1(d7_71__N_1531[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1117_25.INIT0 = 16'hb874;
    defparam add_1117_25.INIT1 = 16'hb874;
    defparam add_1117_25.INJECT1_0 = "NO";
    defparam add_1117_25.INJECT1_1 = "NO";
    CCU2D add_1117_23 (.A0(d_d6[56]), .B0(n6275), .C0(n6276[20]), .D0(d6[56]), 
          .A1(d_d6[57]), .B1(n6275), .C1(n6276[21]), .D1(d6[57]), .CIN(n11264), 
          .COUT(n11265), .S0(d7_71__N_1531[56]), .S1(d7_71__N_1531[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1117_23.INIT0 = 16'hb874;
    defparam add_1117_23.INIT1 = 16'hb874;
    defparam add_1117_23.INJECT1_0 = "NO";
    defparam add_1117_23.INJECT1_1 = "NO";
    CCU2D add_1117_21 (.A0(d_d6[54]), .B0(n6275), .C0(n6276[18]), .D0(d6[54]), 
          .A1(d_d6[55]), .B1(n6275), .C1(n6276[19]), .D1(d6[55]), .CIN(n11263), 
          .COUT(n11264), .S0(d7_71__N_1531[54]), .S1(d7_71__N_1531[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1117_21.INIT0 = 16'hb874;
    defparam add_1117_21.INIT1 = 16'hb874;
    defparam add_1117_21.INJECT1_0 = "NO";
    defparam add_1117_21.INJECT1_1 = "NO";
    CCU2D add_1117_19 (.A0(d_d6[52]), .B0(n6275), .C0(n6276[16]), .D0(d6[52]), 
          .A1(d_d6[53]), .B1(n6275), .C1(n6276[17]), .D1(d6[53]), .CIN(n11262), 
          .COUT(n11263), .S0(d7_71__N_1531[52]), .S1(d7_71__N_1531[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1117_19.INIT0 = 16'hb874;
    defparam add_1117_19.INIT1 = 16'hb874;
    defparam add_1117_19.INJECT1_0 = "NO";
    defparam add_1117_19.INJECT1_1 = "NO";
    CCU2D add_1117_17 (.A0(d_d6[50]), .B0(n6275), .C0(n6276[14]), .D0(d6[50]), 
          .A1(d_d6[51]), .B1(n6275), .C1(n6276[15]), .D1(d6[51]), .CIN(n11261), 
          .COUT(n11262), .S0(d7_71__N_1531[50]), .S1(d7_71__N_1531[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1117_17.INIT0 = 16'hb874;
    defparam add_1117_17.INIT1 = 16'hb874;
    defparam add_1117_17.INJECT1_0 = "NO";
    defparam add_1117_17.INJECT1_1 = "NO";
    CCU2D add_1117_15 (.A0(d_d6[48]), .B0(n6275), .C0(n6276[12]), .D0(d6[48]), 
          .A1(d_d6[49]), .B1(n6275), .C1(n6276[13]), .D1(d6[49]), .CIN(n11260), 
          .COUT(n11261), .S0(d7_71__N_1531[48]), .S1(d7_71__N_1531[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1117_15.INIT0 = 16'hb874;
    defparam add_1117_15.INIT1 = 16'hb874;
    defparam add_1117_15.INJECT1_0 = "NO";
    defparam add_1117_15.INJECT1_1 = "NO";
    CCU2D add_1117_13 (.A0(d_d6[46]), .B0(n6275), .C0(n6276[10]), .D0(d6[46]), 
          .A1(d_d6[47]), .B1(n6275), .C1(n6276[11]), .D1(d6[47]), .CIN(n11259), 
          .COUT(n11260), .S0(d7_71__N_1531[46]), .S1(d7_71__N_1531[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1117_13.INIT0 = 16'hb874;
    defparam add_1117_13.INIT1 = 16'hb874;
    defparam add_1117_13.INJECT1_0 = "NO";
    defparam add_1117_13.INJECT1_1 = "NO";
    CCU2D add_1117_11 (.A0(d_d6[44]), .B0(n6275), .C0(n6276[8]), .D0(d6[44]), 
          .A1(d_d6[45]), .B1(n6275), .C1(n6276[9]), .D1(d6[45]), .CIN(n11258), 
          .COUT(n11259), .S0(d7_71__N_1531[44]), .S1(d7_71__N_1531[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1117_11.INIT0 = 16'hb874;
    defparam add_1117_11.INIT1 = 16'hb874;
    defparam add_1117_11.INJECT1_0 = "NO";
    defparam add_1117_11.INJECT1_1 = "NO";
    CCU2D add_1117_9 (.A0(d_d6[42]), .B0(n6275), .C0(n6276[6]), .D0(d6[42]), 
          .A1(d_d6[43]), .B1(n6275), .C1(n6276[7]), .D1(d6[43]), .CIN(n11257), 
          .COUT(n11258), .S0(d7_71__N_1531[42]), .S1(d7_71__N_1531[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1117_9.INIT0 = 16'hb874;
    defparam add_1117_9.INIT1 = 16'hb874;
    defparam add_1117_9.INJECT1_0 = "NO";
    defparam add_1117_9.INJECT1_1 = "NO";
    CCU2D add_1117_7 (.A0(d_d6[40]), .B0(n6275), .C0(n6276[4]), .D0(d6[40]), 
          .A1(d_d6[41]), .B1(n6275), .C1(n6276[5]), .D1(d6[41]), .CIN(n11256), 
          .COUT(n11257), .S0(d7_71__N_1531[40]), .S1(d7_71__N_1531[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1117_7.INIT0 = 16'hb874;
    defparam add_1117_7.INIT1 = 16'hb874;
    defparam add_1117_7.INJECT1_0 = "NO";
    defparam add_1117_7.INJECT1_1 = "NO";
    CCU2D add_1117_5 (.A0(d_d6[38]), .B0(n6275), .C0(n6276[2]), .D0(d6[38]), 
          .A1(d_d6[39]), .B1(n6275), .C1(n6276[3]), .D1(d6[39]), .CIN(n11255), 
          .COUT(n11256), .S0(d7_71__N_1531[38]), .S1(d7_71__N_1531[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1117_5.INIT0 = 16'hb874;
    defparam add_1117_5.INIT1 = 16'hb874;
    defparam add_1117_5.INJECT1_0 = "NO";
    defparam add_1117_5.INJECT1_1 = "NO";
    CCU2D add_1117_3 (.A0(d_d6[36]), .B0(n6275), .C0(n6276[0]), .D0(d6[36]), 
          .A1(d_d6[37]), .B1(n6275), .C1(n6276[1]), .D1(d6[37]), .CIN(n11254), 
          .COUT(n11255), .S0(d7_71__N_1531[36]), .S1(d7_71__N_1531[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1117_3.INIT0 = 16'hb874;
    defparam add_1117_3.INIT1 = 16'hb874;
    defparam add_1117_3.INJECT1_0 = "NO";
    defparam add_1117_3.INJECT1_1 = "NO";
    CCU2D add_1117_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n6275), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11254));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1117_1.INIT0 = 16'hF000;
    defparam add_1117_1.INIT1 = 16'h0555;
    defparam add_1117_1.INJECT1_0 = "NO";
    defparam add_1117_1.INJECT1_1 = "NO";
    CCU2D add_1121_37 (.A0(d7[71]), .B0(d_d7[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11250), 
          .S0(n6428[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1121_37.INIT0 = 16'h5999;
    defparam add_1121_37.INIT1 = 16'h0000;
    defparam add_1121_37.INJECT1_0 = "NO";
    defparam add_1121_37.INJECT1_1 = "NO";
    CCU2D add_1121_35 (.A0(d7[69]), .B0(d_d7[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[70]), .B1(d_d7[70]), .C1(GND_net), .D1(GND_net), .CIN(n11249), 
          .COUT(n11250), .S0(n6428[33]), .S1(n6428[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1121_35.INIT0 = 16'h5999;
    defparam add_1121_35.INIT1 = 16'h5999;
    defparam add_1121_35.INJECT1_0 = "NO";
    defparam add_1121_35.INJECT1_1 = "NO";
    CCU2D add_1121_33 (.A0(d7[67]), .B0(d_d7[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[68]), .B1(d_d7[68]), .C1(GND_net), .D1(GND_net), .CIN(n11248), 
          .COUT(n11249), .S0(n6428[31]), .S1(n6428[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1121_33.INIT0 = 16'h5999;
    defparam add_1121_33.INIT1 = 16'h5999;
    defparam add_1121_33.INJECT1_0 = "NO";
    defparam add_1121_33.INJECT1_1 = "NO";
    CCU2D add_1121_31 (.A0(d7[65]), .B0(d_d7[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[66]), .B1(d_d7[66]), .C1(GND_net), .D1(GND_net), .CIN(n11247), 
          .COUT(n11248), .S0(n6428[29]), .S1(n6428[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1121_31.INIT0 = 16'h5999;
    defparam add_1121_31.INIT1 = 16'h5999;
    defparam add_1121_31.INJECT1_0 = "NO";
    defparam add_1121_31.INJECT1_1 = "NO";
    CCU2D add_1121_29 (.A0(d7[63]), .B0(d_d7[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[64]), .B1(d_d7[64]), .C1(GND_net), .D1(GND_net), .CIN(n11246), 
          .COUT(n11247), .S0(n6428[27]), .S1(n6428[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1121_29.INIT0 = 16'h5999;
    defparam add_1121_29.INIT1 = 16'h5999;
    defparam add_1121_29.INJECT1_0 = "NO";
    defparam add_1121_29.INJECT1_1 = "NO";
    CCU2D add_1121_27 (.A0(d7[61]), .B0(d_d7[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[62]), .B1(d_d7[62]), .C1(GND_net), .D1(GND_net), .CIN(n11245), 
          .COUT(n11246), .S0(n6428[25]), .S1(n6428[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1121_27.INIT0 = 16'h5999;
    defparam add_1121_27.INIT1 = 16'h5999;
    defparam add_1121_27.INJECT1_0 = "NO";
    defparam add_1121_27.INJECT1_1 = "NO";
    CCU2D add_1121_25 (.A0(d7[59]), .B0(d_d7[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[60]), .B1(d_d7[60]), .C1(GND_net), .D1(GND_net), .CIN(n11244), 
          .COUT(n11245), .S0(n6428[23]), .S1(n6428[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1121_25.INIT0 = 16'h5999;
    defparam add_1121_25.INIT1 = 16'h5999;
    defparam add_1121_25.INJECT1_0 = "NO";
    defparam add_1121_25.INJECT1_1 = "NO";
    CCU2D add_1121_23 (.A0(d7[57]), .B0(d_d7[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[58]), .B1(d_d7[58]), .C1(GND_net), .D1(GND_net), .CIN(n11243), 
          .COUT(n11244), .S0(n6428[21]), .S1(n6428[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1121_23.INIT0 = 16'h5999;
    defparam add_1121_23.INIT1 = 16'h5999;
    defparam add_1121_23.INJECT1_0 = "NO";
    defparam add_1121_23.INJECT1_1 = "NO";
    CCU2D add_1121_21 (.A0(d7[55]), .B0(d_d7[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[56]), .B1(d_d7[56]), .C1(GND_net), .D1(GND_net), .CIN(n11242), 
          .COUT(n11243), .S0(n6428[19]), .S1(n6428[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1121_21.INIT0 = 16'h5999;
    defparam add_1121_21.INIT1 = 16'h5999;
    defparam add_1121_21.INJECT1_0 = "NO";
    defparam add_1121_21.INJECT1_1 = "NO";
    CCU2D add_1121_19 (.A0(d7[53]), .B0(d_d7[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[54]), .B1(d_d7[54]), .C1(GND_net), .D1(GND_net), .CIN(n11241), 
          .COUT(n11242), .S0(n6428[17]), .S1(n6428[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1121_19.INIT0 = 16'h5999;
    defparam add_1121_19.INIT1 = 16'h5999;
    defparam add_1121_19.INJECT1_0 = "NO";
    defparam add_1121_19.INJECT1_1 = "NO";
    CCU2D add_1121_17 (.A0(d7[51]), .B0(d_d7[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[52]), .B1(d_d7[52]), .C1(GND_net), .D1(GND_net), .CIN(n11240), 
          .COUT(n11241), .S0(n6428[15]), .S1(n6428[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1121_17.INIT0 = 16'h5999;
    defparam add_1121_17.INIT1 = 16'h5999;
    defparam add_1121_17.INJECT1_0 = "NO";
    defparam add_1121_17.INJECT1_1 = "NO";
    CCU2D add_1121_15 (.A0(d7[49]), .B0(d_d7[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[50]), .B1(d_d7[50]), .C1(GND_net), .D1(GND_net), .CIN(n11239), 
          .COUT(n11240), .S0(n6428[13]), .S1(n6428[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1121_15.INIT0 = 16'h5999;
    defparam add_1121_15.INIT1 = 16'h5999;
    defparam add_1121_15.INJECT1_0 = "NO";
    defparam add_1121_15.INJECT1_1 = "NO";
    CCU2D add_1121_13 (.A0(d7[47]), .B0(d_d7[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[48]), .B1(d_d7[48]), .C1(GND_net), .D1(GND_net), .CIN(n11238), 
          .COUT(n11239), .S0(n6428[11]), .S1(n6428[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1121_13.INIT0 = 16'h5999;
    defparam add_1121_13.INIT1 = 16'h5999;
    defparam add_1121_13.INJECT1_0 = "NO";
    defparam add_1121_13.INJECT1_1 = "NO";
    CCU2D add_1121_11 (.A0(d7[45]), .B0(d_d7[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[46]), .B1(d_d7[46]), .C1(GND_net), .D1(GND_net), .CIN(n11237), 
          .COUT(n11238), .S0(n6428[9]), .S1(n6428[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1121_11.INIT0 = 16'h5999;
    defparam add_1121_11.INIT1 = 16'h5999;
    defparam add_1121_11.INJECT1_0 = "NO";
    defparam add_1121_11.INJECT1_1 = "NO";
    CCU2D add_1121_9 (.A0(d7[43]), .B0(d_d7[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[44]), .B1(d_d7[44]), .C1(GND_net), .D1(GND_net), .CIN(n11236), 
          .COUT(n11237), .S0(n6428[7]), .S1(n6428[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1121_9.INIT0 = 16'h5999;
    defparam add_1121_9.INIT1 = 16'h5999;
    defparam add_1121_9.INJECT1_0 = "NO";
    defparam add_1121_9.INJECT1_1 = "NO";
    CCU2D add_1121_7 (.A0(d7[41]), .B0(d_d7[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[42]), .B1(d_d7[42]), .C1(GND_net), .D1(GND_net), .CIN(n11235), 
          .COUT(n11236), .S0(n6428[5]), .S1(n6428[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1121_7.INIT0 = 16'h5999;
    defparam add_1121_7.INIT1 = 16'h5999;
    defparam add_1121_7.INJECT1_0 = "NO";
    defparam add_1121_7.INJECT1_1 = "NO";
    CCU2D add_1121_5 (.A0(d7[39]), .B0(d_d7[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[40]), .B1(d_d7[40]), .C1(GND_net), .D1(GND_net), .CIN(n11234), 
          .COUT(n11235), .S0(n6428[3]), .S1(n6428[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1121_5.INIT0 = 16'h5999;
    defparam add_1121_5.INIT1 = 16'h5999;
    defparam add_1121_5.INJECT1_0 = "NO";
    defparam add_1121_5.INJECT1_1 = "NO";
    CCU2D add_1121_3 (.A0(d7[37]), .B0(d_d7[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[38]), .B1(d_d7[38]), .C1(GND_net), .D1(GND_net), .CIN(n11233), 
          .COUT(n11234), .S0(n6428[1]), .S1(n6428[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1121_3.INIT0 = 16'h5999;
    defparam add_1121_3.INIT1 = 16'h5999;
    defparam add_1121_3.INJECT1_0 = "NO";
    defparam add_1121_3.INJECT1_1 = "NO";
    CCU2D add_1121_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d7[36]), .B1(d_d7[36]), .C1(GND_net), .D1(GND_net), .COUT(n11233), 
          .S1(n6428[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1121_1.INIT0 = 16'hF000;
    defparam add_1121_1.INIT1 = 16'h5999;
    defparam add_1121_1.INJECT1_0 = "NO";
    defparam add_1121_1.INJECT1_1 = "NO";
    CCU2D add_1122_37 (.A0(d_d7[70]), .B0(n6427), .C0(n6428[34]), .D0(d7[70]), 
          .A1(d_d7[71]), .B1(n6427), .C1(n6428[35]), .D1(d7[71]), .CIN(n11231), 
          .S0(d8_71__N_1603[70]), .S1(d8_71__N_1603[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1122_37.INIT0 = 16'hb874;
    defparam add_1122_37.INIT1 = 16'hb874;
    defparam add_1122_37.INJECT1_0 = "NO";
    defparam add_1122_37.INJECT1_1 = "NO";
    CCU2D add_1122_35 (.A0(d_d7[68]), .B0(n6427), .C0(n6428[32]), .D0(d7[68]), 
          .A1(d_d7[69]), .B1(n6427), .C1(n6428[33]), .D1(d7[69]), .CIN(n11230), 
          .COUT(n11231), .S0(d8_71__N_1603[68]), .S1(d8_71__N_1603[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1122_35.INIT0 = 16'hb874;
    defparam add_1122_35.INIT1 = 16'hb874;
    defparam add_1122_35.INJECT1_0 = "NO";
    defparam add_1122_35.INJECT1_1 = "NO";
    CCU2D add_1122_33 (.A0(d_d7[66]), .B0(n6427), .C0(n6428[30]), .D0(d7[66]), 
          .A1(d_d7[67]), .B1(n6427), .C1(n6428[31]), .D1(d7[67]), .CIN(n11229), 
          .COUT(n11230), .S0(d8_71__N_1603[66]), .S1(d8_71__N_1603[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1122_33.INIT0 = 16'hb874;
    defparam add_1122_33.INIT1 = 16'hb874;
    defparam add_1122_33.INJECT1_0 = "NO";
    defparam add_1122_33.INJECT1_1 = "NO";
    CCU2D add_1122_31 (.A0(d_d7[64]), .B0(n6427), .C0(n6428[28]), .D0(d7[64]), 
          .A1(d_d7[65]), .B1(n6427), .C1(n6428[29]), .D1(d7[65]), .CIN(n11228), 
          .COUT(n11229), .S0(d8_71__N_1603[64]), .S1(d8_71__N_1603[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1122_31.INIT0 = 16'hb874;
    defparam add_1122_31.INIT1 = 16'hb874;
    defparam add_1122_31.INJECT1_0 = "NO";
    defparam add_1122_31.INJECT1_1 = "NO";
    CCU2D add_1122_29 (.A0(d_d7[62]), .B0(n6427), .C0(n6428[26]), .D0(d7[62]), 
          .A1(d_d7[63]), .B1(n6427), .C1(n6428[27]), .D1(d7[63]), .CIN(n11227), 
          .COUT(n11228), .S0(d8_71__N_1603[62]), .S1(d8_71__N_1603[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1122_29.INIT0 = 16'hb874;
    defparam add_1122_29.INIT1 = 16'hb874;
    defparam add_1122_29.INJECT1_0 = "NO";
    defparam add_1122_29.INJECT1_1 = "NO";
    CCU2D add_1122_27 (.A0(d_d7[60]), .B0(n6427), .C0(n6428[24]), .D0(d7[60]), 
          .A1(d_d7[61]), .B1(n6427), .C1(n6428[25]), .D1(d7[61]), .CIN(n11226), 
          .COUT(n11227), .S0(d8_71__N_1603[60]), .S1(d8_71__N_1603[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1122_27.INIT0 = 16'hb874;
    defparam add_1122_27.INIT1 = 16'hb874;
    defparam add_1122_27.INJECT1_0 = "NO";
    defparam add_1122_27.INJECT1_1 = "NO";
    CCU2D add_1122_25 (.A0(d_d7[58]), .B0(n6427), .C0(n6428[22]), .D0(d7[58]), 
          .A1(d_d7[59]), .B1(n6427), .C1(n6428[23]), .D1(d7[59]), .CIN(n11225), 
          .COUT(n11226), .S0(d8_71__N_1603[58]), .S1(d8_71__N_1603[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1122_25.INIT0 = 16'hb874;
    defparam add_1122_25.INIT1 = 16'hb874;
    defparam add_1122_25.INJECT1_0 = "NO";
    defparam add_1122_25.INJECT1_1 = "NO";
    CCU2D add_1122_23 (.A0(d_d7[56]), .B0(n6427), .C0(n6428[20]), .D0(d7[56]), 
          .A1(d_d7[57]), .B1(n6427), .C1(n6428[21]), .D1(d7[57]), .CIN(n11224), 
          .COUT(n11225), .S0(d8_71__N_1603[56]), .S1(d8_71__N_1603[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1122_23.INIT0 = 16'hb874;
    defparam add_1122_23.INIT1 = 16'hb874;
    defparam add_1122_23.INJECT1_0 = "NO";
    defparam add_1122_23.INJECT1_1 = "NO";
    CCU2D add_1122_21 (.A0(d_d7[54]), .B0(n6427), .C0(n6428[18]), .D0(d7[54]), 
          .A1(d_d7[55]), .B1(n6427), .C1(n6428[19]), .D1(d7[55]), .CIN(n11223), 
          .COUT(n11224), .S0(d8_71__N_1603[54]), .S1(d8_71__N_1603[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1122_21.INIT0 = 16'hb874;
    defparam add_1122_21.INIT1 = 16'hb874;
    defparam add_1122_21.INJECT1_0 = "NO";
    defparam add_1122_21.INJECT1_1 = "NO";
    CCU2D add_1122_19 (.A0(d_d7[52]), .B0(n6427), .C0(n6428[16]), .D0(d7[52]), 
          .A1(d_d7[53]), .B1(n6427), .C1(n6428[17]), .D1(d7[53]), .CIN(n11222), 
          .COUT(n11223), .S0(d8_71__N_1603[52]), .S1(d8_71__N_1603[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1122_19.INIT0 = 16'hb874;
    defparam add_1122_19.INIT1 = 16'hb874;
    defparam add_1122_19.INJECT1_0 = "NO";
    defparam add_1122_19.INJECT1_1 = "NO";
    CCU2D add_1122_17 (.A0(d_d7[50]), .B0(n6427), .C0(n6428[14]), .D0(d7[50]), 
          .A1(d_d7[51]), .B1(n6427), .C1(n6428[15]), .D1(d7[51]), .CIN(n11221), 
          .COUT(n11222), .S0(d8_71__N_1603[50]), .S1(d8_71__N_1603[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1122_17.INIT0 = 16'hb874;
    defparam add_1122_17.INIT1 = 16'hb874;
    defparam add_1122_17.INJECT1_0 = "NO";
    defparam add_1122_17.INJECT1_1 = "NO";
    CCU2D add_1122_15 (.A0(d_d7[48]), .B0(n6427), .C0(n6428[12]), .D0(d7[48]), 
          .A1(d_d7[49]), .B1(n6427), .C1(n6428[13]), .D1(d7[49]), .CIN(n11220), 
          .COUT(n11221), .S0(d8_71__N_1603[48]), .S1(d8_71__N_1603[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1122_15.INIT0 = 16'hb874;
    defparam add_1122_15.INIT1 = 16'hb874;
    defparam add_1122_15.INJECT1_0 = "NO";
    defparam add_1122_15.INJECT1_1 = "NO";
    CCU2D add_1122_13 (.A0(d_d7[46]), .B0(n6427), .C0(n6428[10]), .D0(d7[46]), 
          .A1(d_d7[47]), .B1(n6427), .C1(n6428[11]), .D1(d7[47]), .CIN(n11219), 
          .COUT(n11220), .S0(d8_71__N_1603[46]), .S1(d8_71__N_1603[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1122_13.INIT0 = 16'hb874;
    defparam add_1122_13.INIT1 = 16'hb874;
    defparam add_1122_13.INJECT1_0 = "NO";
    defparam add_1122_13.INJECT1_1 = "NO";
    CCU2D add_1122_11 (.A0(d_d7[44]), .B0(n6427), .C0(n6428[8]), .D0(d7[44]), 
          .A1(d_d7[45]), .B1(n6427), .C1(n6428[9]), .D1(d7[45]), .CIN(n11218), 
          .COUT(n11219), .S0(d8_71__N_1603[44]), .S1(d8_71__N_1603[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1122_11.INIT0 = 16'hb874;
    defparam add_1122_11.INIT1 = 16'hb874;
    defparam add_1122_11.INJECT1_0 = "NO";
    defparam add_1122_11.INJECT1_1 = "NO";
    CCU2D add_1122_9 (.A0(d_d7[42]), .B0(n6427), .C0(n6428[6]), .D0(d7[42]), 
          .A1(d_d7[43]), .B1(n6427), .C1(n6428[7]), .D1(d7[43]), .CIN(n11217), 
          .COUT(n11218), .S0(d8_71__N_1603[42]), .S1(d8_71__N_1603[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1122_9.INIT0 = 16'hb874;
    defparam add_1122_9.INIT1 = 16'hb874;
    defparam add_1122_9.INJECT1_0 = "NO";
    defparam add_1122_9.INJECT1_1 = "NO";
    CCU2D add_1122_7 (.A0(d_d7[40]), .B0(n6427), .C0(n6428[4]), .D0(d7[40]), 
          .A1(d_d7[41]), .B1(n6427), .C1(n6428[5]), .D1(d7[41]), .CIN(n11216), 
          .COUT(n11217), .S0(d8_71__N_1603[40]), .S1(d8_71__N_1603[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1122_7.INIT0 = 16'hb874;
    defparam add_1122_7.INIT1 = 16'hb874;
    defparam add_1122_7.INJECT1_0 = "NO";
    defparam add_1122_7.INJECT1_1 = "NO";
    CCU2D add_1122_5 (.A0(d_d7[38]), .B0(n6427), .C0(n6428[2]), .D0(d7[38]), 
          .A1(d_d7[39]), .B1(n6427), .C1(n6428[3]), .D1(d7[39]), .CIN(n11215), 
          .COUT(n11216), .S0(d8_71__N_1603[38]), .S1(d8_71__N_1603[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1122_5.INIT0 = 16'hb874;
    defparam add_1122_5.INIT1 = 16'hb874;
    defparam add_1122_5.INJECT1_0 = "NO";
    defparam add_1122_5.INJECT1_1 = "NO";
    CCU2D add_1122_3 (.A0(d_d7[36]), .B0(n6427), .C0(n6428[0]), .D0(d7[36]), 
          .A1(d_d7[37]), .B1(n6427), .C1(n6428[1]), .D1(d7[37]), .CIN(n11214), 
          .COUT(n11215), .S0(d8_71__N_1603[36]), .S1(d8_71__N_1603[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1122_3.INIT0 = 16'hb874;
    defparam add_1122_3.INIT1 = 16'hb874;
    defparam add_1122_3.INJECT1_0 = "NO";
    defparam add_1122_3.INJECT1_1 = "NO";
    CCU2D add_1122_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n6427), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11214));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1122_1.INIT0 = 16'hF000;
    defparam add_1122_1.INIT1 = 16'h0555;
    defparam add_1122_1.INJECT1_0 = "NO";
    defparam add_1122_1.INJECT1_1 = "NO";
    CCU2D add_1126_37 (.A0(d8[71]), .B0(d_d8[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11210), 
          .S0(n6580[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1126_37.INIT0 = 16'h5999;
    defparam add_1126_37.INIT1 = 16'h0000;
    defparam add_1126_37.INJECT1_0 = "NO";
    defparam add_1126_37.INJECT1_1 = "NO";
    CCU2D add_1126_35 (.A0(d8[69]), .B0(d_d8[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[70]), .B1(d_d8[70]), .C1(GND_net), .D1(GND_net), .CIN(n11209), 
          .COUT(n11210), .S0(n6580[33]), .S1(n6580[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1126_35.INIT0 = 16'h5999;
    defparam add_1126_35.INIT1 = 16'h5999;
    defparam add_1126_35.INJECT1_0 = "NO";
    defparam add_1126_35.INJECT1_1 = "NO";
    CCU2D add_1126_33 (.A0(d8[67]), .B0(d_d8[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[68]), .B1(d_d8[68]), .C1(GND_net), .D1(GND_net), .CIN(n11208), 
          .COUT(n11209), .S0(n6580[31]), .S1(n6580[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1126_33.INIT0 = 16'h5999;
    defparam add_1126_33.INIT1 = 16'h5999;
    defparam add_1126_33.INJECT1_0 = "NO";
    defparam add_1126_33.INJECT1_1 = "NO";
    CCU2D add_1126_31 (.A0(d8[65]), .B0(d_d8[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[66]), .B1(d_d8[66]), .C1(GND_net), .D1(GND_net), .CIN(n11207), 
          .COUT(n11208), .S0(n6580[29]), .S1(n6580[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1126_31.INIT0 = 16'h5999;
    defparam add_1126_31.INIT1 = 16'h5999;
    defparam add_1126_31.INJECT1_0 = "NO";
    defparam add_1126_31.INJECT1_1 = "NO";
    CCU2D add_1126_29 (.A0(d8[63]), .B0(d_d8[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[64]), .B1(d_d8[64]), .C1(GND_net), .D1(GND_net), .CIN(n11206), 
          .COUT(n11207), .S0(n6580[27]), .S1(n6580[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1126_29.INIT0 = 16'h5999;
    defparam add_1126_29.INIT1 = 16'h5999;
    defparam add_1126_29.INJECT1_0 = "NO";
    defparam add_1126_29.INJECT1_1 = "NO";
    CCU2D add_1126_27 (.A0(d8[61]), .B0(d_d8[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[62]), .B1(d_d8[62]), .C1(GND_net), .D1(GND_net), .CIN(n11205), 
          .COUT(n11206), .S0(n6580[25]), .S1(n6580[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1126_27.INIT0 = 16'h5999;
    defparam add_1126_27.INIT1 = 16'h5999;
    defparam add_1126_27.INJECT1_0 = "NO";
    defparam add_1126_27.INJECT1_1 = "NO";
    CCU2D add_1126_25 (.A0(d8[59]), .B0(d_d8[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[60]), .B1(d_d8[60]), .C1(GND_net), .D1(GND_net), .CIN(n11204), 
          .COUT(n11205), .S0(n6580[23]), .S1(n6580[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1126_25.INIT0 = 16'h5999;
    defparam add_1126_25.INIT1 = 16'h5999;
    defparam add_1126_25.INJECT1_0 = "NO";
    defparam add_1126_25.INJECT1_1 = "NO";
    CCU2D add_1126_23 (.A0(d8[57]), .B0(d_d8[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[58]), .B1(d_d8[58]), .C1(GND_net), .D1(GND_net), .CIN(n11203), 
          .COUT(n11204), .S0(n6580[21]), .S1(n6580[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1126_23.INIT0 = 16'h5999;
    defparam add_1126_23.INIT1 = 16'h5999;
    defparam add_1126_23.INJECT1_0 = "NO";
    defparam add_1126_23.INJECT1_1 = "NO";
    CCU2D add_1126_21 (.A0(d8[55]), .B0(d_d8[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[56]), .B1(d_d8[56]), .C1(GND_net), .D1(GND_net), .CIN(n11202), 
          .COUT(n11203), .S0(n6580[19]), .S1(n6580[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1126_21.INIT0 = 16'h5999;
    defparam add_1126_21.INIT1 = 16'h5999;
    defparam add_1126_21.INJECT1_0 = "NO";
    defparam add_1126_21.INJECT1_1 = "NO";
    CCU2D add_1126_19 (.A0(d8[53]), .B0(d_d8[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[54]), .B1(d_d8[54]), .C1(GND_net), .D1(GND_net), .CIN(n11201), 
          .COUT(n11202), .S0(n6580[17]), .S1(n6580[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1126_19.INIT0 = 16'h5999;
    defparam add_1126_19.INIT1 = 16'h5999;
    defparam add_1126_19.INJECT1_0 = "NO";
    defparam add_1126_19.INJECT1_1 = "NO";
    CCU2D add_1126_17 (.A0(d8[51]), .B0(d_d8[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[52]), .B1(d_d8[52]), .C1(GND_net), .D1(GND_net), .CIN(n11200), 
          .COUT(n11201), .S0(n6580[15]), .S1(n6580[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1126_17.INIT0 = 16'h5999;
    defparam add_1126_17.INIT1 = 16'h5999;
    defparam add_1126_17.INJECT1_0 = "NO";
    defparam add_1126_17.INJECT1_1 = "NO";
    CCU2D add_1126_15 (.A0(d8[49]), .B0(d_d8[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[50]), .B1(d_d8[50]), .C1(GND_net), .D1(GND_net), .CIN(n11199), 
          .COUT(n11200), .S0(n6580[13]), .S1(n6580[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1126_15.INIT0 = 16'h5999;
    defparam add_1126_15.INIT1 = 16'h5999;
    defparam add_1126_15.INJECT1_0 = "NO";
    defparam add_1126_15.INJECT1_1 = "NO";
    CCU2D add_1126_13 (.A0(d8[47]), .B0(d_d8[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[48]), .B1(d_d8[48]), .C1(GND_net), .D1(GND_net), .CIN(n11198), 
          .COUT(n11199), .S0(n6580[11]), .S1(n6580[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1126_13.INIT0 = 16'h5999;
    defparam add_1126_13.INIT1 = 16'h5999;
    defparam add_1126_13.INJECT1_0 = "NO";
    defparam add_1126_13.INJECT1_1 = "NO";
    CCU2D add_1126_11 (.A0(d8[45]), .B0(d_d8[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[46]), .B1(d_d8[46]), .C1(GND_net), .D1(GND_net), .CIN(n11197), 
          .COUT(n11198), .S0(n6580[9]), .S1(n6580[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1126_11.INIT0 = 16'h5999;
    defparam add_1126_11.INIT1 = 16'h5999;
    defparam add_1126_11.INJECT1_0 = "NO";
    defparam add_1126_11.INJECT1_1 = "NO";
    CCU2D add_1126_9 (.A0(d8[43]), .B0(d_d8[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[44]), .B1(d_d8[44]), .C1(GND_net), .D1(GND_net), .CIN(n11196), 
          .COUT(n11197), .S0(n6580[7]), .S1(n6580[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1126_9.INIT0 = 16'h5999;
    defparam add_1126_9.INIT1 = 16'h5999;
    defparam add_1126_9.INJECT1_0 = "NO";
    defparam add_1126_9.INJECT1_1 = "NO";
    CCU2D add_1126_7 (.A0(d8[41]), .B0(d_d8[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[42]), .B1(d_d8[42]), .C1(GND_net), .D1(GND_net), .CIN(n11195), 
          .COUT(n11196), .S0(n6580[5]), .S1(n6580[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1126_7.INIT0 = 16'h5999;
    defparam add_1126_7.INIT1 = 16'h5999;
    defparam add_1126_7.INJECT1_0 = "NO";
    defparam add_1126_7.INJECT1_1 = "NO";
    CCU2D add_1126_5 (.A0(d8[39]), .B0(d_d8[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[40]), .B1(d_d8[40]), .C1(GND_net), .D1(GND_net), .CIN(n11194), 
          .COUT(n11195), .S0(n6580[3]), .S1(n6580[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1126_5.INIT0 = 16'h5999;
    defparam add_1126_5.INIT1 = 16'h5999;
    defparam add_1126_5.INJECT1_0 = "NO";
    defparam add_1126_5.INJECT1_1 = "NO";
    CCU2D add_1126_3 (.A0(d8[37]), .B0(d_d8[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[38]), .B1(d_d8[38]), .C1(GND_net), .D1(GND_net), .CIN(n11193), 
          .COUT(n11194), .S0(n6580[1]), .S1(n6580[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1126_3.INIT0 = 16'h5999;
    defparam add_1126_3.INIT1 = 16'h5999;
    defparam add_1126_3.INJECT1_0 = "NO";
    defparam add_1126_3.INJECT1_1 = "NO";
    CCU2D add_1126_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d8[36]), .B1(d_d8[36]), .C1(GND_net), .D1(GND_net), .COUT(n11193), 
          .S1(n6580[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1126_1.INIT0 = 16'hF000;
    defparam add_1126_1.INIT1 = 16'h5999;
    defparam add_1126_1.INJECT1_0 = "NO";
    defparam add_1126_1.INJECT1_1 = "NO";
    CCU2D add_1127_37 (.A0(d_d8[70]), .B0(n6579), .C0(n6580[34]), .D0(d8[70]), 
          .A1(d_d8[71]), .B1(n6579), .C1(n6580[35]), .D1(d8[71]), .CIN(n11191), 
          .S0(d9_71__N_1675[70]), .S1(d9_71__N_1675[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1127_37.INIT0 = 16'hb874;
    defparam add_1127_37.INIT1 = 16'hb874;
    defparam add_1127_37.INJECT1_0 = "NO";
    defparam add_1127_37.INJECT1_1 = "NO";
    CCU2D add_1127_35 (.A0(d_d8[68]), .B0(n6579), .C0(n6580[32]), .D0(d8[68]), 
          .A1(d_d8[69]), .B1(n6579), .C1(n6580[33]), .D1(d8[69]), .CIN(n11190), 
          .COUT(n11191), .S0(d9_71__N_1675[68]), .S1(d9_71__N_1675[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1127_35.INIT0 = 16'hb874;
    defparam add_1127_35.INIT1 = 16'hb874;
    defparam add_1127_35.INJECT1_0 = "NO";
    defparam add_1127_35.INJECT1_1 = "NO";
    CCU2D add_1127_33 (.A0(d_d8[66]), .B0(n6579), .C0(n6580[30]), .D0(d8[66]), 
          .A1(d_d8[67]), .B1(n6579), .C1(n6580[31]), .D1(d8[67]), .CIN(n11189), 
          .COUT(n11190), .S0(d9_71__N_1675[66]), .S1(d9_71__N_1675[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1127_33.INIT0 = 16'hb874;
    defparam add_1127_33.INIT1 = 16'hb874;
    defparam add_1127_33.INJECT1_0 = "NO";
    defparam add_1127_33.INJECT1_1 = "NO";
    CCU2D add_1127_31 (.A0(d_d8[64]), .B0(n6579), .C0(n6580[28]), .D0(d8[64]), 
          .A1(d_d8[65]), .B1(n6579), .C1(n6580[29]), .D1(d8[65]), .CIN(n11188), 
          .COUT(n11189), .S0(d9_71__N_1675[64]), .S1(d9_71__N_1675[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1127_31.INIT0 = 16'hb874;
    defparam add_1127_31.INIT1 = 16'hb874;
    defparam add_1127_31.INJECT1_0 = "NO";
    defparam add_1127_31.INJECT1_1 = "NO";
    CCU2D add_1127_29 (.A0(d_d8[62]), .B0(n6579), .C0(n6580[26]), .D0(d8[62]), 
          .A1(d_d8[63]), .B1(n6579), .C1(n6580[27]), .D1(d8[63]), .CIN(n11187), 
          .COUT(n11188), .S0(d9_71__N_1675[62]), .S1(d9_71__N_1675[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1127_29.INIT0 = 16'hb874;
    defparam add_1127_29.INIT1 = 16'hb874;
    defparam add_1127_29.INJECT1_0 = "NO";
    defparam add_1127_29.INJECT1_1 = "NO";
    CCU2D add_1127_27 (.A0(d_d8[60]), .B0(n6579), .C0(n6580[24]), .D0(d8[60]), 
          .A1(d_d8[61]), .B1(n6579), .C1(n6580[25]), .D1(d8[61]), .CIN(n11186), 
          .COUT(n11187), .S0(d9_71__N_1675[60]), .S1(d9_71__N_1675[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1127_27.INIT0 = 16'hb874;
    defparam add_1127_27.INIT1 = 16'hb874;
    defparam add_1127_27.INJECT1_0 = "NO";
    defparam add_1127_27.INJECT1_1 = "NO";
    CCU2D add_1127_25 (.A0(d_d8[58]), .B0(n6579), .C0(n6580[22]), .D0(d8[58]), 
          .A1(d_d8[59]), .B1(n6579), .C1(n6580[23]), .D1(d8[59]), .CIN(n11185), 
          .COUT(n11186), .S0(d9_71__N_1675[58]), .S1(d9_71__N_1675[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1127_25.INIT0 = 16'hb874;
    defparam add_1127_25.INIT1 = 16'hb874;
    defparam add_1127_25.INJECT1_0 = "NO";
    defparam add_1127_25.INJECT1_1 = "NO";
    CCU2D add_1127_23 (.A0(d_d8[56]), .B0(n6579), .C0(n6580[20]), .D0(d8[56]), 
          .A1(d_d8[57]), .B1(n6579), .C1(n6580[21]), .D1(d8[57]), .CIN(n11184), 
          .COUT(n11185), .S0(d9_71__N_1675[56]), .S1(d9_71__N_1675[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1127_23.INIT0 = 16'hb874;
    defparam add_1127_23.INIT1 = 16'hb874;
    defparam add_1127_23.INJECT1_0 = "NO";
    defparam add_1127_23.INJECT1_1 = "NO";
    CCU2D add_1127_21 (.A0(d_d8[54]), .B0(n6579), .C0(n6580[18]), .D0(d8[54]), 
          .A1(d_d8[55]), .B1(n6579), .C1(n6580[19]), .D1(d8[55]), .CIN(n11183), 
          .COUT(n11184), .S0(d9_71__N_1675[54]), .S1(d9_71__N_1675[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1127_21.INIT0 = 16'hb874;
    defparam add_1127_21.INIT1 = 16'hb874;
    defparam add_1127_21.INJECT1_0 = "NO";
    defparam add_1127_21.INJECT1_1 = "NO";
    CCU2D add_1127_19 (.A0(d_d8[52]), .B0(n6579), .C0(n6580[16]), .D0(d8[52]), 
          .A1(d_d8[53]), .B1(n6579), .C1(n6580[17]), .D1(d8[53]), .CIN(n11182), 
          .COUT(n11183), .S0(d9_71__N_1675[52]), .S1(d9_71__N_1675[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1127_19.INIT0 = 16'hb874;
    defparam add_1127_19.INIT1 = 16'hb874;
    defparam add_1127_19.INJECT1_0 = "NO";
    defparam add_1127_19.INJECT1_1 = "NO";
    CCU2D add_1127_17 (.A0(d_d8[50]), .B0(n6579), .C0(n6580[14]), .D0(d8[50]), 
          .A1(d_d8[51]), .B1(n6579), .C1(n6580[15]), .D1(d8[51]), .CIN(n11181), 
          .COUT(n11182), .S0(d9_71__N_1675[50]), .S1(d9_71__N_1675[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1127_17.INIT0 = 16'hb874;
    defparam add_1127_17.INIT1 = 16'hb874;
    defparam add_1127_17.INJECT1_0 = "NO";
    defparam add_1127_17.INJECT1_1 = "NO";
    CCU2D add_1127_15 (.A0(d_d8[48]), .B0(n6579), .C0(n6580[12]), .D0(d8[48]), 
          .A1(d_d8[49]), .B1(n6579), .C1(n6580[13]), .D1(d8[49]), .CIN(n11180), 
          .COUT(n11181), .S0(d9_71__N_1675[48]), .S1(d9_71__N_1675[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1127_15.INIT0 = 16'hb874;
    defparam add_1127_15.INIT1 = 16'hb874;
    defparam add_1127_15.INJECT1_0 = "NO";
    defparam add_1127_15.INJECT1_1 = "NO";
    CCU2D add_1127_13 (.A0(d_d8[46]), .B0(n6579), .C0(n6580[10]), .D0(d8[46]), 
          .A1(d_d8[47]), .B1(n6579), .C1(n6580[11]), .D1(d8[47]), .CIN(n11179), 
          .COUT(n11180), .S0(d9_71__N_1675[46]), .S1(d9_71__N_1675[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1127_13.INIT0 = 16'hb874;
    defparam add_1127_13.INIT1 = 16'hb874;
    defparam add_1127_13.INJECT1_0 = "NO";
    defparam add_1127_13.INJECT1_1 = "NO";
    CCU2D add_1127_11 (.A0(d_d8[44]), .B0(n6579), .C0(n6580[8]), .D0(d8[44]), 
          .A1(d_d8[45]), .B1(n6579), .C1(n6580[9]), .D1(d8[45]), .CIN(n11178), 
          .COUT(n11179), .S0(d9_71__N_1675[44]), .S1(d9_71__N_1675[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1127_11.INIT0 = 16'hb874;
    defparam add_1127_11.INIT1 = 16'hb874;
    defparam add_1127_11.INJECT1_0 = "NO";
    defparam add_1127_11.INJECT1_1 = "NO";
    CCU2D add_1127_9 (.A0(d_d8[42]), .B0(n6579), .C0(n6580[6]), .D0(d8[42]), 
          .A1(d_d8[43]), .B1(n6579), .C1(n6580[7]), .D1(d8[43]), .CIN(n11177), 
          .COUT(n11178), .S0(d9_71__N_1675[42]), .S1(d9_71__N_1675[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1127_9.INIT0 = 16'hb874;
    defparam add_1127_9.INIT1 = 16'hb874;
    defparam add_1127_9.INJECT1_0 = "NO";
    defparam add_1127_9.INJECT1_1 = "NO";
    CCU2D add_1127_7 (.A0(d_d8[40]), .B0(n6579), .C0(n6580[4]), .D0(d8[40]), 
          .A1(d_d8[41]), .B1(n6579), .C1(n6580[5]), .D1(d8[41]), .CIN(n11176), 
          .COUT(n11177), .S0(d9_71__N_1675[40]), .S1(d9_71__N_1675[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1127_7.INIT0 = 16'hb874;
    defparam add_1127_7.INIT1 = 16'hb874;
    defparam add_1127_7.INJECT1_0 = "NO";
    defparam add_1127_7.INJECT1_1 = "NO";
    CCU2D add_1127_5 (.A0(d_d8[38]), .B0(n6579), .C0(n6580[2]), .D0(d8[38]), 
          .A1(d_d8[39]), .B1(n6579), .C1(n6580[3]), .D1(d8[39]), .CIN(n11175), 
          .COUT(n11176), .S0(d9_71__N_1675[38]), .S1(d9_71__N_1675[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1127_5.INIT0 = 16'hb874;
    defparam add_1127_5.INIT1 = 16'hb874;
    defparam add_1127_5.INJECT1_0 = "NO";
    defparam add_1127_5.INJECT1_1 = "NO";
    CCU2D add_1127_3 (.A0(d_d8[36]), .B0(n6579), .C0(n6580[0]), .D0(d8[36]), 
          .A1(d_d8[37]), .B1(n6579), .C1(n6580[1]), .D1(d8[37]), .CIN(n11174), 
          .COUT(n11175), .S0(d9_71__N_1675[36]), .S1(d9_71__N_1675[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1127_3.INIT0 = 16'hb874;
    defparam add_1127_3.INIT1 = 16'hb874;
    defparam add_1127_3.INJECT1_0 = "NO";
    defparam add_1127_3.INJECT1_1 = "NO";
    CCU2D add_1127_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n6579), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11174));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1127_1.INIT0 = 16'hF000;
    defparam add_1127_1.INIT1 = 16'h0555;
    defparam add_1127_1.INJECT1_0 = "NO";
    defparam add_1127_1.INJECT1_1 = "NO";
    CCU2D add_1131_37 (.A0(d9[71]), .B0(d_d9[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11170), 
          .S0(n6732[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1131_37.INIT0 = 16'h5999;
    defparam add_1131_37.INIT1 = 16'h0000;
    defparam add_1131_37.INJECT1_0 = "NO";
    defparam add_1131_37.INJECT1_1 = "NO";
    CCU2D add_1131_35 (.A0(d9[69]), .B0(d_d9[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[70]), .B1(d_d9[70]), .C1(GND_net), .D1(GND_net), .CIN(n11169), 
          .COUT(n11170), .S0(n6732[33]), .S1(n6732[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1131_35.INIT0 = 16'h5999;
    defparam add_1131_35.INIT1 = 16'h5999;
    defparam add_1131_35.INJECT1_0 = "NO";
    defparam add_1131_35.INJECT1_1 = "NO";
    CCU2D add_1131_33 (.A0(d9[67]), .B0(d_d9[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[68]), .B1(d_d9[68]), .C1(GND_net), .D1(GND_net), .CIN(n11168), 
          .COUT(n11169), .S0(n6732[31]), .S1(n6732[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1131_33.INIT0 = 16'h5999;
    defparam add_1131_33.INIT1 = 16'h5999;
    defparam add_1131_33.INJECT1_0 = "NO";
    defparam add_1131_33.INJECT1_1 = "NO";
    CCU2D add_1131_31 (.A0(d9[65]), .B0(d_d9[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[66]), .B1(d_d9[66]), .C1(GND_net), .D1(GND_net), .CIN(n11167), 
          .COUT(n11168), .S0(n6732[29]), .S1(n6732[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1131_31.INIT0 = 16'h5999;
    defparam add_1131_31.INIT1 = 16'h5999;
    defparam add_1131_31.INJECT1_0 = "NO";
    defparam add_1131_31.INJECT1_1 = "NO";
    CCU2D add_1131_29 (.A0(d9[63]), .B0(d_d9[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[64]), .B1(d_d9[64]), .C1(GND_net), .D1(GND_net), .CIN(n11166), 
          .COUT(n11167), .S0(n6732[27]), .S1(n6732[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1131_29.INIT0 = 16'h5999;
    defparam add_1131_29.INIT1 = 16'h5999;
    defparam add_1131_29.INJECT1_0 = "NO";
    defparam add_1131_29.INJECT1_1 = "NO";
    CCU2D add_1131_27 (.A0(d9[61]), .B0(d_d9[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[62]), .B1(d_d9[62]), .C1(GND_net), .D1(GND_net), .CIN(n11165), 
          .COUT(n11166), .S0(n6732[25]), .S1(n6732[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1131_27.INIT0 = 16'h5999;
    defparam add_1131_27.INIT1 = 16'h5999;
    defparam add_1131_27.INJECT1_0 = "NO";
    defparam add_1131_27.INJECT1_1 = "NO";
    CCU2D add_1131_25 (.A0(d9[59]), .B0(d_d9[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[60]), .B1(d_d9[60]), .C1(GND_net), .D1(GND_net), .CIN(n11164), 
          .COUT(n11165), .S0(n6732[23]), .S1(n6732[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1131_25.INIT0 = 16'h5999;
    defparam add_1131_25.INIT1 = 16'h5999;
    defparam add_1131_25.INJECT1_0 = "NO";
    defparam add_1131_25.INJECT1_1 = "NO";
    CCU2D add_1131_23 (.A0(d9[57]), .B0(d_d9[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[58]), .B1(d_d9[58]), .C1(GND_net), .D1(GND_net), .CIN(n11163), 
          .COUT(n11164), .S0(n6732[21]), .S1(n6732[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1131_23.INIT0 = 16'h5999;
    defparam add_1131_23.INIT1 = 16'h5999;
    defparam add_1131_23.INJECT1_0 = "NO";
    defparam add_1131_23.INJECT1_1 = "NO";
    CCU2D add_1131_21 (.A0(d9[55]), .B0(d_d9[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[56]), .B1(d_d9[56]), .C1(GND_net), .D1(GND_net), .CIN(n11162), 
          .COUT(n11163));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1131_21.INIT0 = 16'h5999;
    defparam add_1131_21.INIT1 = 16'h5999;
    defparam add_1131_21.INJECT1_0 = "NO";
    defparam add_1131_21.INJECT1_1 = "NO";
    CCU2D add_1131_19 (.A0(d9[53]), .B0(d_d9[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[54]), .B1(d_d9[54]), .C1(GND_net), .D1(GND_net), .CIN(n11161), 
          .COUT(n11162));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1131_19.INIT0 = 16'h5999;
    defparam add_1131_19.INIT1 = 16'h5999;
    defparam add_1131_19.INJECT1_0 = "NO";
    defparam add_1131_19.INJECT1_1 = "NO";
    CCU2D add_1131_17 (.A0(d9[51]), .B0(d_d9[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[52]), .B1(d_d9[52]), .C1(GND_net), .D1(GND_net), .CIN(n11160), 
          .COUT(n11161));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1131_17.INIT0 = 16'h5999;
    defparam add_1131_17.INIT1 = 16'h5999;
    defparam add_1131_17.INJECT1_0 = "NO";
    defparam add_1131_17.INJECT1_1 = "NO";
    CCU2D add_1131_15 (.A0(d9[49]), .B0(d_d9[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[50]), .B1(d_d9[50]), .C1(GND_net), .D1(GND_net), .CIN(n11159), 
          .COUT(n11160));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1131_15.INIT0 = 16'h5999;
    defparam add_1131_15.INIT1 = 16'h5999;
    defparam add_1131_15.INJECT1_0 = "NO";
    defparam add_1131_15.INJECT1_1 = "NO";
    CCU2D add_1131_13 (.A0(d9[47]), .B0(d_d9[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[48]), .B1(d_d9[48]), .C1(GND_net), .D1(GND_net), .CIN(n11158), 
          .COUT(n11159));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1131_13.INIT0 = 16'h5999;
    defparam add_1131_13.INIT1 = 16'h5999;
    defparam add_1131_13.INJECT1_0 = "NO";
    defparam add_1131_13.INJECT1_1 = "NO";
    CCU2D add_1131_11 (.A0(d9[45]), .B0(d_d9[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[46]), .B1(d_d9[46]), .C1(GND_net), .D1(GND_net), .CIN(n11157), 
          .COUT(n11158));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1131_11.INIT0 = 16'h5999;
    defparam add_1131_11.INIT1 = 16'h5999;
    defparam add_1131_11.INJECT1_0 = "NO";
    defparam add_1131_11.INJECT1_1 = "NO";
    CCU2D add_1131_9 (.A0(d9[43]), .B0(d_d9[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[44]), .B1(d_d9[44]), .C1(GND_net), .D1(GND_net), .CIN(n11156), 
          .COUT(n11157));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1131_9.INIT0 = 16'h5999;
    defparam add_1131_9.INIT1 = 16'h5999;
    defparam add_1131_9.INJECT1_0 = "NO";
    defparam add_1131_9.INJECT1_1 = "NO";
    CCU2D add_1131_7 (.A0(d9[41]), .B0(d_d9[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[42]), .B1(d_d9[42]), .C1(GND_net), .D1(GND_net), .CIN(n11155), 
          .COUT(n11156));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1131_7.INIT0 = 16'h5999;
    defparam add_1131_7.INIT1 = 16'h5999;
    defparam add_1131_7.INJECT1_0 = "NO";
    defparam add_1131_7.INJECT1_1 = "NO";
    CCU2D add_1131_5 (.A0(d9[39]), .B0(d_d9[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[40]), .B1(d_d9[40]), .C1(GND_net), .D1(GND_net), .CIN(n11154), 
          .COUT(n11155));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1131_5.INIT0 = 16'h5999;
    defparam add_1131_5.INIT1 = 16'h5999;
    defparam add_1131_5.INJECT1_0 = "NO";
    defparam add_1131_5.INJECT1_1 = "NO";
    CCU2D add_1131_3 (.A0(d9[37]), .B0(d_d9[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[38]), .B1(d_d9[38]), .C1(GND_net), .D1(GND_net), .CIN(n11153), 
          .COUT(n11154));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1131_3.INIT0 = 16'h5999;
    defparam add_1131_3.INIT1 = 16'h5999;
    defparam add_1131_3.INJECT1_0 = "NO";
    defparam add_1131_3.INJECT1_1 = "NO";
    CCU2D add_1131_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d9[36]), .B1(d_d9[36]), .C1(GND_net), .D1(GND_net), .COUT(n11153));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1131_1.INIT0 = 16'hF000;
    defparam add_1131_1.INIT1 = 16'h5999;
    defparam add_1131_1.INJECT1_0 = "NO";
    defparam add_1131_1.INJECT1_1 = "NO";
    CCU2D add_1132_37 (.A0(d9[71]), .B0(d_d9[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11152), 
          .S0(n6770[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1132_37.INIT0 = 16'h5999;
    defparam add_1132_37.INIT1 = 16'h0000;
    defparam add_1132_37.INJECT1_0 = "NO";
    defparam add_1132_37.INJECT1_1 = "NO";
    CCU2D add_1132_35 (.A0(d9[69]), .B0(d_d9[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[70]), .B1(d_d9[70]), .C1(GND_net), .D1(GND_net), .CIN(n11151), 
          .COUT(n11152), .S0(n6770[33]), .S1(n6770[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1132_35.INIT0 = 16'h5999;
    defparam add_1132_35.INIT1 = 16'h5999;
    defparam add_1132_35.INJECT1_0 = "NO";
    defparam add_1132_35.INJECT1_1 = "NO";
    CCU2D add_1132_33 (.A0(d9[67]), .B0(d_d9[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[68]), .B1(d_d9[68]), .C1(GND_net), .D1(GND_net), .CIN(n11150), 
          .COUT(n11151), .S0(n6770[31]), .S1(n6770[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1132_33.INIT0 = 16'h5999;
    defparam add_1132_33.INIT1 = 16'h5999;
    defparam add_1132_33.INJECT1_0 = "NO";
    defparam add_1132_33.INJECT1_1 = "NO";
    CCU2D add_1132_31 (.A0(d9[65]), .B0(d_d9[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[66]), .B1(d_d9[66]), .C1(GND_net), .D1(GND_net), .CIN(n11149), 
          .COUT(n11150), .S0(n6770[29]), .S1(n6770[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1132_31.INIT0 = 16'h5999;
    defparam add_1132_31.INIT1 = 16'h5999;
    defparam add_1132_31.INJECT1_0 = "NO";
    defparam add_1132_31.INJECT1_1 = "NO";
    CCU2D add_1132_29 (.A0(d9[63]), .B0(d_d9[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[64]), .B1(d_d9[64]), .C1(GND_net), .D1(GND_net), .CIN(n11148), 
          .COUT(n11149), .S0(n6770[27]), .S1(n6770[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1132_29.INIT0 = 16'h5999;
    defparam add_1132_29.INIT1 = 16'h5999;
    defparam add_1132_29.INJECT1_0 = "NO";
    defparam add_1132_29.INJECT1_1 = "NO";
    CCU2D add_1132_27 (.A0(d9[61]), .B0(d_d9[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[62]), .B1(d_d9[62]), .C1(GND_net), .D1(GND_net), .CIN(n11147), 
          .COUT(n11148), .S0(n6770[25]), .S1(n6770[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1132_27.INIT0 = 16'h5999;
    defparam add_1132_27.INIT1 = 16'h5999;
    defparam add_1132_27.INJECT1_0 = "NO";
    defparam add_1132_27.INJECT1_1 = "NO";
    CCU2D add_1132_25 (.A0(d9[59]), .B0(d_d9[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[60]), .B1(d_d9[60]), .C1(GND_net), .D1(GND_net), .CIN(n11146), 
          .COUT(n11147), .S0(n6770[23]), .S1(n6770[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1132_25.INIT0 = 16'h5999;
    defparam add_1132_25.INIT1 = 16'h5999;
    defparam add_1132_25.INJECT1_0 = "NO";
    defparam add_1132_25.INJECT1_1 = "NO";
    CCU2D add_1132_23 (.A0(d9[57]), .B0(d_d9[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[58]), .B1(d_d9[58]), .C1(GND_net), .D1(GND_net), .CIN(n11145), 
          .COUT(n11146), .S0(n6770[21]), .S1(n6770[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1132_23.INIT0 = 16'h5999;
    defparam add_1132_23.INIT1 = 16'h5999;
    defparam add_1132_23.INJECT1_0 = "NO";
    defparam add_1132_23.INJECT1_1 = "NO";
    CCU2D add_1132_21 (.A0(d9[55]), .B0(d_d9[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[56]), .B1(d_d9[56]), .C1(GND_net), .D1(GND_net), .CIN(n11144), 
          .COUT(n11145));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1132_21.INIT0 = 16'h5999;
    defparam add_1132_21.INIT1 = 16'h5999;
    defparam add_1132_21.INJECT1_0 = "NO";
    defparam add_1132_21.INJECT1_1 = "NO";
    CCU2D add_1132_19 (.A0(d9[53]), .B0(d_d9[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[54]), .B1(d_d9[54]), .C1(GND_net), .D1(GND_net), .CIN(n11143), 
          .COUT(n11144));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1132_19.INIT0 = 16'h5999;
    defparam add_1132_19.INIT1 = 16'h5999;
    defparam add_1132_19.INJECT1_0 = "NO";
    defparam add_1132_19.INJECT1_1 = "NO";
    CCU2D add_1132_17 (.A0(d9[51]), .B0(d_d9[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[52]), .B1(d_d9[52]), .C1(GND_net), .D1(GND_net), .CIN(n11142), 
          .COUT(n11143));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1132_17.INIT0 = 16'h5999;
    defparam add_1132_17.INIT1 = 16'h5999;
    defparam add_1132_17.INJECT1_0 = "NO";
    defparam add_1132_17.INJECT1_1 = "NO";
    CCU2D add_1132_15 (.A0(d9[49]), .B0(d_d9[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[50]), .B1(d_d9[50]), .C1(GND_net), .D1(GND_net), .CIN(n11141), 
          .COUT(n11142));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1132_15.INIT0 = 16'h5999;
    defparam add_1132_15.INIT1 = 16'h5999;
    defparam add_1132_15.INJECT1_0 = "NO";
    defparam add_1132_15.INJECT1_1 = "NO";
    CCU2D add_1132_13 (.A0(d9[47]), .B0(d_d9[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[48]), .B1(d_d9[48]), .C1(GND_net), .D1(GND_net), .CIN(n11140), 
          .COUT(n11141));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1132_13.INIT0 = 16'h5999;
    defparam add_1132_13.INIT1 = 16'h5999;
    defparam add_1132_13.INJECT1_0 = "NO";
    defparam add_1132_13.INJECT1_1 = "NO";
    CCU2D add_1132_11 (.A0(d9[45]), .B0(d_d9[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[46]), .B1(d_d9[46]), .C1(GND_net), .D1(GND_net), .CIN(n11139), 
          .COUT(n11140));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1132_11.INIT0 = 16'h5999;
    defparam add_1132_11.INIT1 = 16'h5999;
    defparam add_1132_11.INJECT1_0 = "NO";
    defparam add_1132_11.INJECT1_1 = "NO";
    CCU2D add_1132_9 (.A0(d9[43]), .B0(d_d9[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[44]), .B1(d_d9[44]), .C1(GND_net), .D1(GND_net), .CIN(n11138), 
          .COUT(n11139));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1132_9.INIT0 = 16'h5999;
    defparam add_1132_9.INIT1 = 16'h5999;
    defparam add_1132_9.INJECT1_0 = "NO";
    defparam add_1132_9.INJECT1_1 = "NO";
    CCU2D add_1132_7 (.A0(d9[41]), .B0(d_d9[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[42]), .B1(d_d9[42]), .C1(GND_net), .D1(GND_net), .CIN(n11137), 
          .COUT(n11138));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1132_7.INIT0 = 16'h5999;
    defparam add_1132_7.INIT1 = 16'h5999;
    defparam add_1132_7.INJECT1_0 = "NO";
    defparam add_1132_7.INJECT1_1 = "NO";
    CCU2D add_1132_5 (.A0(d9[39]), .B0(d_d9[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[40]), .B1(d_d9[40]), .C1(GND_net), .D1(GND_net), .CIN(n11136), 
          .COUT(n11137));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1132_5.INIT0 = 16'h5999;
    defparam add_1132_5.INIT1 = 16'h5999;
    defparam add_1132_5.INJECT1_0 = "NO";
    defparam add_1132_5.INJECT1_1 = "NO";
    CCU2D add_1132_3 (.A0(d9[37]), .B0(d_d9[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[38]), .B1(d_d9[38]), .C1(GND_net), .D1(GND_net), .CIN(n11135), 
          .COUT(n11136));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1132_3.INIT0 = 16'h5999;
    defparam add_1132_3.INIT1 = 16'h5999;
    defparam add_1132_3.INJECT1_0 = "NO";
    defparam add_1132_3.INJECT1_1 = "NO";
    CCU2D add_1132_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d9[36]), .B1(d_d9[36]), .C1(GND_net), .D1(GND_net), .COUT(n11135));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1132_1.INIT0 = 16'h0000;
    defparam add_1132_1.INIT1 = 16'h5999;
    defparam add_1132_1.INJECT1_0 = "NO";
    defparam add_1132_1.INJECT1_1 = "NO";
    FD1S3IX count__i2 (.D(n375[2]), .CK(osc_clk), .CD(n8436), .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n375[3]), .CK(osc_clk), .CD(n8436), .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n375[4]), .CK(osc_clk), .CD(n8436), .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n375[5]), .CK(osc_clk), .CD(n8436), .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n375[6]), .CK(osc_clk), .CD(n8436), .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n375[7]), .CK(osc_clk), .CD(n8436), .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n375[8]), .CK(osc_clk), .CD(n8436), .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n375[9]), .CK(osc_clk), .CD(n8436), .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n375[10]), .CK(osc_clk), .CD(n8436), .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_15__N_1442[11]), .CK(osc_clk), .CD(count_15__N_1458), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(n375[12]), .CK(osc_clk), .CD(n8436), .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(n375[13]), .CK(osc_clk), .CD(n8436), .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(n375[14]), .CK(osc_clk), .CD(n8436), .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(n375[15]), .CK(osc_clk), .CD(n8436), .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i15.GSR = "ENABLED";
    CCU2D add_10_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10938), 
          .S0(n375[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_17.INIT0 = 16'h5aaa;
    defparam add_10_17.INIT1 = 16'h0000;
    defparam add_10_17.INJECT1_0 = "NO";
    defparam add_10_17.INJECT1_1 = "NO";
    CCU2D add_10_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n10937), .COUT(n10938), .S0(n375[13]), .S1(n375[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_15.INIT0 = 16'h5aaa;
    defparam add_10_15.INIT1 = 16'h5aaa;
    defparam add_10_15.INJECT1_0 = "NO";
    defparam add_10_15.INJECT1_1 = "NO";
    CCU2D add_10_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n10936), .COUT(n10937), .S0(n375[11]), .S1(n375[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_13.INIT0 = 16'h5aaa;
    defparam add_10_13.INIT1 = 16'h5aaa;
    defparam add_10_13.INJECT1_0 = "NO";
    defparam add_10_13.INJECT1_1 = "NO";
    CCU2D add_10_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n10935), .COUT(n10936), .S0(n375[9]), .S1(n375[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_11.INIT0 = 16'h5aaa;
    defparam add_10_11.INIT1 = 16'h5aaa;
    defparam add_10_11.INJECT1_0 = "NO";
    defparam add_10_11.INJECT1_1 = "NO";
    CCU2D add_10_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10934), 
          .COUT(n10935), .S0(n375[7]), .S1(n375[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_9.INIT0 = 16'h5aaa;
    defparam add_10_9.INIT1 = 16'h5aaa;
    defparam add_10_9.INJECT1_0 = "NO";
    defparam add_10_9.INJECT1_1 = "NO";
    CCU2D add_10_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10933), 
          .COUT(n10934), .S0(n375[5]), .S1(n375[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_7.INIT0 = 16'h5aaa;
    defparam add_10_7.INIT1 = 16'h5aaa;
    defparam add_10_7.INJECT1_0 = "NO";
    defparam add_10_7.INJECT1_1 = "NO";
    CCU2D add_10_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10932), 
          .COUT(n10933), .S0(n375[3]), .S1(n375[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_5.INIT0 = 16'h5aaa;
    defparam add_10_5.INIT1 = 16'h5aaa;
    defparam add_10_5.INJECT1_0 = "NO";
    defparam add_10_5.INJECT1_1 = "NO";
    CCU2D add_10_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10931), 
          .COUT(n10932), .S0(n375[1]), .S1(n375[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_3.INIT0 = 16'h5aaa;
    defparam add_10_3.INIT1 = 16'h5aaa;
    defparam add_10_3.INJECT1_0 = "NO";
    defparam add_10_3.INJECT1_1 = "NO";
    CCU2D add_10_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n10931), 
          .S1(n375[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_1.INIT0 = 16'hF000;
    defparam add_10_1.INIT1 = 16'h5555;
    defparam add_10_1.INJECT1_0 = "NO";
    defparam add_10_1.INJECT1_1 = "NO";
    CCU2D add_1095_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10912), 
          .S0(n5667));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1095_cout.INIT0 = 16'h0000;
    defparam add_1095_cout.INIT1 = 16'h0000;
    defparam add_1095_cout.INJECT1_0 = "NO";
    defparam add_1095_cout.INJECT1_1 = "NO";
    CCU2D add_1095_36 (.A0(d4[34]), .B0(d5[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[35]), .B1(d5[35]), .C1(GND_net), .D1(GND_net), .CIN(n10911), 
          .COUT(n10912), .S0(d5_71__N_706[34]), .S1(d5_71__N_706[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1095_36.INIT0 = 16'h5666;
    defparam add_1095_36.INIT1 = 16'h5666;
    defparam add_1095_36.INJECT1_0 = "NO";
    defparam add_1095_36.INJECT1_1 = "NO";
    CCU2D add_1095_34 (.A0(d4[32]), .B0(d5[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[33]), .B1(d5[33]), .C1(GND_net), .D1(GND_net), .CIN(n10910), 
          .COUT(n10911), .S0(d5_71__N_706[32]), .S1(d5_71__N_706[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1095_34.INIT0 = 16'h5666;
    defparam add_1095_34.INIT1 = 16'h5666;
    defparam add_1095_34.INJECT1_0 = "NO";
    defparam add_1095_34.INJECT1_1 = "NO";
    CCU2D add_1095_32 (.A0(d4[30]), .B0(d5[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[31]), .B1(d5[31]), .C1(GND_net), .D1(GND_net), .CIN(n10909), 
          .COUT(n10910), .S0(d5_71__N_706[30]), .S1(d5_71__N_706[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1095_32.INIT0 = 16'h5666;
    defparam add_1095_32.INIT1 = 16'h5666;
    defparam add_1095_32.INJECT1_0 = "NO";
    defparam add_1095_32.INJECT1_1 = "NO";
    CCU2D add_1095_30 (.A0(d4[28]), .B0(d5[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[29]), .B1(d5[29]), .C1(GND_net), .D1(GND_net), .CIN(n10908), 
          .COUT(n10909), .S0(d5_71__N_706[28]), .S1(d5_71__N_706[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1095_30.INIT0 = 16'h5666;
    defparam add_1095_30.INIT1 = 16'h5666;
    defparam add_1095_30.INJECT1_0 = "NO";
    defparam add_1095_30.INJECT1_1 = "NO";
    CCU2D add_1095_28 (.A0(d4[26]), .B0(d5[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[27]), .B1(d5[27]), .C1(GND_net), .D1(GND_net), .CIN(n10907), 
          .COUT(n10908), .S0(d5_71__N_706[26]), .S1(d5_71__N_706[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1095_28.INIT0 = 16'h5666;
    defparam add_1095_28.INIT1 = 16'h5666;
    defparam add_1095_28.INJECT1_0 = "NO";
    defparam add_1095_28.INJECT1_1 = "NO";
    CCU2D add_1095_26 (.A0(d4[24]), .B0(d5[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[25]), .B1(d5[25]), .C1(GND_net), .D1(GND_net), .CIN(n10906), 
          .COUT(n10907), .S0(d5_71__N_706[24]), .S1(d5_71__N_706[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1095_26.INIT0 = 16'h5666;
    defparam add_1095_26.INIT1 = 16'h5666;
    defparam add_1095_26.INJECT1_0 = "NO";
    defparam add_1095_26.INJECT1_1 = "NO";
    CCU2D add_1095_24 (.A0(d4[22]), .B0(d5[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[23]), .B1(d5[23]), .C1(GND_net), .D1(GND_net), .CIN(n10905), 
          .COUT(n10906), .S0(d5_71__N_706[22]), .S1(d5_71__N_706[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1095_24.INIT0 = 16'h5666;
    defparam add_1095_24.INIT1 = 16'h5666;
    defparam add_1095_24.INJECT1_0 = "NO";
    defparam add_1095_24.INJECT1_1 = "NO";
    CCU2D add_1095_22 (.A0(d4[20]), .B0(d5[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[21]), .B1(d5[21]), .C1(GND_net), .D1(GND_net), .CIN(n10904), 
          .COUT(n10905), .S0(d5_71__N_706[20]), .S1(d5_71__N_706[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1095_22.INIT0 = 16'h5666;
    defparam add_1095_22.INIT1 = 16'h5666;
    defparam add_1095_22.INJECT1_0 = "NO";
    defparam add_1095_22.INJECT1_1 = "NO";
    CCU2D add_1095_20 (.A0(d4[18]), .B0(d5[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[19]), .B1(d5[19]), .C1(GND_net), .D1(GND_net), .CIN(n10903), 
          .COUT(n10904), .S0(d5_71__N_706[18]), .S1(d5_71__N_706[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1095_20.INIT0 = 16'h5666;
    defparam add_1095_20.INIT1 = 16'h5666;
    defparam add_1095_20.INJECT1_0 = "NO";
    defparam add_1095_20.INJECT1_1 = "NO";
    CCU2D add_1095_18 (.A0(d4[16]), .B0(d5[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[17]), .B1(d5[17]), .C1(GND_net), .D1(GND_net), .CIN(n10902), 
          .COUT(n10903), .S0(d5_71__N_706[16]), .S1(d5_71__N_706[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1095_18.INIT0 = 16'h5666;
    defparam add_1095_18.INIT1 = 16'h5666;
    defparam add_1095_18.INJECT1_0 = "NO";
    defparam add_1095_18.INJECT1_1 = "NO";
    CCU2D add_1095_16 (.A0(d4[14]), .B0(d5[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[15]), .B1(d5[15]), .C1(GND_net), .D1(GND_net), .CIN(n10901), 
          .COUT(n10902), .S0(d5_71__N_706[14]), .S1(d5_71__N_706[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1095_16.INIT0 = 16'h5666;
    defparam add_1095_16.INIT1 = 16'h5666;
    defparam add_1095_16.INJECT1_0 = "NO";
    defparam add_1095_16.INJECT1_1 = "NO";
    CCU2D add_1095_14 (.A0(d4[12]), .B0(d5[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[13]), .B1(d5[13]), .C1(GND_net), .D1(GND_net), .CIN(n10900), 
          .COUT(n10901), .S0(d5_71__N_706[12]), .S1(d5_71__N_706[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1095_14.INIT0 = 16'h5666;
    defparam add_1095_14.INIT1 = 16'h5666;
    defparam add_1095_14.INJECT1_0 = "NO";
    defparam add_1095_14.INJECT1_1 = "NO";
    CCU2D add_1095_12 (.A0(d4[10]), .B0(d5[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[11]), .B1(d5[11]), .C1(GND_net), .D1(GND_net), .CIN(n10899), 
          .COUT(n10900), .S0(d5_71__N_706[10]), .S1(d5_71__N_706[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1095_12.INIT0 = 16'h5666;
    defparam add_1095_12.INIT1 = 16'h5666;
    defparam add_1095_12.INJECT1_0 = "NO";
    defparam add_1095_12.INJECT1_1 = "NO";
    CCU2D add_1095_10 (.A0(d4[8]), .B0(d5[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[9]), .B1(d5[9]), .C1(GND_net), .D1(GND_net), .CIN(n10898), 
          .COUT(n10899), .S0(d5_71__N_706[8]), .S1(d5_71__N_706[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1095_10.INIT0 = 16'h5666;
    defparam add_1095_10.INIT1 = 16'h5666;
    defparam add_1095_10.INJECT1_0 = "NO";
    defparam add_1095_10.INJECT1_1 = "NO";
    CCU2D add_1095_8 (.A0(d4[6]), .B0(d5[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[7]), .B1(d5[7]), .C1(GND_net), .D1(GND_net), .CIN(n10897), 
          .COUT(n10898), .S0(d5_71__N_706[6]), .S1(d5_71__N_706[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1095_8.INIT0 = 16'h5666;
    defparam add_1095_8.INIT1 = 16'h5666;
    defparam add_1095_8.INJECT1_0 = "NO";
    defparam add_1095_8.INJECT1_1 = "NO";
    CCU2D add_1095_6 (.A0(d4[4]), .B0(d5[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[5]), .B1(d5[5]), .C1(GND_net), .D1(GND_net), .CIN(n10896), 
          .COUT(n10897), .S0(d5_71__N_706[4]), .S1(d5_71__N_706[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1095_6.INIT0 = 16'h5666;
    defparam add_1095_6.INIT1 = 16'h5666;
    defparam add_1095_6.INJECT1_0 = "NO";
    defparam add_1095_6.INJECT1_1 = "NO";
    CCU2D add_1095_4 (.A0(d4[2]), .B0(d5[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[3]), .B1(d5[3]), .C1(GND_net), .D1(GND_net), .CIN(n10895), 
          .COUT(n10896), .S0(d5_71__N_706[2]), .S1(d5_71__N_706[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1095_4.INIT0 = 16'h5666;
    defparam add_1095_4.INIT1 = 16'h5666;
    defparam add_1095_4.INJECT1_0 = "NO";
    defparam add_1095_4.INJECT1_1 = "NO";
    CCU2D add_1095_2 (.A0(d4[0]), .B0(d5[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[1]), .B1(d5[1]), .C1(GND_net), .D1(GND_net), .COUT(n10895), 
          .S1(d5_71__N_706[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1095_2.INIT0 = 16'h7000;
    defparam add_1095_2.INIT1 = 16'h5666;
    defparam add_1095_2.INJECT1_0 = "NO";
    defparam add_1095_2.INJECT1_1 = "NO";
    CCU2D add_1090_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10893), 
          .S0(n5515));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1090_cout.INIT0 = 16'h0000;
    defparam add_1090_cout.INIT1 = 16'h0000;
    defparam add_1090_cout.INJECT1_0 = "NO";
    defparam add_1090_cout.INJECT1_1 = "NO";
    CCU2D add_1090_36 (.A0(d3[34]), .B0(d4[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[35]), .B1(d4[35]), .C1(GND_net), .D1(GND_net), .CIN(n10892), 
          .COUT(n10893), .S0(d4_71__N_634[34]), .S1(d4_71__N_634[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1090_36.INIT0 = 16'h5666;
    defparam add_1090_36.INIT1 = 16'h5666;
    defparam add_1090_36.INJECT1_0 = "NO";
    defparam add_1090_36.INJECT1_1 = "NO";
    CCU2D add_1090_34 (.A0(d3[32]), .B0(d4[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[33]), .B1(d4[33]), .C1(GND_net), .D1(GND_net), .CIN(n10891), 
          .COUT(n10892), .S0(d4_71__N_634[32]), .S1(d4_71__N_634[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1090_34.INIT0 = 16'h5666;
    defparam add_1090_34.INIT1 = 16'h5666;
    defparam add_1090_34.INJECT1_0 = "NO";
    defparam add_1090_34.INJECT1_1 = "NO";
    CCU2D add_1090_32 (.A0(d3[30]), .B0(d4[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[31]), .B1(d4[31]), .C1(GND_net), .D1(GND_net), .CIN(n10890), 
          .COUT(n10891), .S0(d4_71__N_634[30]), .S1(d4_71__N_634[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1090_32.INIT0 = 16'h5666;
    defparam add_1090_32.INIT1 = 16'h5666;
    defparam add_1090_32.INJECT1_0 = "NO";
    defparam add_1090_32.INJECT1_1 = "NO";
    CCU2D add_1090_30 (.A0(d3[28]), .B0(d4[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[29]), .B1(d4[29]), .C1(GND_net), .D1(GND_net), .CIN(n10889), 
          .COUT(n10890), .S0(d4_71__N_634[28]), .S1(d4_71__N_634[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1090_30.INIT0 = 16'h5666;
    defparam add_1090_30.INIT1 = 16'h5666;
    defparam add_1090_30.INJECT1_0 = "NO";
    defparam add_1090_30.INJECT1_1 = "NO";
    CCU2D add_1090_28 (.A0(d3[26]), .B0(d4[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[27]), .B1(d4[27]), .C1(GND_net), .D1(GND_net), .CIN(n10888), 
          .COUT(n10889), .S0(d4_71__N_634[26]), .S1(d4_71__N_634[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1090_28.INIT0 = 16'h5666;
    defparam add_1090_28.INIT1 = 16'h5666;
    defparam add_1090_28.INJECT1_0 = "NO";
    defparam add_1090_28.INJECT1_1 = "NO";
    CCU2D add_1090_26 (.A0(d3[24]), .B0(d4[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[25]), .B1(d4[25]), .C1(GND_net), .D1(GND_net), .CIN(n10887), 
          .COUT(n10888), .S0(d4_71__N_634[24]), .S1(d4_71__N_634[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1090_26.INIT0 = 16'h5666;
    defparam add_1090_26.INIT1 = 16'h5666;
    defparam add_1090_26.INJECT1_0 = "NO";
    defparam add_1090_26.INJECT1_1 = "NO";
    CCU2D add_1090_24 (.A0(d3[22]), .B0(d4[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[23]), .B1(d4[23]), .C1(GND_net), .D1(GND_net), .CIN(n10886), 
          .COUT(n10887), .S0(d4_71__N_634[22]), .S1(d4_71__N_634[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1090_24.INIT0 = 16'h5666;
    defparam add_1090_24.INIT1 = 16'h5666;
    defparam add_1090_24.INJECT1_0 = "NO";
    defparam add_1090_24.INJECT1_1 = "NO";
    CCU2D add_1090_22 (.A0(d3[20]), .B0(d4[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[21]), .B1(d4[21]), .C1(GND_net), .D1(GND_net), .CIN(n10885), 
          .COUT(n10886), .S0(d4_71__N_634[20]), .S1(d4_71__N_634[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1090_22.INIT0 = 16'h5666;
    defparam add_1090_22.INIT1 = 16'h5666;
    defparam add_1090_22.INJECT1_0 = "NO";
    defparam add_1090_22.INJECT1_1 = "NO";
    CCU2D add_1090_20 (.A0(d3[18]), .B0(d4[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[19]), .B1(d4[19]), .C1(GND_net), .D1(GND_net), .CIN(n10884), 
          .COUT(n10885), .S0(d4_71__N_634[18]), .S1(d4_71__N_634[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1090_20.INIT0 = 16'h5666;
    defparam add_1090_20.INIT1 = 16'h5666;
    defparam add_1090_20.INJECT1_0 = "NO";
    defparam add_1090_20.INJECT1_1 = "NO";
    CCU2D add_1090_18 (.A0(d3[16]), .B0(d4[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[17]), .B1(d4[17]), .C1(GND_net), .D1(GND_net), .CIN(n10883), 
          .COUT(n10884), .S0(d4_71__N_634[16]), .S1(d4_71__N_634[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1090_18.INIT0 = 16'h5666;
    defparam add_1090_18.INIT1 = 16'h5666;
    defparam add_1090_18.INJECT1_0 = "NO";
    defparam add_1090_18.INJECT1_1 = "NO";
    CCU2D add_1090_16 (.A0(d3[14]), .B0(d4[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[15]), .B1(d4[15]), .C1(GND_net), .D1(GND_net), .CIN(n10882), 
          .COUT(n10883), .S0(d4_71__N_634[14]), .S1(d4_71__N_634[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1090_16.INIT0 = 16'h5666;
    defparam add_1090_16.INIT1 = 16'h5666;
    defparam add_1090_16.INJECT1_0 = "NO";
    defparam add_1090_16.INJECT1_1 = "NO";
    CCU2D add_1090_14 (.A0(d3[12]), .B0(d4[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[13]), .B1(d4[13]), .C1(GND_net), .D1(GND_net), .CIN(n10881), 
          .COUT(n10882), .S0(d4_71__N_634[12]), .S1(d4_71__N_634[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1090_14.INIT0 = 16'h5666;
    defparam add_1090_14.INIT1 = 16'h5666;
    defparam add_1090_14.INJECT1_0 = "NO";
    defparam add_1090_14.INJECT1_1 = "NO";
    CCU2D add_1090_12 (.A0(d3[10]), .B0(d4[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[11]), .B1(d4[11]), .C1(GND_net), .D1(GND_net), .CIN(n10880), 
          .COUT(n10881), .S0(d4_71__N_634[10]), .S1(d4_71__N_634[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1090_12.INIT0 = 16'h5666;
    defparam add_1090_12.INIT1 = 16'h5666;
    defparam add_1090_12.INJECT1_0 = "NO";
    defparam add_1090_12.INJECT1_1 = "NO";
    CCU2D add_1090_10 (.A0(d3[8]), .B0(d4[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[9]), .B1(d4[9]), .C1(GND_net), .D1(GND_net), .CIN(n10879), 
          .COUT(n10880), .S0(d4_71__N_634[8]), .S1(d4_71__N_634[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1090_10.INIT0 = 16'h5666;
    defparam add_1090_10.INIT1 = 16'h5666;
    defparam add_1090_10.INJECT1_0 = "NO";
    defparam add_1090_10.INJECT1_1 = "NO";
    CCU2D add_1090_8 (.A0(d3[6]), .B0(d4[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[7]), .B1(d4[7]), .C1(GND_net), .D1(GND_net), .CIN(n10878), 
          .COUT(n10879), .S0(d4_71__N_634[6]), .S1(d4_71__N_634[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1090_8.INIT0 = 16'h5666;
    defparam add_1090_8.INIT1 = 16'h5666;
    defparam add_1090_8.INJECT1_0 = "NO";
    defparam add_1090_8.INJECT1_1 = "NO";
    CCU2D add_1090_6 (.A0(d3[4]), .B0(d4[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[5]), .B1(d4[5]), .C1(GND_net), .D1(GND_net), .CIN(n10877), 
          .COUT(n10878), .S0(d4_71__N_634[4]), .S1(d4_71__N_634[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1090_6.INIT0 = 16'h5666;
    defparam add_1090_6.INIT1 = 16'h5666;
    defparam add_1090_6.INJECT1_0 = "NO";
    defparam add_1090_6.INJECT1_1 = "NO";
    CCU2D add_1090_4 (.A0(d3[2]), .B0(d4[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[3]), .B1(d4[3]), .C1(GND_net), .D1(GND_net), .CIN(n10876), 
          .COUT(n10877), .S0(d4_71__N_634[2]), .S1(d4_71__N_634[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1090_4.INIT0 = 16'h5666;
    defparam add_1090_4.INIT1 = 16'h5666;
    defparam add_1090_4.INJECT1_0 = "NO";
    defparam add_1090_4.INJECT1_1 = "NO";
    CCU2D add_1090_2 (.A0(d3[0]), .B0(d4[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[1]), .B1(d4[1]), .C1(GND_net), .D1(GND_net), .COUT(n10876), 
          .S1(d4_71__N_634[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1090_2.INIT0 = 16'h7000;
    defparam add_1090_2.INIT1 = 16'h5666;
    defparam add_1090_2.INJECT1_0 = "NO";
    defparam add_1090_2.INJECT1_1 = "NO";
    CCU2D add_1085_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10874), 
          .S0(n5363));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1085_cout.INIT0 = 16'h0000;
    defparam add_1085_cout.INIT1 = 16'h0000;
    defparam add_1085_cout.INJECT1_0 = "NO";
    defparam add_1085_cout.INJECT1_1 = "NO";
    CCU2D add_1085_36 (.A0(d2[34]), .B0(d3[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[35]), .B1(d3[35]), .C1(GND_net), .D1(GND_net), .CIN(n10873), 
          .COUT(n10874), .S0(d3_71__N_562[34]), .S1(d3_71__N_562[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1085_36.INIT0 = 16'h5666;
    defparam add_1085_36.INIT1 = 16'h5666;
    defparam add_1085_36.INJECT1_0 = "NO";
    defparam add_1085_36.INJECT1_1 = "NO";
    CCU2D add_1085_34 (.A0(d2[32]), .B0(d3[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[33]), .B1(d3[33]), .C1(GND_net), .D1(GND_net), .CIN(n10872), 
          .COUT(n10873), .S0(d3_71__N_562[32]), .S1(d3_71__N_562[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1085_34.INIT0 = 16'h5666;
    defparam add_1085_34.INIT1 = 16'h5666;
    defparam add_1085_34.INJECT1_0 = "NO";
    defparam add_1085_34.INJECT1_1 = "NO";
    CCU2D add_1085_32 (.A0(d2[30]), .B0(d3[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[31]), .B1(d3[31]), .C1(GND_net), .D1(GND_net), .CIN(n10871), 
          .COUT(n10872), .S0(d3_71__N_562[30]), .S1(d3_71__N_562[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1085_32.INIT0 = 16'h5666;
    defparam add_1085_32.INIT1 = 16'h5666;
    defparam add_1085_32.INJECT1_0 = "NO";
    defparam add_1085_32.INJECT1_1 = "NO";
    CCU2D add_1085_30 (.A0(d2[28]), .B0(d3[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[29]), .B1(d3[29]), .C1(GND_net), .D1(GND_net), .CIN(n10870), 
          .COUT(n10871), .S0(d3_71__N_562[28]), .S1(d3_71__N_562[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1085_30.INIT0 = 16'h5666;
    defparam add_1085_30.INIT1 = 16'h5666;
    defparam add_1085_30.INJECT1_0 = "NO";
    defparam add_1085_30.INJECT1_1 = "NO";
    CCU2D add_1085_28 (.A0(d2[26]), .B0(d3[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[27]), .B1(d3[27]), .C1(GND_net), .D1(GND_net), .CIN(n10869), 
          .COUT(n10870), .S0(d3_71__N_562[26]), .S1(d3_71__N_562[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1085_28.INIT0 = 16'h5666;
    defparam add_1085_28.INIT1 = 16'h5666;
    defparam add_1085_28.INJECT1_0 = "NO";
    defparam add_1085_28.INJECT1_1 = "NO";
    CCU2D add_1085_26 (.A0(d2[24]), .B0(d3[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[25]), .B1(d3[25]), .C1(GND_net), .D1(GND_net), .CIN(n10868), 
          .COUT(n10869), .S0(d3_71__N_562[24]), .S1(d3_71__N_562[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1085_26.INIT0 = 16'h5666;
    defparam add_1085_26.INIT1 = 16'h5666;
    defparam add_1085_26.INJECT1_0 = "NO";
    defparam add_1085_26.INJECT1_1 = "NO";
    CCU2D add_1085_24 (.A0(d2[22]), .B0(d3[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[23]), .B1(d3[23]), .C1(GND_net), .D1(GND_net), .CIN(n10867), 
          .COUT(n10868), .S0(d3_71__N_562[22]), .S1(d3_71__N_562[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1085_24.INIT0 = 16'h5666;
    defparam add_1085_24.INIT1 = 16'h5666;
    defparam add_1085_24.INJECT1_0 = "NO";
    defparam add_1085_24.INJECT1_1 = "NO";
    CCU2D add_1085_22 (.A0(d2[20]), .B0(d3[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[21]), .B1(d3[21]), .C1(GND_net), .D1(GND_net), .CIN(n10866), 
          .COUT(n10867), .S0(d3_71__N_562[20]), .S1(d3_71__N_562[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1085_22.INIT0 = 16'h5666;
    defparam add_1085_22.INIT1 = 16'h5666;
    defparam add_1085_22.INJECT1_0 = "NO";
    defparam add_1085_22.INJECT1_1 = "NO";
    CCU2D add_1085_20 (.A0(d2[18]), .B0(d3[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[19]), .B1(d3[19]), .C1(GND_net), .D1(GND_net), .CIN(n10865), 
          .COUT(n10866), .S0(d3_71__N_562[18]), .S1(d3_71__N_562[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1085_20.INIT0 = 16'h5666;
    defparam add_1085_20.INIT1 = 16'h5666;
    defparam add_1085_20.INJECT1_0 = "NO";
    defparam add_1085_20.INJECT1_1 = "NO";
    CCU2D add_1085_18 (.A0(d2[16]), .B0(d3[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[17]), .B1(d3[17]), .C1(GND_net), .D1(GND_net), .CIN(n10864), 
          .COUT(n10865), .S0(d3_71__N_562[16]), .S1(d3_71__N_562[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1085_18.INIT0 = 16'h5666;
    defparam add_1085_18.INIT1 = 16'h5666;
    defparam add_1085_18.INJECT1_0 = "NO";
    defparam add_1085_18.INJECT1_1 = "NO";
    CCU2D add_1085_16 (.A0(d2[14]), .B0(d3[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[15]), .B1(d3[15]), .C1(GND_net), .D1(GND_net), .CIN(n10863), 
          .COUT(n10864), .S0(d3_71__N_562[14]), .S1(d3_71__N_562[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1085_16.INIT0 = 16'h5666;
    defparam add_1085_16.INIT1 = 16'h5666;
    defparam add_1085_16.INJECT1_0 = "NO";
    defparam add_1085_16.INJECT1_1 = "NO";
    CCU2D add_1085_14 (.A0(d2[12]), .B0(d3[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[13]), .B1(d3[13]), .C1(GND_net), .D1(GND_net), .CIN(n10862), 
          .COUT(n10863), .S0(d3_71__N_562[12]), .S1(d3_71__N_562[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1085_14.INIT0 = 16'h5666;
    defparam add_1085_14.INIT1 = 16'h5666;
    defparam add_1085_14.INJECT1_0 = "NO";
    defparam add_1085_14.INJECT1_1 = "NO";
    CCU2D add_1085_12 (.A0(d2[10]), .B0(d3[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[11]), .B1(d3[11]), .C1(GND_net), .D1(GND_net), .CIN(n10861), 
          .COUT(n10862), .S0(d3_71__N_562[10]), .S1(d3_71__N_562[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1085_12.INIT0 = 16'h5666;
    defparam add_1085_12.INIT1 = 16'h5666;
    defparam add_1085_12.INJECT1_0 = "NO";
    defparam add_1085_12.INJECT1_1 = "NO";
    CCU2D add_1085_10 (.A0(d2[8]), .B0(d3[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[9]), .B1(d3[9]), .C1(GND_net), .D1(GND_net), .CIN(n10860), 
          .COUT(n10861), .S0(d3_71__N_562[8]), .S1(d3_71__N_562[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1085_10.INIT0 = 16'h5666;
    defparam add_1085_10.INIT1 = 16'h5666;
    defparam add_1085_10.INJECT1_0 = "NO";
    defparam add_1085_10.INJECT1_1 = "NO";
    CCU2D add_1085_8 (.A0(d2[6]), .B0(d3[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[7]), .B1(d3[7]), .C1(GND_net), .D1(GND_net), .CIN(n10859), 
          .COUT(n10860), .S0(d3_71__N_562[6]), .S1(d3_71__N_562[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1085_8.INIT0 = 16'h5666;
    defparam add_1085_8.INIT1 = 16'h5666;
    defparam add_1085_8.INJECT1_0 = "NO";
    defparam add_1085_8.INJECT1_1 = "NO";
    CCU2D add_1085_6 (.A0(d2[4]), .B0(d3[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[5]), .B1(d3[5]), .C1(GND_net), .D1(GND_net), .CIN(n10858), 
          .COUT(n10859), .S0(d3_71__N_562[4]), .S1(d3_71__N_562[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1085_6.INIT0 = 16'h5666;
    defparam add_1085_6.INIT1 = 16'h5666;
    defparam add_1085_6.INJECT1_0 = "NO";
    defparam add_1085_6.INJECT1_1 = "NO";
    CCU2D add_1085_4 (.A0(d2[2]), .B0(d3[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[3]), .B1(d3[3]), .C1(GND_net), .D1(GND_net), .CIN(n10857), 
          .COUT(n10858), .S0(d3_71__N_562[2]), .S1(d3_71__N_562[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1085_4.INIT0 = 16'h5666;
    defparam add_1085_4.INIT1 = 16'h5666;
    defparam add_1085_4.INJECT1_0 = "NO";
    defparam add_1085_4.INJECT1_1 = "NO";
    CCU2D add_1085_2 (.A0(d2[0]), .B0(d3[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[1]), .B1(d3[1]), .C1(GND_net), .D1(GND_net), .COUT(n10857), 
          .S1(d3_71__N_562[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1085_2.INIT0 = 16'h7000;
    defparam add_1085_2.INIT1 = 16'h5666;
    defparam add_1085_2.INJECT1_0 = "NO";
    defparam add_1085_2.INJECT1_1 = "NO";
    CCU2D add_1080_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10855), 
          .S0(n5211));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1080_cout.INIT0 = 16'h0000;
    defparam add_1080_cout.INIT1 = 16'h0000;
    defparam add_1080_cout.INJECT1_0 = "NO";
    defparam add_1080_cout.INJECT1_1 = "NO";
    CCU2D add_1080_36 (.A0(d1[34]), .B0(d2[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[35]), .B1(d2[35]), .C1(GND_net), .D1(GND_net), .CIN(n10854), 
          .COUT(n10855), .S0(d2_71__N_490[34]), .S1(d2_71__N_490[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1080_36.INIT0 = 16'h5666;
    defparam add_1080_36.INIT1 = 16'h5666;
    defparam add_1080_36.INJECT1_0 = "NO";
    defparam add_1080_36.INJECT1_1 = "NO";
    CCU2D add_1080_34 (.A0(d1[32]), .B0(d2[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[33]), .B1(d2[33]), .C1(GND_net), .D1(GND_net), .CIN(n10853), 
          .COUT(n10854), .S0(d2_71__N_490[32]), .S1(d2_71__N_490[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1080_34.INIT0 = 16'h5666;
    defparam add_1080_34.INIT1 = 16'h5666;
    defparam add_1080_34.INJECT1_0 = "NO";
    defparam add_1080_34.INJECT1_1 = "NO";
    CCU2D add_1080_32 (.A0(d1[30]), .B0(d2[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[31]), .B1(d2[31]), .C1(GND_net), .D1(GND_net), .CIN(n10852), 
          .COUT(n10853), .S0(d2_71__N_490[30]), .S1(d2_71__N_490[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1080_32.INIT0 = 16'h5666;
    defparam add_1080_32.INIT1 = 16'h5666;
    defparam add_1080_32.INJECT1_0 = "NO";
    defparam add_1080_32.INJECT1_1 = "NO";
    CCU2D add_1080_30 (.A0(d1[28]), .B0(d2[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[29]), .B1(d2[29]), .C1(GND_net), .D1(GND_net), .CIN(n10851), 
          .COUT(n10852), .S0(d2_71__N_490[28]), .S1(d2_71__N_490[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1080_30.INIT0 = 16'h5666;
    defparam add_1080_30.INIT1 = 16'h5666;
    defparam add_1080_30.INJECT1_0 = "NO";
    defparam add_1080_30.INJECT1_1 = "NO";
    CCU2D add_1080_28 (.A0(d1[26]), .B0(d2[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[27]), .B1(d2[27]), .C1(GND_net), .D1(GND_net), .CIN(n10850), 
          .COUT(n10851), .S0(d2_71__N_490[26]), .S1(d2_71__N_490[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1080_28.INIT0 = 16'h5666;
    defparam add_1080_28.INIT1 = 16'h5666;
    defparam add_1080_28.INJECT1_0 = "NO";
    defparam add_1080_28.INJECT1_1 = "NO";
    CCU2D add_1080_26 (.A0(d1[24]), .B0(d2[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[25]), .B1(d2[25]), .C1(GND_net), .D1(GND_net), .CIN(n10849), 
          .COUT(n10850), .S0(d2_71__N_490[24]), .S1(d2_71__N_490[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1080_26.INIT0 = 16'h5666;
    defparam add_1080_26.INIT1 = 16'h5666;
    defparam add_1080_26.INJECT1_0 = "NO";
    defparam add_1080_26.INJECT1_1 = "NO";
    CCU2D add_1080_24 (.A0(d1[22]), .B0(d2[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[23]), .B1(d2[23]), .C1(GND_net), .D1(GND_net), .CIN(n10848), 
          .COUT(n10849), .S0(d2_71__N_490[22]), .S1(d2_71__N_490[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1080_24.INIT0 = 16'h5666;
    defparam add_1080_24.INIT1 = 16'h5666;
    defparam add_1080_24.INJECT1_0 = "NO";
    defparam add_1080_24.INJECT1_1 = "NO";
    CCU2D add_1080_22 (.A0(d1[20]), .B0(d2[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[21]), .B1(d2[21]), .C1(GND_net), .D1(GND_net), .CIN(n10847), 
          .COUT(n10848), .S0(d2_71__N_490[20]), .S1(d2_71__N_490[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1080_22.INIT0 = 16'h5666;
    defparam add_1080_22.INIT1 = 16'h5666;
    defparam add_1080_22.INJECT1_0 = "NO";
    defparam add_1080_22.INJECT1_1 = "NO";
    CCU2D add_1080_20 (.A0(d1[18]), .B0(d2[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[19]), .B1(d2[19]), .C1(GND_net), .D1(GND_net), .CIN(n10846), 
          .COUT(n10847), .S0(d2_71__N_490[18]), .S1(d2_71__N_490[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1080_20.INIT0 = 16'h5666;
    defparam add_1080_20.INIT1 = 16'h5666;
    defparam add_1080_20.INJECT1_0 = "NO";
    defparam add_1080_20.INJECT1_1 = "NO";
    CCU2D add_1080_18 (.A0(d1[16]), .B0(d2[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[17]), .B1(d2[17]), .C1(GND_net), .D1(GND_net), .CIN(n10845), 
          .COUT(n10846), .S0(d2_71__N_490[16]), .S1(d2_71__N_490[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1080_18.INIT0 = 16'h5666;
    defparam add_1080_18.INIT1 = 16'h5666;
    defparam add_1080_18.INJECT1_0 = "NO";
    defparam add_1080_18.INJECT1_1 = "NO";
    CCU2D add_1080_16 (.A0(d1[14]), .B0(d2[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[15]), .B1(d2[15]), .C1(GND_net), .D1(GND_net), .CIN(n10844), 
          .COUT(n10845), .S0(d2_71__N_490[14]), .S1(d2_71__N_490[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1080_16.INIT0 = 16'h5666;
    defparam add_1080_16.INIT1 = 16'h5666;
    defparam add_1080_16.INJECT1_0 = "NO";
    defparam add_1080_16.INJECT1_1 = "NO";
    CCU2D add_1080_14 (.A0(d1[12]), .B0(d2[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[13]), .B1(d2[13]), .C1(GND_net), .D1(GND_net), .CIN(n10843), 
          .COUT(n10844), .S0(d2_71__N_490[12]), .S1(d2_71__N_490[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1080_14.INIT0 = 16'h5666;
    defparam add_1080_14.INIT1 = 16'h5666;
    defparam add_1080_14.INJECT1_0 = "NO";
    defparam add_1080_14.INJECT1_1 = "NO";
    CCU2D add_1080_12 (.A0(d1[10]), .B0(d2[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[11]), .B1(d2[11]), .C1(GND_net), .D1(GND_net), .CIN(n10842), 
          .COUT(n10843), .S0(d2_71__N_490[10]), .S1(d2_71__N_490[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1080_12.INIT0 = 16'h5666;
    defparam add_1080_12.INIT1 = 16'h5666;
    defparam add_1080_12.INJECT1_0 = "NO";
    defparam add_1080_12.INJECT1_1 = "NO";
    CCU2D add_1080_10 (.A0(d1[8]), .B0(d2[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[9]), .B1(d2[9]), .C1(GND_net), .D1(GND_net), .CIN(n10841), 
          .COUT(n10842), .S0(d2_71__N_490[8]), .S1(d2_71__N_490[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1080_10.INIT0 = 16'h5666;
    defparam add_1080_10.INIT1 = 16'h5666;
    defparam add_1080_10.INJECT1_0 = "NO";
    defparam add_1080_10.INJECT1_1 = "NO";
    CCU2D add_1080_8 (.A0(d1[6]), .B0(d2[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[7]), .B1(d2[7]), .C1(GND_net), .D1(GND_net), .CIN(n10840), 
          .COUT(n10841), .S0(d2_71__N_490[6]), .S1(d2_71__N_490[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1080_8.INIT0 = 16'h5666;
    defparam add_1080_8.INIT1 = 16'h5666;
    defparam add_1080_8.INJECT1_0 = "NO";
    defparam add_1080_8.INJECT1_1 = "NO";
    CCU2D add_1080_6 (.A0(d1[4]), .B0(d2[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[5]), .B1(d2[5]), .C1(GND_net), .D1(GND_net), .CIN(n10839), 
          .COUT(n10840), .S0(d2_71__N_490[4]), .S1(d2_71__N_490[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1080_6.INIT0 = 16'h5666;
    defparam add_1080_6.INIT1 = 16'h5666;
    defparam add_1080_6.INJECT1_0 = "NO";
    defparam add_1080_6.INJECT1_1 = "NO";
    CCU2D add_1080_4 (.A0(d1[2]), .B0(d2[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[3]), .B1(d2[3]), .C1(GND_net), .D1(GND_net), .CIN(n10838), 
          .COUT(n10839), .S0(d2_71__N_490[2]), .S1(d2_71__N_490[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1080_4.INIT0 = 16'h5666;
    defparam add_1080_4.INIT1 = 16'h5666;
    defparam add_1080_4.INJECT1_0 = "NO";
    defparam add_1080_4.INJECT1_1 = "NO";
    CCU2D add_1080_2 (.A0(d1[0]), .B0(d2[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[1]), .B1(d2[1]), .C1(GND_net), .D1(GND_net), .COUT(n10838), 
          .S1(d2_71__N_490[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1080_2.INIT0 = 16'h7000;
    defparam add_1080_2.INIT1 = 16'h5666;
    defparam add_1080_2.INJECT1_0 = "NO";
    defparam add_1080_2.INJECT1_1 = "NO";
    CCU2D add_1075_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10798), 
          .S0(n5059));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1075_cout.INIT0 = 16'h0000;
    defparam add_1075_cout.INIT1 = 16'h0000;
    defparam add_1075_cout.INJECT1_0 = "NO";
    defparam add_1075_cout.INJECT1_1 = "NO";
    CCU2D add_1075_36 (.A0(MixerOutCos[11]), .B0(d1[34]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[35]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10797), .COUT(n10798), .S0(d1_71__N_418[34]), 
          .S1(d1_71__N_418[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1075_36.INIT0 = 16'h5666;
    defparam add_1075_36.INIT1 = 16'h5666;
    defparam add_1075_36.INJECT1_0 = "NO";
    defparam add_1075_36.INJECT1_1 = "NO";
    CCU2D add_1075_34 (.A0(MixerOutCos[11]), .B0(d1[32]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[33]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10796), .COUT(n10797), .S0(d1_71__N_418[32]), 
          .S1(d1_71__N_418[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1075_34.INIT0 = 16'h5666;
    defparam add_1075_34.INIT1 = 16'h5666;
    defparam add_1075_34.INJECT1_0 = "NO";
    defparam add_1075_34.INJECT1_1 = "NO";
    CCU2D add_1075_32 (.A0(MixerOutCos[11]), .B0(d1[30]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10795), .COUT(n10796), .S0(d1_71__N_418[30]), 
          .S1(d1_71__N_418[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1075_32.INIT0 = 16'h5666;
    defparam add_1075_32.INIT1 = 16'h5666;
    defparam add_1075_32.INJECT1_0 = "NO";
    defparam add_1075_32.INJECT1_1 = "NO";
    CCU2D add_1075_30 (.A0(MixerOutCos[11]), .B0(d1[28]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10794), .COUT(n10795), .S0(d1_71__N_418[28]), 
          .S1(d1_71__N_418[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1075_30.INIT0 = 16'h5666;
    defparam add_1075_30.INIT1 = 16'h5666;
    defparam add_1075_30.INJECT1_0 = "NO";
    defparam add_1075_30.INJECT1_1 = "NO";
    CCU2D add_1075_28 (.A0(MixerOutCos[11]), .B0(d1[26]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10793), .COUT(n10794), .S0(d1_71__N_418[26]), 
          .S1(d1_71__N_418[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1075_28.INIT0 = 16'h5666;
    defparam add_1075_28.INIT1 = 16'h5666;
    defparam add_1075_28.INJECT1_0 = "NO";
    defparam add_1075_28.INJECT1_1 = "NO";
    CCU2D add_1075_26 (.A0(MixerOutCos[11]), .B0(d1[24]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10792), .COUT(n10793), .S0(d1_71__N_418[24]), 
          .S1(d1_71__N_418[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1075_26.INIT0 = 16'h5666;
    defparam add_1075_26.INIT1 = 16'h5666;
    defparam add_1075_26.INJECT1_0 = "NO";
    defparam add_1075_26.INJECT1_1 = "NO";
    CCU2D add_1075_24 (.A0(MixerOutCos[11]), .B0(d1[22]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10791), .COUT(n10792), .S0(d1_71__N_418[22]), 
          .S1(d1_71__N_418[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1075_24.INIT0 = 16'h5666;
    defparam add_1075_24.INIT1 = 16'h5666;
    defparam add_1075_24.INJECT1_0 = "NO";
    defparam add_1075_24.INJECT1_1 = "NO";
    CCU2D add_1075_22 (.A0(MixerOutCos[11]), .B0(d1[20]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10790), .COUT(n10791), .S0(d1_71__N_418[20]), 
          .S1(d1_71__N_418[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1075_22.INIT0 = 16'h5666;
    defparam add_1075_22.INIT1 = 16'h5666;
    defparam add_1075_22.INJECT1_0 = "NO";
    defparam add_1075_22.INJECT1_1 = "NO";
    CCU2D add_1075_20 (.A0(MixerOutCos[11]), .B0(d1[18]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10789), .COUT(n10790), .S0(d1_71__N_418[18]), 
          .S1(d1_71__N_418[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1075_20.INIT0 = 16'h5666;
    defparam add_1075_20.INIT1 = 16'h5666;
    defparam add_1075_20.INJECT1_0 = "NO";
    defparam add_1075_20.INJECT1_1 = "NO";
    CCU2D add_1075_18 (.A0(MixerOutCos[11]), .B0(d1[16]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10788), .COUT(n10789), .S0(d1_71__N_418[16]), 
          .S1(d1_71__N_418[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1075_18.INIT0 = 16'h5666;
    defparam add_1075_18.INIT1 = 16'h5666;
    defparam add_1075_18.INJECT1_0 = "NO";
    defparam add_1075_18.INJECT1_1 = "NO";
    CCU2D add_1075_16 (.A0(MixerOutCos[11]), .B0(d1[14]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10787), .COUT(n10788), .S0(d1_71__N_418[14]), 
          .S1(d1_71__N_418[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1075_16.INIT0 = 16'h5666;
    defparam add_1075_16.INIT1 = 16'h5666;
    defparam add_1075_16.INJECT1_0 = "NO";
    defparam add_1075_16.INJECT1_1 = "NO";
    CCU2D add_1075_14 (.A0(MixerOutCos[11]), .B0(d1[12]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10786), .COUT(n10787), .S0(d1_71__N_418[12]), 
          .S1(d1_71__N_418[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1075_14.INIT0 = 16'h5666;
    defparam add_1075_14.INIT1 = 16'h5666;
    defparam add_1075_14.INJECT1_0 = "NO";
    defparam add_1075_14.INJECT1_1 = "NO";
    CCU2D add_1075_12 (.A0(MixerOutCos[10]), .B0(d1[10]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10785), .COUT(n10786), .S0(d1_71__N_418[10]), 
          .S1(d1_71__N_418[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1075_12.INIT0 = 16'h5666;
    defparam add_1075_12.INIT1 = 16'h5666;
    defparam add_1075_12.INJECT1_0 = "NO";
    defparam add_1075_12.INJECT1_1 = "NO";
    CCU2D add_1075_10 (.A0(MixerOutCos[8]), .B0(d1[8]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[9]), .B1(d1[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10784), .COUT(n10785), .S0(d1_71__N_418[8]), 
          .S1(d1_71__N_418[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1075_10.INIT0 = 16'h5666;
    defparam add_1075_10.INIT1 = 16'h5666;
    defparam add_1075_10.INJECT1_0 = "NO";
    defparam add_1075_10.INJECT1_1 = "NO";
    CCU2D add_1075_8 (.A0(MixerOutCos[6]), .B0(d1[6]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutCos[7]), .B1(d1[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10783), .COUT(n10784), .S0(d1_71__N_418[6]), .S1(d1_71__N_418[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1075_8.INIT0 = 16'h5666;
    defparam add_1075_8.INIT1 = 16'h5666;
    defparam add_1075_8.INJECT1_0 = "NO";
    defparam add_1075_8.INJECT1_1 = "NO";
    CCU2D add_1075_6 (.A0(MixerOutCos[4]), .B0(d1[4]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutCos[5]), .B1(d1[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10782), .COUT(n10783), .S0(d1_71__N_418[4]), .S1(d1_71__N_418[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1075_6.INIT0 = 16'h5666;
    defparam add_1075_6.INIT1 = 16'h5666;
    defparam add_1075_6.INJECT1_0 = "NO";
    defparam add_1075_6.INJECT1_1 = "NO";
    CCU2D add_1075_4 (.A0(MixerOutCos[2]), .B0(d1[2]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutCos[3]), .B1(d1[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10781), .COUT(n10782), .S0(d1_71__N_418[2]), .S1(d1_71__N_418[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1075_4.INIT0 = 16'h5666;
    defparam add_1075_4.INIT1 = 16'h5666;
    defparam add_1075_4.INJECT1_0 = "NO";
    defparam add_1075_4.INJECT1_1 = "NO";
    CCU2D add_1075_2 (.A0(MixerOutCos[0]), .B0(d1[0]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutCos[1]), .B1(d1[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n10781), .S1(d1_71__N_418[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1075_2.INIT0 = 16'h7000;
    defparam add_1075_2.INIT1 = 16'h5666;
    defparam add_1075_2.INJECT1_0 = "NO";
    defparam add_1075_2.INJECT1_1 = "NO";
    CCU2D add_1130_37 (.A0(d9[35]), .B0(d_d9[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11452), 
          .S1(n6731));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1130_37.INIT0 = 16'h5999;
    defparam add_1130_37.INIT1 = 16'h0000;
    defparam add_1130_37.INJECT1_0 = "NO";
    defparam add_1130_37.INJECT1_1 = "NO";
    CCU2D add_1130_35 (.A0(d9[33]), .B0(d_d9[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[34]), .B1(d_d9[34]), .C1(GND_net), .D1(GND_net), .CIN(n11451), 
          .COUT(n11452));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1130_35.INIT0 = 16'h5999;
    defparam add_1130_35.INIT1 = 16'h5999;
    defparam add_1130_35.INJECT1_0 = "NO";
    defparam add_1130_35.INJECT1_1 = "NO";
    CCU2D add_1130_33 (.A0(d9[31]), .B0(d_d9[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[32]), .B1(d_d9[32]), .C1(GND_net), .D1(GND_net), .CIN(n11450), 
          .COUT(n11451));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1130_33.INIT0 = 16'h5999;
    defparam add_1130_33.INIT1 = 16'h5999;
    defparam add_1130_33.INJECT1_0 = "NO";
    defparam add_1130_33.INJECT1_1 = "NO";
    CCU2D add_1130_31 (.A0(d9[29]), .B0(d_d9[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[30]), .B1(d_d9[30]), .C1(GND_net), .D1(GND_net), .CIN(n11449), 
          .COUT(n11450));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1130_31.INIT0 = 16'h5999;
    defparam add_1130_31.INIT1 = 16'h5999;
    defparam add_1130_31.INJECT1_0 = "NO";
    defparam add_1130_31.INJECT1_1 = "NO";
    CCU2D add_1130_29 (.A0(d9[27]), .B0(d_d9[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[28]), .B1(d_d9[28]), .C1(GND_net), .D1(GND_net), .CIN(n11448), 
          .COUT(n11449));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1130_29.INIT0 = 16'h5999;
    defparam add_1130_29.INIT1 = 16'h5999;
    defparam add_1130_29.INJECT1_0 = "NO";
    defparam add_1130_29.INJECT1_1 = "NO";
    CCU2D add_1130_27 (.A0(d9[25]), .B0(d_d9[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[26]), .B1(d_d9[26]), .C1(GND_net), .D1(GND_net), .CIN(n11447), 
          .COUT(n11448));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1130_27.INIT0 = 16'h5999;
    defparam add_1130_27.INIT1 = 16'h5999;
    defparam add_1130_27.INJECT1_0 = "NO";
    defparam add_1130_27.INJECT1_1 = "NO";
    CCU2D add_1130_25 (.A0(d9[23]), .B0(d_d9[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[24]), .B1(d_d9[24]), .C1(GND_net), .D1(GND_net), .CIN(n11446), 
          .COUT(n11447));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1130_25.INIT0 = 16'h5999;
    defparam add_1130_25.INIT1 = 16'h5999;
    defparam add_1130_25.INJECT1_0 = "NO";
    defparam add_1130_25.INJECT1_1 = "NO";
    CCU2D add_1130_23 (.A0(d9[21]), .B0(d_d9[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[22]), .B1(d_d9[22]), .C1(GND_net), .D1(GND_net), .CIN(n11445), 
          .COUT(n11446));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1130_23.INIT0 = 16'h5999;
    defparam add_1130_23.INIT1 = 16'h5999;
    defparam add_1130_23.INJECT1_0 = "NO";
    defparam add_1130_23.INJECT1_1 = "NO";
    CCU2D add_1130_21 (.A0(d9[19]), .B0(d_d9[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[20]), .B1(d_d9[20]), .C1(GND_net), .D1(GND_net), .CIN(n11444), 
          .COUT(n11445));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1130_21.INIT0 = 16'h5999;
    defparam add_1130_21.INIT1 = 16'h5999;
    defparam add_1130_21.INJECT1_0 = "NO";
    defparam add_1130_21.INJECT1_1 = "NO";
    CCU2D add_1130_19 (.A0(d9[17]), .B0(d_d9[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[18]), .B1(d_d9[18]), .C1(GND_net), .D1(GND_net), .CIN(n11443), 
          .COUT(n11444));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1130_19.INIT0 = 16'h5999;
    defparam add_1130_19.INIT1 = 16'h5999;
    defparam add_1130_19.INJECT1_0 = "NO";
    defparam add_1130_19.INJECT1_1 = "NO";
    CCU2D add_1130_17 (.A0(d9[15]), .B0(d_d9[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[16]), .B1(d_d9[16]), .C1(GND_net), .D1(GND_net), .CIN(n11442), 
          .COUT(n11443));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1130_17.INIT0 = 16'h5999;
    defparam add_1130_17.INIT1 = 16'h5999;
    defparam add_1130_17.INJECT1_0 = "NO";
    defparam add_1130_17.INJECT1_1 = "NO";
    CCU2D add_1130_15 (.A0(d9[13]), .B0(d_d9[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[14]), .B1(d_d9[14]), .C1(GND_net), .D1(GND_net), .CIN(n11441), 
          .COUT(n11442));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1130_15.INIT0 = 16'h5999;
    defparam add_1130_15.INIT1 = 16'h5999;
    defparam add_1130_15.INJECT1_0 = "NO";
    defparam add_1130_15.INJECT1_1 = "NO";
    CCU2D add_1130_13 (.A0(d9[11]), .B0(d_d9[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[12]), .B1(d_d9[12]), .C1(GND_net), .D1(GND_net), .CIN(n11440), 
          .COUT(n11441));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1130_13.INIT0 = 16'h5999;
    defparam add_1130_13.INIT1 = 16'h5999;
    defparam add_1130_13.INJECT1_0 = "NO";
    defparam add_1130_13.INJECT1_1 = "NO";
    CCU2D add_1130_11 (.A0(d9[9]), .B0(d_d9[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[10]), .B1(d_d9[10]), .C1(GND_net), .D1(GND_net), .CIN(n11439), 
          .COUT(n11440));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1130_11.INIT0 = 16'h5999;
    defparam add_1130_11.INIT1 = 16'h5999;
    defparam add_1130_11.INJECT1_0 = "NO";
    defparam add_1130_11.INJECT1_1 = "NO";
    CCU2D add_1130_9 (.A0(d9[7]), .B0(d_d9[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[8]), .B1(d_d9[8]), .C1(GND_net), .D1(GND_net), .CIN(n11438), 
          .COUT(n11439));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1130_9.INIT0 = 16'h5999;
    defparam add_1130_9.INIT1 = 16'h5999;
    defparam add_1130_9.INJECT1_0 = "NO";
    defparam add_1130_9.INJECT1_1 = "NO";
    CCU2D add_1130_7 (.A0(d9[5]), .B0(d_d9[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[6]), .B1(d_d9[6]), .C1(GND_net), .D1(GND_net), .CIN(n11437), 
          .COUT(n11438));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1130_7.INIT0 = 16'h5999;
    defparam add_1130_7.INIT1 = 16'h5999;
    defparam add_1130_7.INJECT1_0 = "NO";
    defparam add_1130_7.INJECT1_1 = "NO";
    CCU2D add_1130_5 (.A0(d9[3]), .B0(d_d9[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[4]), .B1(d_d9[4]), .C1(GND_net), .D1(GND_net), .CIN(n11436), 
          .COUT(n11437));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1130_5.INIT0 = 16'h5999;
    defparam add_1130_5.INIT1 = 16'h5999;
    defparam add_1130_5.INJECT1_0 = "NO";
    defparam add_1130_5.INJECT1_1 = "NO";
    CCU2D add_1130_3 (.A0(d9[1]), .B0(d_d9[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[2]), .B1(d_d9[2]), .C1(GND_net), .D1(GND_net), .CIN(n11435), 
          .COUT(n11436));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1130_3.INIT0 = 16'h5999;
    defparam add_1130_3.INIT1 = 16'h5999;
    defparam add_1130_3.INJECT1_0 = "NO";
    defparam add_1130_3.INJECT1_1 = "NO";
    CCU2D add_1130_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d9[0]), .B1(d_d9[0]), .C1(GND_net), .D1(GND_net), .COUT(n11435));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1130_1.INIT0 = 16'h0000;
    defparam add_1130_1.INIT1 = 16'h5999;
    defparam add_1130_1.INJECT1_0 = "NO";
    defparam add_1130_1.INJECT1_1 = "NO";
    CCU2D add_1125_37 (.A0(d8[35]), .B0(d_d8[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11434), 
          .S0(d9_71__N_1675[35]), .S1(n6579));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1125_37.INIT0 = 16'h5999;
    defparam add_1125_37.INIT1 = 16'h0000;
    defparam add_1125_37.INJECT1_0 = "NO";
    defparam add_1125_37.INJECT1_1 = "NO";
    CCU2D add_1125_35 (.A0(d8[33]), .B0(d_d8[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[34]), .B1(d_d8[34]), .C1(GND_net), .D1(GND_net), .CIN(n11433), 
          .COUT(n11434), .S0(d9_71__N_1675[33]), .S1(d9_71__N_1675[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1125_35.INIT0 = 16'h5999;
    defparam add_1125_35.INIT1 = 16'h5999;
    defparam add_1125_35.INJECT1_0 = "NO";
    defparam add_1125_35.INJECT1_1 = "NO";
    CCU2D add_1125_33 (.A0(d8[31]), .B0(d_d8[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[32]), .B1(d_d8[32]), .C1(GND_net), .D1(GND_net), .CIN(n11432), 
          .COUT(n11433), .S0(d9_71__N_1675[31]), .S1(d9_71__N_1675[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1125_33.INIT0 = 16'h5999;
    defparam add_1125_33.INIT1 = 16'h5999;
    defparam add_1125_33.INJECT1_0 = "NO";
    defparam add_1125_33.INJECT1_1 = "NO";
    CCU2D add_1125_31 (.A0(d8[29]), .B0(d_d8[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[30]), .B1(d_d8[30]), .C1(GND_net), .D1(GND_net), .CIN(n11431), 
          .COUT(n11432), .S0(d9_71__N_1675[29]), .S1(d9_71__N_1675[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1125_31.INIT0 = 16'h5999;
    defparam add_1125_31.INIT1 = 16'h5999;
    defparam add_1125_31.INJECT1_0 = "NO";
    defparam add_1125_31.INJECT1_1 = "NO";
    CCU2D add_1125_29 (.A0(d8[27]), .B0(d_d8[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[28]), .B1(d_d8[28]), .C1(GND_net), .D1(GND_net), .CIN(n11430), 
          .COUT(n11431), .S0(d9_71__N_1675[27]), .S1(d9_71__N_1675[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1125_29.INIT0 = 16'h5999;
    defparam add_1125_29.INIT1 = 16'h5999;
    defparam add_1125_29.INJECT1_0 = "NO";
    defparam add_1125_29.INJECT1_1 = "NO";
    CCU2D add_1125_27 (.A0(d8[25]), .B0(d_d8[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[26]), .B1(d_d8[26]), .C1(GND_net), .D1(GND_net), .CIN(n11429), 
          .COUT(n11430), .S0(d9_71__N_1675[25]), .S1(d9_71__N_1675[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1125_27.INIT0 = 16'h5999;
    defparam add_1125_27.INIT1 = 16'h5999;
    defparam add_1125_27.INJECT1_0 = "NO";
    defparam add_1125_27.INJECT1_1 = "NO";
    CCU2D add_1125_25 (.A0(d8[23]), .B0(d_d8[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[24]), .B1(d_d8[24]), .C1(GND_net), .D1(GND_net), .CIN(n11428), 
          .COUT(n11429), .S0(d9_71__N_1675[23]), .S1(d9_71__N_1675[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1125_25.INIT0 = 16'h5999;
    defparam add_1125_25.INIT1 = 16'h5999;
    defparam add_1125_25.INJECT1_0 = "NO";
    defparam add_1125_25.INJECT1_1 = "NO";
    CCU2D add_1125_23 (.A0(d8[21]), .B0(d_d8[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[22]), .B1(d_d8[22]), .C1(GND_net), .D1(GND_net), .CIN(n11427), 
          .COUT(n11428), .S0(d9_71__N_1675[21]), .S1(d9_71__N_1675[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1125_23.INIT0 = 16'h5999;
    defparam add_1125_23.INIT1 = 16'h5999;
    defparam add_1125_23.INJECT1_0 = "NO";
    defparam add_1125_23.INJECT1_1 = "NO";
    CCU2D add_1125_21 (.A0(d8[19]), .B0(d_d8[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[20]), .B1(d_d8[20]), .C1(GND_net), .D1(GND_net), .CIN(n11426), 
          .COUT(n11427), .S0(d9_71__N_1675[19]), .S1(d9_71__N_1675[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1125_21.INIT0 = 16'h5999;
    defparam add_1125_21.INIT1 = 16'h5999;
    defparam add_1125_21.INJECT1_0 = "NO";
    defparam add_1125_21.INJECT1_1 = "NO";
    CCU2D add_1125_19 (.A0(d8[17]), .B0(d_d8[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[18]), .B1(d_d8[18]), .C1(GND_net), .D1(GND_net), .CIN(n11425), 
          .COUT(n11426), .S0(d9_71__N_1675[17]), .S1(d9_71__N_1675[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1125_19.INIT0 = 16'h5999;
    defparam add_1125_19.INIT1 = 16'h5999;
    defparam add_1125_19.INJECT1_0 = "NO";
    defparam add_1125_19.INJECT1_1 = "NO";
    CCU2D add_1125_17 (.A0(d8[15]), .B0(d_d8[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[16]), .B1(d_d8[16]), .C1(GND_net), .D1(GND_net), .CIN(n11424), 
          .COUT(n11425), .S0(d9_71__N_1675[15]), .S1(d9_71__N_1675[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1125_17.INIT0 = 16'h5999;
    defparam add_1125_17.INIT1 = 16'h5999;
    defparam add_1125_17.INJECT1_0 = "NO";
    defparam add_1125_17.INJECT1_1 = "NO";
    CCU2D add_1125_15 (.A0(d8[13]), .B0(d_d8[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[14]), .B1(d_d8[14]), .C1(GND_net), .D1(GND_net), .CIN(n11423), 
          .COUT(n11424), .S0(d9_71__N_1675[13]), .S1(d9_71__N_1675[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1125_15.INIT0 = 16'h5999;
    defparam add_1125_15.INIT1 = 16'h5999;
    defparam add_1125_15.INJECT1_0 = "NO";
    defparam add_1125_15.INJECT1_1 = "NO";
    CCU2D add_1125_13 (.A0(d8[11]), .B0(d_d8[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[12]), .B1(d_d8[12]), .C1(GND_net), .D1(GND_net), .CIN(n11422), 
          .COUT(n11423), .S0(d9_71__N_1675[11]), .S1(d9_71__N_1675[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1125_13.INIT0 = 16'h5999;
    defparam add_1125_13.INIT1 = 16'h5999;
    defparam add_1125_13.INJECT1_0 = "NO";
    defparam add_1125_13.INJECT1_1 = "NO";
    CCU2D add_1125_11 (.A0(d8[9]), .B0(d_d8[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[10]), .B1(d_d8[10]), .C1(GND_net), .D1(GND_net), .CIN(n11421), 
          .COUT(n11422), .S0(d9_71__N_1675[9]), .S1(d9_71__N_1675[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1125_11.INIT0 = 16'h5999;
    defparam add_1125_11.INIT1 = 16'h5999;
    defparam add_1125_11.INJECT1_0 = "NO";
    defparam add_1125_11.INJECT1_1 = "NO";
    CCU2D add_1125_9 (.A0(d8[7]), .B0(d_d8[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[8]), .B1(d_d8[8]), .C1(GND_net), .D1(GND_net), .CIN(n11420), 
          .COUT(n11421), .S0(d9_71__N_1675[7]), .S1(d9_71__N_1675[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1125_9.INIT0 = 16'h5999;
    defparam add_1125_9.INIT1 = 16'h5999;
    defparam add_1125_9.INJECT1_0 = "NO";
    defparam add_1125_9.INJECT1_1 = "NO";
    CCU2D add_1125_7 (.A0(d8[5]), .B0(d_d8[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[6]), .B1(d_d8[6]), .C1(GND_net), .D1(GND_net), .CIN(n11419), 
          .COUT(n11420), .S0(d9_71__N_1675[5]), .S1(d9_71__N_1675[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1125_7.INIT0 = 16'h5999;
    defparam add_1125_7.INIT1 = 16'h5999;
    defparam add_1125_7.INJECT1_0 = "NO";
    defparam add_1125_7.INJECT1_1 = "NO";
    CCU2D add_1125_5 (.A0(d8[3]), .B0(d_d8[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[4]), .B1(d_d8[4]), .C1(GND_net), .D1(GND_net), .CIN(n11418), 
          .COUT(n11419), .S0(d9_71__N_1675[3]), .S1(d9_71__N_1675[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1125_5.INIT0 = 16'h5999;
    defparam add_1125_5.INIT1 = 16'h5999;
    defparam add_1125_5.INJECT1_0 = "NO";
    defparam add_1125_5.INJECT1_1 = "NO";
    CCU2D add_1125_3 (.A0(d8[1]), .B0(d_d8[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[2]), .B1(d_d8[2]), .C1(GND_net), .D1(GND_net), .CIN(n11417), 
          .COUT(n11418), .S0(d9_71__N_1675[1]), .S1(d9_71__N_1675[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1125_3.INIT0 = 16'h5999;
    defparam add_1125_3.INIT1 = 16'h5999;
    defparam add_1125_3.INJECT1_0 = "NO";
    defparam add_1125_3.INJECT1_1 = "NO";
    CCU2D add_1125_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d8[0]), .B1(d_d8[0]), .C1(GND_net), .D1(GND_net), .COUT(n11417), 
          .S1(d9_71__N_1675[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1125_1.INIT0 = 16'h0000;
    defparam add_1125_1.INIT1 = 16'h5999;
    defparam add_1125_1.INJECT1_0 = "NO";
    defparam add_1125_1.INJECT1_1 = "NO";
    CCU2D add_1120_37 (.A0(d7[35]), .B0(d_d7[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11416), 
          .S0(d8_71__N_1603[35]), .S1(n6427));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1120_37.INIT0 = 16'h5999;
    defparam add_1120_37.INIT1 = 16'h0000;
    defparam add_1120_37.INJECT1_0 = "NO";
    defparam add_1120_37.INJECT1_1 = "NO";
    CCU2D add_1120_35 (.A0(d7[33]), .B0(d_d7[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[34]), .B1(d_d7[34]), .C1(GND_net), .D1(GND_net), .CIN(n11415), 
          .COUT(n11416), .S0(d8_71__N_1603[33]), .S1(d8_71__N_1603[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1120_35.INIT0 = 16'h5999;
    defparam add_1120_35.INIT1 = 16'h5999;
    defparam add_1120_35.INJECT1_0 = "NO";
    defparam add_1120_35.INJECT1_1 = "NO";
    CCU2D add_1120_33 (.A0(d7[31]), .B0(d_d7[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[32]), .B1(d_d7[32]), .C1(GND_net), .D1(GND_net), .CIN(n11414), 
          .COUT(n11415), .S0(d8_71__N_1603[31]), .S1(d8_71__N_1603[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1120_33.INIT0 = 16'h5999;
    defparam add_1120_33.INIT1 = 16'h5999;
    defparam add_1120_33.INJECT1_0 = "NO";
    defparam add_1120_33.INJECT1_1 = "NO";
    CCU2D add_1120_31 (.A0(d7[29]), .B0(d_d7[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[30]), .B1(d_d7[30]), .C1(GND_net), .D1(GND_net), .CIN(n11413), 
          .COUT(n11414), .S0(d8_71__N_1603[29]), .S1(d8_71__N_1603[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1120_31.INIT0 = 16'h5999;
    defparam add_1120_31.INIT1 = 16'h5999;
    defparam add_1120_31.INJECT1_0 = "NO";
    defparam add_1120_31.INJECT1_1 = "NO";
    CCU2D add_1120_29 (.A0(d7[27]), .B0(d_d7[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[28]), .B1(d_d7[28]), .C1(GND_net), .D1(GND_net), .CIN(n11412), 
          .COUT(n11413), .S0(d8_71__N_1603[27]), .S1(d8_71__N_1603[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1120_29.INIT0 = 16'h5999;
    defparam add_1120_29.INIT1 = 16'h5999;
    defparam add_1120_29.INJECT1_0 = "NO";
    defparam add_1120_29.INJECT1_1 = "NO";
    CCU2D add_1120_27 (.A0(d7[25]), .B0(d_d7[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[26]), .B1(d_d7[26]), .C1(GND_net), .D1(GND_net), .CIN(n11411), 
          .COUT(n11412), .S0(d8_71__N_1603[25]), .S1(d8_71__N_1603[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1120_27.INIT0 = 16'h5999;
    defparam add_1120_27.INIT1 = 16'h5999;
    defparam add_1120_27.INJECT1_0 = "NO";
    defparam add_1120_27.INJECT1_1 = "NO";
    CCU2D add_1120_25 (.A0(d7[23]), .B0(d_d7[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[24]), .B1(d_d7[24]), .C1(GND_net), .D1(GND_net), .CIN(n11410), 
          .COUT(n11411), .S0(d8_71__N_1603[23]), .S1(d8_71__N_1603[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1120_25.INIT0 = 16'h5999;
    defparam add_1120_25.INIT1 = 16'h5999;
    defparam add_1120_25.INJECT1_0 = "NO";
    defparam add_1120_25.INJECT1_1 = "NO";
    CCU2D add_1120_23 (.A0(d7[21]), .B0(d_d7[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[22]), .B1(d_d7[22]), .C1(GND_net), .D1(GND_net), .CIN(n11409), 
          .COUT(n11410), .S0(d8_71__N_1603[21]), .S1(d8_71__N_1603[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1120_23.INIT0 = 16'h5999;
    defparam add_1120_23.INIT1 = 16'h5999;
    defparam add_1120_23.INJECT1_0 = "NO";
    defparam add_1120_23.INJECT1_1 = "NO";
    CCU2D add_1120_21 (.A0(d7[19]), .B0(d_d7[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[20]), .B1(d_d7[20]), .C1(GND_net), .D1(GND_net), .CIN(n11408), 
          .COUT(n11409), .S0(d8_71__N_1603[19]), .S1(d8_71__N_1603[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1120_21.INIT0 = 16'h5999;
    defparam add_1120_21.INIT1 = 16'h5999;
    defparam add_1120_21.INJECT1_0 = "NO";
    defparam add_1120_21.INJECT1_1 = "NO";
    CCU2D add_1120_19 (.A0(d7[17]), .B0(d_d7[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[18]), .B1(d_d7[18]), .C1(GND_net), .D1(GND_net), .CIN(n11407), 
          .COUT(n11408), .S0(d8_71__N_1603[17]), .S1(d8_71__N_1603[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1120_19.INIT0 = 16'h5999;
    defparam add_1120_19.INIT1 = 16'h5999;
    defparam add_1120_19.INJECT1_0 = "NO";
    defparam add_1120_19.INJECT1_1 = "NO";
    CCU2D add_1120_17 (.A0(d7[15]), .B0(d_d7[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[16]), .B1(d_d7[16]), .C1(GND_net), .D1(GND_net), .CIN(n11406), 
          .COUT(n11407), .S0(d8_71__N_1603[15]), .S1(d8_71__N_1603[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1120_17.INIT0 = 16'h5999;
    defparam add_1120_17.INIT1 = 16'h5999;
    defparam add_1120_17.INJECT1_0 = "NO";
    defparam add_1120_17.INJECT1_1 = "NO";
    CCU2D add_1120_15 (.A0(d7[13]), .B0(d_d7[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[14]), .B1(d_d7[14]), .C1(GND_net), .D1(GND_net), .CIN(n11405), 
          .COUT(n11406), .S0(d8_71__N_1603[13]), .S1(d8_71__N_1603[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1120_15.INIT0 = 16'h5999;
    defparam add_1120_15.INIT1 = 16'h5999;
    defparam add_1120_15.INJECT1_0 = "NO";
    defparam add_1120_15.INJECT1_1 = "NO";
    CCU2D add_1120_13 (.A0(d7[11]), .B0(d_d7[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[12]), .B1(d_d7[12]), .C1(GND_net), .D1(GND_net), .CIN(n11404), 
          .COUT(n11405), .S0(d8_71__N_1603[11]), .S1(d8_71__N_1603[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1120_13.INIT0 = 16'h5999;
    defparam add_1120_13.INIT1 = 16'h5999;
    defparam add_1120_13.INJECT1_0 = "NO";
    defparam add_1120_13.INJECT1_1 = "NO";
    CCU2D add_1120_11 (.A0(d7[9]), .B0(d_d7[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[10]), .B1(d_d7[10]), .C1(GND_net), .D1(GND_net), .CIN(n11403), 
          .COUT(n11404), .S0(d8_71__N_1603[9]), .S1(d8_71__N_1603[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1120_11.INIT0 = 16'h5999;
    defparam add_1120_11.INIT1 = 16'h5999;
    defparam add_1120_11.INJECT1_0 = "NO";
    defparam add_1120_11.INJECT1_1 = "NO";
    CCU2D add_1120_9 (.A0(d7[7]), .B0(d_d7[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[8]), .B1(d_d7[8]), .C1(GND_net), .D1(GND_net), .CIN(n11402), 
          .COUT(n11403), .S0(d8_71__N_1603[7]), .S1(d8_71__N_1603[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1120_9.INIT0 = 16'h5999;
    defparam add_1120_9.INIT1 = 16'h5999;
    defparam add_1120_9.INJECT1_0 = "NO";
    defparam add_1120_9.INJECT1_1 = "NO";
    CCU2D add_1120_7 (.A0(d7[5]), .B0(d_d7[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[6]), .B1(d_d7[6]), .C1(GND_net), .D1(GND_net), .CIN(n11401), 
          .COUT(n11402), .S0(d8_71__N_1603[5]), .S1(d8_71__N_1603[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1120_7.INIT0 = 16'h5999;
    defparam add_1120_7.INIT1 = 16'h5999;
    defparam add_1120_7.INJECT1_0 = "NO";
    defparam add_1120_7.INJECT1_1 = "NO";
    CCU2D add_1120_5 (.A0(d7[3]), .B0(d_d7[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[4]), .B1(d_d7[4]), .C1(GND_net), .D1(GND_net), .CIN(n11400), 
          .COUT(n11401), .S0(d8_71__N_1603[3]), .S1(d8_71__N_1603[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1120_5.INIT0 = 16'h5999;
    defparam add_1120_5.INIT1 = 16'h5999;
    defparam add_1120_5.INJECT1_0 = "NO";
    defparam add_1120_5.INJECT1_1 = "NO";
    CCU2D add_1120_3 (.A0(d7[1]), .B0(d_d7[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[2]), .B1(d_d7[2]), .C1(GND_net), .D1(GND_net), .CIN(n11399), 
          .COUT(n11400), .S0(d8_71__N_1603[1]), .S1(d8_71__N_1603[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1120_3.INIT0 = 16'h5999;
    defparam add_1120_3.INIT1 = 16'h5999;
    defparam add_1120_3.INJECT1_0 = "NO";
    defparam add_1120_3.INJECT1_1 = "NO";
    CCU2D add_1120_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d7[0]), .B1(d_d7[0]), .C1(GND_net), .D1(GND_net), .COUT(n11399), 
          .S1(d8_71__N_1603[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1120_1.INIT0 = 16'h0000;
    defparam add_1120_1.INIT1 = 16'h5999;
    defparam add_1120_1.INJECT1_0 = "NO";
    defparam add_1120_1.INJECT1_1 = "NO";
    CCU2D add_1115_37 (.A0(d6[35]), .B0(d_d6[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11398), 
          .S0(d7_71__N_1531[35]), .S1(n6275));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1115_37.INIT0 = 16'h5999;
    defparam add_1115_37.INIT1 = 16'h0000;
    defparam add_1115_37.INJECT1_0 = "NO";
    defparam add_1115_37.INJECT1_1 = "NO";
    CCU2D add_1115_35 (.A0(d6[33]), .B0(d_d6[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[34]), .B1(d_d6[34]), .C1(GND_net), .D1(GND_net), .CIN(n11397), 
          .COUT(n11398), .S0(d7_71__N_1531[33]), .S1(d7_71__N_1531[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1115_35.INIT0 = 16'h5999;
    defparam add_1115_35.INIT1 = 16'h5999;
    defparam add_1115_35.INJECT1_0 = "NO";
    defparam add_1115_35.INJECT1_1 = "NO";
    CCU2D add_1115_33 (.A0(d6[31]), .B0(d_d6[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[32]), .B1(d_d6[32]), .C1(GND_net), .D1(GND_net), .CIN(n11396), 
          .COUT(n11397), .S0(d7_71__N_1531[31]), .S1(d7_71__N_1531[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1115_33.INIT0 = 16'h5999;
    defparam add_1115_33.INIT1 = 16'h5999;
    defparam add_1115_33.INJECT1_0 = "NO";
    defparam add_1115_33.INJECT1_1 = "NO";
    CCU2D add_1115_31 (.A0(d6[29]), .B0(d_d6[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[30]), .B1(d_d6[30]), .C1(GND_net), .D1(GND_net), .CIN(n11395), 
          .COUT(n11396), .S0(d7_71__N_1531[29]), .S1(d7_71__N_1531[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1115_31.INIT0 = 16'h5999;
    defparam add_1115_31.INIT1 = 16'h5999;
    defparam add_1115_31.INJECT1_0 = "NO";
    defparam add_1115_31.INJECT1_1 = "NO";
    CCU2D add_1115_29 (.A0(d6[27]), .B0(d_d6[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[28]), .B1(d_d6[28]), .C1(GND_net), .D1(GND_net), .CIN(n11394), 
          .COUT(n11395), .S0(d7_71__N_1531[27]), .S1(d7_71__N_1531[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1115_29.INIT0 = 16'h5999;
    defparam add_1115_29.INIT1 = 16'h5999;
    defparam add_1115_29.INJECT1_0 = "NO";
    defparam add_1115_29.INJECT1_1 = "NO";
    CCU2D add_1115_27 (.A0(d6[25]), .B0(d_d6[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[26]), .B1(d_d6[26]), .C1(GND_net), .D1(GND_net), .CIN(n11393), 
          .COUT(n11394), .S0(d7_71__N_1531[25]), .S1(d7_71__N_1531[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1115_27.INIT0 = 16'h5999;
    defparam add_1115_27.INIT1 = 16'h5999;
    defparam add_1115_27.INJECT1_0 = "NO";
    defparam add_1115_27.INJECT1_1 = "NO";
    CCU2D add_1115_25 (.A0(d6[23]), .B0(d_d6[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[24]), .B1(d_d6[24]), .C1(GND_net), .D1(GND_net), .CIN(n11392), 
          .COUT(n11393), .S0(d7_71__N_1531[23]), .S1(d7_71__N_1531[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1115_25.INIT0 = 16'h5999;
    defparam add_1115_25.INIT1 = 16'h5999;
    defparam add_1115_25.INJECT1_0 = "NO";
    defparam add_1115_25.INJECT1_1 = "NO";
    CCU2D add_1115_23 (.A0(d6[21]), .B0(d_d6[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[22]), .B1(d_d6[22]), .C1(GND_net), .D1(GND_net), .CIN(n11391), 
          .COUT(n11392), .S0(d7_71__N_1531[21]), .S1(d7_71__N_1531[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1115_23.INIT0 = 16'h5999;
    defparam add_1115_23.INIT1 = 16'h5999;
    defparam add_1115_23.INJECT1_0 = "NO";
    defparam add_1115_23.INJECT1_1 = "NO";
    CCU2D add_1115_21 (.A0(d6[19]), .B0(d_d6[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[20]), .B1(d_d6[20]), .C1(GND_net), .D1(GND_net), .CIN(n11390), 
          .COUT(n11391), .S0(d7_71__N_1531[19]), .S1(d7_71__N_1531[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1115_21.INIT0 = 16'h5999;
    defparam add_1115_21.INIT1 = 16'h5999;
    defparam add_1115_21.INJECT1_0 = "NO";
    defparam add_1115_21.INJECT1_1 = "NO";
    CCU2D add_1115_19 (.A0(d6[17]), .B0(d_d6[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[18]), .B1(d_d6[18]), .C1(GND_net), .D1(GND_net), .CIN(n11389), 
          .COUT(n11390), .S0(d7_71__N_1531[17]), .S1(d7_71__N_1531[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1115_19.INIT0 = 16'h5999;
    defparam add_1115_19.INIT1 = 16'h5999;
    defparam add_1115_19.INJECT1_0 = "NO";
    defparam add_1115_19.INJECT1_1 = "NO";
    CCU2D add_1115_17 (.A0(d6[15]), .B0(d_d6[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[16]), .B1(d_d6[16]), .C1(GND_net), .D1(GND_net), .CIN(n11388), 
          .COUT(n11389), .S0(d7_71__N_1531[15]), .S1(d7_71__N_1531[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1115_17.INIT0 = 16'h5999;
    defparam add_1115_17.INIT1 = 16'h5999;
    defparam add_1115_17.INJECT1_0 = "NO";
    defparam add_1115_17.INJECT1_1 = "NO";
    CCU2D add_1115_15 (.A0(d6[13]), .B0(d_d6[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[14]), .B1(d_d6[14]), .C1(GND_net), .D1(GND_net), .CIN(n11387), 
          .COUT(n11388), .S0(d7_71__N_1531[13]), .S1(d7_71__N_1531[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1115_15.INIT0 = 16'h5999;
    defparam add_1115_15.INIT1 = 16'h5999;
    defparam add_1115_15.INJECT1_0 = "NO";
    defparam add_1115_15.INJECT1_1 = "NO";
    CCU2D add_1115_13 (.A0(d6[11]), .B0(d_d6[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[12]), .B1(d_d6[12]), .C1(GND_net), .D1(GND_net), .CIN(n11386), 
          .COUT(n11387), .S0(d7_71__N_1531[11]), .S1(d7_71__N_1531[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1115_13.INIT0 = 16'h5999;
    defparam add_1115_13.INIT1 = 16'h5999;
    defparam add_1115_13.INJECT1_0 = "NO";
    defparam add_1115_13.INJECT1_1 = "NO";
    CCU2D add_1115_11 (.A0(d6[9]), .B0(d_d6[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[10]), .B1(d_d6[10]), .C1(GND_net), .D1(GND_net), .CIN(n11385), 
          .COUT(n11386), .S0(d7_71__N_1531[9]), .S1(d7_71__N_1531[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1115_11.INIT0 = 16'h5999;
    defparam add_1115_11.INIT1 = 16'h5999;
    defparam add_1115_11.INJECT1_0 = "NO";
    defparam add_1115_11.INJECT1_1 = "NO";
    CCU2D add_1115_9 (.A0(d6[7]), .B0(d_d6[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[8]), .B1(d_d6[8]), .C1(GND_net), .D1(GND_net), .CIN(n11384), 
          .COUT(n11385), .S0(d7_71__N_1531[7]), .S1(d7_71__N_1531[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1115_9.INIT0 = 16'h5999;
    defparam add_1115_9.INIT1 = 16'h5999;
    defparam add_1115_9.INJECT1_0 = "NO";
    defparam add_1115_9.INJECT1_1 = "NO";
    CCU2D add_1115_7 (.A0(d6[5]), .B0(d_d6[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[6]), .B1(d_d6[6]), .C1(GND_net), .D1(GND_net), .CIN(n11383), 
          .COUT(n11384), .S0(d7_71__N_1531[5]), .S1(d7_71__N_1531[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1115_7.INIT0 = 16'h5999;
    defparam add_1115_7.INIT1 = 16'h5999;
    defparam add_1115_7.INJECT1_0 = "NO";
    defparam add_1115_7.INJECT1_1 = "NO";
    CCU2D add_1115_5 (.A0(d6[3]), .B0(d_d6[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[4]), .B1(d_d6[4]), .C1(GND_net), .D1(GND_net), .CIN(n11382), 
          .COUT(n11383), .S0(d7_71__N_1531[3]), .S1(d7_71__N_1531[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1115_5.INIT0 = 16'h5999;
    defparam add_1115_5.INIT1 = 16'h5999;
    defparam add_1115_5.INJECT1_0 = "NO";
    defparam add_1115_5.INJECT1_1 = "NO";
    CCU2D add_1115_3 (.A0(d6[1]), .B0(d_d6[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[2]), .B1(d_d6[2]), .C1(GND_net), .D1(GND_net), .CIN(n11381), 
          .COUT(n11382), .S0(d7_71__N_1531[1]), .S1(d7_71__N_1531[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1115_3.INIT0 = 16'h5999;
    defparam add_1115_3.INIT1 = 16'h5999;
    defparam add_1115_3.INJECT1_0 = "NO";
    defparam add_1115_3.INJECT1_1 = "NO";
    CCU2D add_1115_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d6[0]), .B1(d_d6[0]), .C1(GND_net), .D1(GND_net), .COUT(n11381), 
          .S1(d7_71__N_1531[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1115_1.INIT0 = 16'h0000;
    defparam add_1115_1.INIT1 = 16'h5999;
    defparam add_1115_1.INJECT1_0 = "NO";
    defparam add_1115_1.INJECT1_1 = "NO";
    CCU2D add_1110_37 (.A0(d_tmp[35]), .B0(d_d_tmp[35]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11380), .S0(d6_71__N_1459[35]), .S1(n6123));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1110_37.INIT0 = 16'h5999;
    defparam add_1110_37.INIT1 = 16'h0000;
    defparam add_1110_37.INJECT1_0 = "NO";
    defparam add_1110_37.INJECT1_1 = "NO";
    CCU2D add_1110_35 (.A0(d_tmp[33]), .B0(d_d_tmp[33]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[34]), .B1(d_d_tmp[34]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11379), .COUT(n11380), .S0(d6_71__N_1459[33]), 
          .S1(d6_71__N_1459[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1110_35.INIT0 = 16'h5999;
    defparam add_1110_35.INIT1 = 16'h5999;
    defparam add_1110_35.INJECT1_0 = "NO";
    defparam add_1110_35.INJECT1_1 = "NO";
    CCU2D add_1110_33 (.A0(d_tmp[31]), .B0(d_d_tmp[31]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[32]), .B1(d_d_tmp[32]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11378), .COUT(n11379), .S0(d6_71__N_1459[31]), 
          .S1(d6_71__N_1459[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1110_33.INIT0 = 16'h5999;
    defparam add_1110_33.INIT1 = 16'h5999;
    defparam add_1110_33.INJECT1_0 = "NO";
    defparam add_1110_33.INJECT1_1 = "NO";
    CCU2D add_1110_31 (.A0(d_tmp[29]), .B0(d_d_tmp[29]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[30]), .B1(d_d_tmp[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11377), .COUT(n11378), .S0(d6_71__N_1459[29]), 
          .S1(d6_71__N_1459[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1110_31.INIT0 = 16'h5999;
    defparam add_1110_31.INIT1 = 16'h5999;
    defparam add_1110_31.INJECT1_0 = "NO";
    defparam add_1110_31.INJECT1_1 = "NO";
    CCU2D add_1110_29 (.A0(d_tmp[27]), .B0(d_d_tmp[27]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[28]), .B1(d_d_tmp[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11376), .COUT(n11377), .S0(d6_71__N_1459[27]), 
          .S1(d6_71__N_1459[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1110_29.INIT0 = 16'h5999;
    defparam add_1110_29.INIT1 = 16'h5999;
    defparam add_1110_29.INJECT1_0 = "NO";
    defparam add_1110_29.INJECT1_1 = "NO";
    CCU2D add_1110_27 (.A0(d_tmp[25]), .B0(d_d_tmp[25]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[26]), .B1(d_d_tmp[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11375), .COUT(n11376), .S0(d6_71__N_1459[25]), 
          .S1(d6_71__N_1459[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1110_27.INIT0 = 16'h5999;
    defparam add_1110_27.INIT1 = 16'h5999;
    defparam add_1110_27.INJECT1_0 = "NO";
    defparam add_1110_27.INJECT1_1 = "NO";
    CCU2D add_1110_25 (.A0(d_tmp[23]), .B0(d_d_tmp[23]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[24]), .B1(d_d_tmp[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11374), .COUT(n11375), .S0(d6_71__N_1459[23]), 
          .S1(d6_71__N_1459[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1110_25.INIT0 = 16'h5999;
    defparam add_1110_25.INIT1 = 16'h5999;
    defparam add_1110_25.INJECT1_0 = "NO";
    defparam add_1110_25.INJECT1_1 = "NO";
    CCU2D add_1110_23 (.A0(d_tmp[21]), .B0(d_d_tmp[21]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[22]), .B1(d_d_tmp[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11373), .COUT(n11374), .S0(d6_71__N_1459[21]), 
          .S1(d6_71__N_1459[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1110_23.INIT0 = 16'h5999;
    defparam add_1110_23.INIT1 = 16'h5999;
    defparam add_1110_23.INJECT1_0 = "NO";
    defparam add_1110_23.INJECT1_1 = "NO";
    CCU2D add_1110_21 (.A0(d_tmp[19]), .B0(d_d_tmp[19]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[20]), .B1(d_d_tmp[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11372), .COUT(n11373), .S0(d6_71__N_1459[19]), 
          .S1(d6_71__N_1459[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1110_21.INIT0 = 16'h5999;
    defparam add_1110_21.INIT1 = 16'h5999;
    defparam add_1110_21.INJECT1_0 = "NO";
    defparam add_1110_21.INJECT1_1 = "NO";
    CCU2D add_1110_19 (.A0(d_tmp[17]), .B0(d_d_tmp[17]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[18]), .B1(d_d_tmp[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11371), .COUT(n11372), .S0(d6_71__N_1459[17]), 
          .S1(d6_71__N_1459[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1110_19.INIT0 = 16'h5999;
    defparam add_1110_19.INIT1 = 16'h5999;
    defparam add_1110_19.INJECT1_0 = "NO";
    defparam add_1110_19.INJECT1_1 = "NO";
    CCU2D add_1110_17 (.A0(d_tmp[15]), .B0(d_d_tmp[15]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[16]), .B1(d_d_tmp[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11370), .COUT(n11371), .S0(d6_71__N_1459[15]), 
          .S1(d6_71__N_1459[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1110_17.INIT0 = 16'h5999;
    defparam add_1110_17.INIT1 = 16'h5999;
    defparam add_1110_17.INJECT1_0 = "NO";
    defparam add_1110_17.INJECT1_1 = "NO";
    CCU2D add_1110_15 (.A0(d_tmp[13]), .B0(d_d_tmp[13]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[14]), .B1(d_d_tmp[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11369), .COUT(n11370), .S0(d6_71__N_1459[13]), 
          .S1(d6_71__N_1459[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1110_15.INIT0 = 16'h5999;
    defparam add_1110_15.INIT1 = 16'h5999;
    defparam add_1110_15.INJECT1_0 = "NO";
    defparam add_1110_15.INJECT1_1 = "NO";
    CCU2D add_1110_13 (.A0(d_tmp[11]), .B0(d_d_tmp[11]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[12]), .B1(d_d_tmp[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11368), .COUT(n11369), .S0(d6_71__N_1459[11]), 
          .S1(d6_71__N_1459[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1110_13.INIT0 = 16'h5999;
    defparam add_1110_13.INIT1 = 16'h5999;
    defparam add_1110_13.INJECT1_0 = "NO";
    defparam add_1110_13.INJECT1_1 = "NO";
    CCU2D add_1110_11 (.A0(d_tmp[9]), .B0(d_d_tmp[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[10]), .B1(d_d_tmp[10]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11367), .COUT(n11368), .S0(d6_71__N_1459[9]), .S1(d6_71__N_1459[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1110_11.INIT0 = 16'h5999;
    defparam add_1110_11.INIT1 = 16'h5999;
    defparam add_1110_11.INJECT1_0 = "NO";
    defparam add_1110_11.INJECT1_1 = "NO";
    CCU2D add_1110_9 (.A0(d_tmp[7]), .B0(d_d_tmp[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[8]), .B1(d_d_tmp[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11366), .COUT(n11367), .S0(d6_71__N_1459[7]), .S1(d6_71__N_1459[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1110_9.INIT0 = 16'h5999;
    defparam add_1110_9.INIT1 = 16'h5999;
    defparam add_1110_9.INJECT1_0 = "NO";
    defparam add_1110_9.INJECT1_1 = "NO";
    CCU2D add_1110_7 (.A0(d_tmp[5]), .B0(d_d_tmp[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[6]), .B1(d_d_tmp[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11365), .COUT(n11366), .S0(d6_71__N_1459[5]), .S1(d6_71__N_1459[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1110_7.INIT0 = 16'h5999;
    defparam add_1110_7.INIT1 = 16'h5999;
    defparam add_1110_7.INJECT1_0 = "NO";
    defparam add_1110_7.INJECT1_1 = "NO";
    CCU2D add_1110_5 (.A0(d_tmp[3]), .B0(d_d_tmp[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[4]), .B1(d_d_tmp[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11364), .COUT(n11365), .S0(d6_71__N_1459[3]), .S1(d6_71__N_1459[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1110_5.INIT0 = 16'h5999;
    defparam add_1110_5.INIT1 = 16'h5999;
    defparam add_1110_5.INJECT1_0 = "NO";
    defparam add_1110_5.INJECT1_1 = "NO";
    CCU2D add_1110_3 (.A0(d_tmp[1]), .B0(d_d_tmp[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[2]), .B1(d_d_tmp[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11363), .COUT(n11364), .S0(d6_71__N_1459[1]), .S1(d6_71__N_1459[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1110_3.INIT0 = 16'h5999;
    defparam add_1110_3.INIT1 = 16'h5999;
    defparam add_1110_3.INJECT1_0 = "NO";
    defparam add_1110_3.INJECT1_1 = "NO";
    CCU2D add_1110_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[0]), .B1(d_d_tmp[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n11363), .S1(d6_71__N_1459[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1110_1.INIT0 = 16'h0000;
    defparam add_1110_1.INIT1 = 16'h5999;
    defparam add_1110_1.INJECT1_0 = "NO";
    defparam add_1110_1.INJECT1_1 = "NO";
    LUT4 i5330_4_lut (.A(n12778), .B(n12503), .C(n12780), .D(count[3]), 
         .Z(count_15__N_1458)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i5330_4_lut.init = 16'h2000;
    LUT4 mux_1243_i2_3_lut (.A(n6732[21]), .B(n6770[21]), .C(n6731), .Z(d10_71__N_1747[57])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1243_i2_3_lut.init = 16'hcaca;
    LUT4 i5294_2_lut (.A(count[1]), .B(count[8]), .Z(n12778)) /* synthesis lut_function=(A (B)) */ ;
    defparam i5294_2_lut.init = 16'h8888;
    LUT4 mux_1243_i3_3_lut (.A(n6732[22]), .B(n6770[22]), .C(n6731), .Z(d10_71__N_1747[58])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1243_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1243_i4_3_lut (.A(n6732[23]), .B(n6770[23]), .C(n6731), .Z(d10_71__N_1747[59])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1243_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1243_i5_3_lut (.A(n6732[24]), .B(n6770[24]), .C(n6731), .Z(d10_71__N_1747[60])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1243_i5_3_lut.init = 16'hcaca;
    LUT4 i5296_4_lut (.A(count[0]), .B(count[2]), .C(n12), .D(n8), .Z(n12780)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5296_4_lut.init = 16'h8000;
    LUT4 mux_1243_i6_3_lut (.A(n6732[25]), .B(n6770[25]), .C(n6731), .Z(d10_71__N_1747[61])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1243_i6_3_lut.init = 16'hcaca;
    LUT4 i5_4_lut (.A(count[9]), .B(count[4]), .C(count[7]), .D(count[6]), 
         .Z(n12)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut.init = 16'h8000;
    LUT4 mux_1243_i7_3_lut (.A(n6732[26]), .B(n6770[26]), .C(n6731), .Z(d10_71__N_1747[62])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1243_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1243_i8_3_lut (.A(n6732[27]), .B(n6770[27]), .C(n6731), .Z(d10_71__N_1747[63])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1243_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1243_i9_3_lut (.A(n6732[28]), .B(n6770[28]), .C(n6731), .Z(d10_71__N_1747[64])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1243_i9_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut (.A(count[10]), .B(count[5]), .Z(n8)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i4604_2_lut (.A(d3[0]), .B(d4[0]), .Z(d4_71__N_634[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4604_2_lut.init = 16'h6666;
    LUT4 mux_1243_i10_3_lut (.A(n6732[29]), .B(n6770[29]), .C(n6731), 
         .Z(d10_71__N_1747[65])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1243_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1243_i11_3_lut (.A(n6732[30]), .B(n6770[30]), .C(n6731), 
         .Z(d10_71__N_1747[66])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1243_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1243_i12_3_lut (.A(n6732[31]), .B(n6770[31]), .C(n6731), 
         .Z(d10_71__N_1747[67])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1243_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1243_i13_3_lut (.A(n6732[32]), .B(n6770[32]), .C(n6731), 
         .Z(d10_71__N_1747[68])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1243_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1243_i14_3_lut (.A(n6732[33]), .B(n6770[33]), .C(n6731), 
         .Z(d10_71__N_1747[69])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1243_i14_3_lut.init = 16'hcaca;
    LUT4 i5361_2_lut (.A(n31), .B(n13196), .Z(n8436)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam i5361_2_lut.init = 16'hdddd;
    LUT4 i2608_2_lut (.A(n375[11]), .B(n31), .Z(count_15__N_1442[11])) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(86[13] 89[16])
    defparam i2608_2_lut.init = 16'hbbbb;
    FD1S3AX v_comb_66_rep_130 (.D(osc_clk_enable_757), .CK(osc_clk), .Q(osc_clk_enable_1397)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_130.GSR = "ENABLED";
    LUT4 i4634_2_lut (.A(d3[36]), .B(d4[36]), .Z(n5516[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4634_2_lut.init = 16'h6666;
    LUT4 i4602_2_lut (.A(d1[0]), .B(d2[0]), .Z(d2_71__N_490[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4602_2_lut.init = 16'h6666;
    LUT4 i4603_2_lut (.A(d2[0]), .B(d3[0]), .Z(d3_71__N_562[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4603_2_lut.init = 16'h6666;
    FD1S3AX v_comb_66_rep_129 (.D(osc_clk_enable_757), .CK(osc_clk), .Q(osc_clk_enable_1347)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_129.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_128 (.D(osc_clk_enable_757), .CK(osc_clk), .Q(osc_clk_enable_1297)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_128.GSR = "ENABLED";
    CCU2D add_1077_7 (.A0(d1[40]), .B0(n5059), .C0(n5060[4]), .D0(MixerOutCos[11]), 
          .A1(d1[41]), .B1(n5059), .C1(n5060[5]), .D1(MixerOutCos[11]), 
          .CIN(n11757), .COUT(n11758), .S0(d1_71__N_418[40]), .S1(d1_71__N_418[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1077_7.INIT0 = 16'h74b8;
    defparam add_1077_7.INIT1 = 16'h74b8;
    defparam add_1077_7.INJECT1_0 = "NO";
    defparam add_1077_7.INJECT1_1 = "NO";
    CCU2D add_1097_21 (.A0(d5[54]), .B0(n5667), .C0(n5668[18]), .D0(d4[54]), 
          .A1(d5[55]), .B1(n5667), .C1(n5668[19]), .D1(d4[55]), .CIN(n11600), 
          .COUT(n11601), .S0(d5_71__N_706[54]), .S1(d5_71__N_706[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1097_21.INIT0 = 16'h74b8;
    defparam add_1097_21.INIT1 = 16'h74b8;
    defparam add_1097_21.INJECT1_0 = "NO";
    defparam add_1097_21.INJECT1_1 = "NO";
    LUT4 i4640_2_lut (.A(d1[36]), .B(d2[36]), .Z(n5212[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4640_2_lut.init = 16'h6666;
    CCU2D add_1077_15 (.A0(d1[48]), .B0(n5059), .C0(n5060[12]), .D0(MixerOutCos[11]), 
          .A1(d1[49]), .B1(n5059), .C1(n5060[13]), .D1(MixerOutCos[11]), 
          .CIN(n11761), .COUT(n11762), .S0(d1_71__N_418[48]), .S1(d1_71__N_418[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1077_15.INIT0 = 16'h74b8;
    defparam add_1077_15.INIT1 = 16'h74b8;
    defparam add_1077_15.INJECT1_0 = "NO";
    defparam add_1077_15.INJECT1_1 = "NO";
    CCU2D add_1096_2 (.A0(d4[36]), .B0(d5[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[37]), .B1(d5[37]), .C1(GND_net), .D1(GND_net), .COUT(n11611), 
          .S1(n5668[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1096_2.INIT0 = 16'h7000;
    defparam add_1096_2.INIT1 = 16'h5666;
    defparam add_1096_2.INJECT1_0 = "NO";
    defparam add_1096_2.INJECT1_1 = "NO";
    FD1S3AX v_comb_66_rep_127 (.D(osc_clk_enable_757), .CK(osc_clk), .Q(osc_clk_enable_1247)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_127.GSR = "ENABLED";
    CCU2D add_1077_37 (.A0(d1[70]), .B0(n5059), .C0(n5060[34]), .D0(MixerOutCos[11]), 
          .A1(d1[71]), .B1(n5059), .C1(n5060[35]), .D1(MixerOutCos[11]), 
          .CIN(n11772), .S0(d1_71__N_418[70]), .S1(d1_71__N_418[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1077_37.INIT0 = 16'h74b8;
    defparam add_1077_37.INIT1 = 16'h74b8;
    defparam add_1077_37.INJECT1_0 = "NO";
    defparam add_1077_37.INJECT1_1 = "NO";
    CCU2D add_1077_35 (.A0(d1[68]), .B0(n5059), .C0(n5060[32]), .D0(MixerOutCos[11]), 
          .A1(d1[69]), .B1(n5059), .C1(n5060[33]), .D1(MixerOutCos[11]), 
          .CIN(n11771), .COUT(n11772), .S0(d1_71__N_418[68]), .S1(d1_71__N_418[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1077_35.INIT0 = 16'h74b8;
    defparam add_1077_35.INIT1 = 16'h74b8;
    defparam add_1077_35.INJECT1_0 = "NO";
    defparam add_1077_35.INJECT1_1 = "NO";
    CCU2D add_1077_33 (.A0(d1[66]), .B0(n5059), .C0(n5060[30]), .D0(MixerOutCos[11]), 
          .A1(d1[67]), .B1(n5059), .C1(n5060[31]), .D1(MixerOutCos[11]), 
          .CIN(n11770), .COUT(n11771), .S0(d1_71__N_418[66]), .S1(d1_71__N_418[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1077_33.INIT0 = 16'h74b8;
    defparam add_1077_33.INIT1 = 16'h74b8;
    defparam add_1077_33.INJECT1_0 = "NO";
    defparam add_1077_33.INJECT1_1 = "NO";
    FD1S3AX v_comb_66_rep_126 (.D(osc_clk_enable_757), .CK(osc_clk), .Q(osc_clk_enable_1197)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_126.GSR = "ENABLED";
    CCU2D add_1077_31 (.A0(d1[64]), .B0(n5059), .C0(n5060[28]), .D0(MixerOutCos[11]), 
          .A1(d1[65]), .B1(n5059), .C1(n5060[29]), .D1(MixerOutCos[11]), 
          .CIN(n11769), .COUT(n11770), .S0(d1_71__N_418[64]), .S1(d1_71__N_418[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1077_31.INIT0 = 16'h74b8;
    defparam add_1077_31.INIT1 = 16'h74b8;
    defparam add_1077_31.INJECT1_0 = "NO";
    defparam add_1077_31.INJECT1_1 = "NO";
    CCU2D add_1077_29 (.A0(d1[62]), .B0(n5059), .C0(n5060[26]), .D0(MixerOutCos[11]), 
          .A1(d1[63]), .B1(n5059), .C1(n5060[27]), .D1(MixerOutCos[11]), 
          .CIN(n11768), .COUT(n11769), .S0(d1_71__N_418[62]), .S1(d1_71__N_418[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1077_29.INIT0 = 16'h74b8;
    defparam add_1077_29.INIT1 = 16'h74b8;
    defparam add_1077_29.INJECT1_0 = "NO";
    defparam add_1077_29.INJECT1_1 = "NO";
    CCU2D add_1077_27 (.A0(d1[60]), .B0(n5059), .C0(n5060[24]), .D0(MixerOutCos[11]), 
          .A1(d1[61]), .B1(n5059), .C1(n5060[25]), .D1(MixerOutCos[11]), 
          .CIN(n11767), .COUT(n11768), .S0(d1_71__N_418[60]), .S1(d1_71__N_418[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1077_27.INIT0 = 16'h74b8;
    defparam add_1077_27.INIT1 = 16'h74b8;
    defparam add_1077_27.INJECT1_0 = "NO";
    defparam add_1077_27.INJECT1_1 = "NO";
    CCU2D add_1077_25 (.A0(d1[58]), .B0(n5059), .C0(n5060[22]), .D0(MixerOutCos[11]), 
          .A1(d1[59]), .B1(n5059), .C1(n5060[23]), .D1(MixerOutCos[11]), 
          .CIN(n11766), .COUT(n11767), .S0(d1_71__N_418[58]), .S1(d1_71__N_418[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1077_25.INIT0 = 16'h74b8;
    defparam add_1077_25.INIT1 = 16'h74b8;
    defparam add_1077_25.INJECT1_0 = "NO";
    defparam add_1077_25.INJECT1_1 = "NO";
    FD1S3AX v_comb_66_rep_125 (.D(osc_clk_enable_757), .CK(osc_clk), .Q(osc_clk_enable_1147)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_125.GSR = "ENABLED";
    PFUMX i5444 (.BLUT(n13089), .ALUT(n13090), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[0]));
    FD1S3AX v_comb_66_rep_124 (.D(osc_clk_enable_757), .CK(osc_clk), .Q(osc_clk_enable_1097)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_124.GSR = "ENABLED";
    LUT4 i5409_then_3_lut (.A(\CICGain[1] ), .B(\d10[60] ), .C(d10[58]), 
         .Z(n13087)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i5409_then_3_lut.init = 16'he4e4;
    LUT4 i5409_else_3_lut (.A(n62), .B(\CICGain[1] ), .C(\d10[59] ), .Z(n13086)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i5409_else_3_lut.init = 16'he2e2;
    FD1S3IX count__i1 (.D(n375[1]), .CK(osc_clk), .CD(n8436), .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i1.GSR = "ENABLED";
    LUT4 i5406_then_3_lut (.A(\CICGain[1] ), .B(\d10[59] ), .C(d10[57]), 
         .Z(n13090)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i5406_then_3_lut.init = 16'he4e4;
    PFUMX i5442 (.BLUT(n13086), .ALUT(n13087), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[1]));
    LUT4 i5406_else_3_lut (.A(n61), .B(\CICGain[1] ), .C(d10[58]), .Z(n13089)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i5406_else_3_lut.init = 16'he2e2;
    FD1S3AX v_comb_66_rep_123 (.D(osc_clk_enable_757), .CK(osc_clk), .Q(osc_clk_enable_1047)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_123.GSR = "ENABLED";
    LUT4 i5330_4_lut_rep_116 (.A(n12778), .B(n12503), .C(n12780), .D(count[3]), 
         .Z(osc_clk_enable_757)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i5330_4_lut_rep_116.init = 16'h2000;
    FD1S3AX v_comb_66_rep_122 (.D(osc_clk_enable_757), .CK(osc_clk), .Q(osc_clk_enable_997)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_122.GSR = "ENABLED";
    CCU2D add_1077_23 (.A0(d1[56]), .B0(n5059), .C0(n5060[20]), .D0(MixerOutCos[11]), 
          .A1(d1[57]), .B1(n5059), .C1(n5060[21]), .D1(MixerOutCos[11]), 
          .CIN(n11765), .COUT(n11766), .S0(d1_71__N_418[56]), .S1(d1_71__N_418[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1077_23.INIT0 = 16'h74b8;
    defparam add_1077_23.INIT1 = 16'h74b8;
    defparam add_1077_23.INJECT1_0 = "NO";
    defparam add_1077_23.INJECT1_1 = "NO";
    CCU2D add_1077_21 (.A0(d1[54]), .B0(n5059), .C0(n5060[18]), .D0(MixerOutCos[11]), 
          .A1(d1[55]), .B1(n5059), .C1(n5060[19]), .D1(MixerOutCos[11]), 
          .CIN(n11764), .COUT(n11765), .S0(d1_71__N_418[54]), .S1(d1_71__N_418[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1077_21.INIT0 = 16'h74b8;
    defparam add_1077_21.INIT1 = 16'h74b8;
    defparam add_1077_21.INJECT1_0 = "NO";
    defparam add_1077_21.INJECT1_1 = "NO";
    FD1S3AX v_comb_66_rep_121 (.D(osc_clk_enable_757), .CK(osc_clk), .Q(osc_clk_enable_947)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_121.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_120 (.D(osc_clk_enable_757), .CK(osc_clk), .Q(osc_clk_enable_897)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_120.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_119 (.D(osc_clk_enable_757), .CK(osc_clk), .Q(osc_clk_enable_847)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_119.GSR = "ENABLED";
    CCU2D add_1077_13 (.A0(d1[46]), .B0(n5059), .C0(n5060[10]), .D0(MixerOutCos[11]), 
          .A1(d1[47]), .B1(n5059), .C1(n5060[11]), .D1(MixerOutCos[11]), 
          .CIN(n11760), .COUT(n11761), .S0(d1_71__N_418[46]), .S1(d1_71__N_418[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1077_13.INIT0 = 16'h74b8;
    defparam add_1077_13.INIT1 = 16'h74b8;
    defparam add_1077_13.INJECT1_0 = "NO";
    defparam add_1077_13.INJECT1_1 = "NO";
    FD1S3AX v_comb_66_rep_118 (.D(osc_clk_enable_757), .CK(osc_clk), .Q(osc_clk_enable_797)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=180, LSE_RLINE=186 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_118.GSR = "ENABLED";
    CCU2D add_1077_11 (.A0(d1[44]), .B0(n5059), .C0(n5060[8]), .D0(MixerOutCos[11]), 
          .A1(d1[45]), .B1(n5059), .C1(n5060[9]), .D1(MixerOutCos[11]), 
          .CIN(n11759), .COUT(n11760), .S0(d1_71__N_418[44]), .S1(d1_71__N_418[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1077_11.INIT0 = 16'h74b8;
    defparam add_1077_11.INIT1 = 16'h74b8;
    defparam add_1077_11.INJECT1_0 = "NO";
    defparam add_1077_11.INJECT1_1 = "NO";
    CCU2D add_1077_9 (.A0(d1[42]), .B0(n5059), .C0(n5060[6]), .D0(MixerOutCos[11]), 
          .A1(d1[43]), .B1(n5059), .C1(n5060[7]), .D1(MixerOutCos[11]), 
          .CIN(n11758), .COUT(n11759), .S0(d1_71__N_418[42]), .S1(d1_71__N_418[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1077_9.INIT0 = 16'h74b8;
    defparam add_1077_9.INIT1 = 16'h74b8;
    defparam add_1077_9.INJECT1_0 = "NO";
    defparam add_1077_9.INJECT1_1 = "NO";
    CCU2D add_1077_19 (.A0(d1[52]), .B0(n5059), .C0(n5060[16]), .D0(MixerOutCos[11]), 
          .A1(d1[53]), .B1(n5059), .C1(n5060[17]), .D1(MixerOutCos[11]), 
          .CIN(n11763), .COUT(n11764), .S0(d1_71__N_418[52]), .S1(d1_71__N_418[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1077_19.INIT0 = 16'h74b8;
    defparam add_1077_19.INIT1 = 16'h74b8;
    defparam add_1077_19.INJECT1_0 = "NO";
    defparam add_1077_19.INJECT1_1 = "NO";
    CCU2D add_1077_17 (.A0(d1[50]), .B0(n5059), .C0(n5060[14]), .D0(MixerOutCos[11]), 
          .A1(d1[51]), .B1(n5059), .C1(n5060[15]), .D1(MixerOutCos[11]), 
          .CIN(n11762), .COUT(n11763), .S0(d1_71__N_418[50]), .S1(d1_71__N_418[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1077_17.INIT0 = 16'h74b8;
    defparam add_1077_17.INIT1 = 16'h74b8;
    defparam add_1077_17.INJECT1_0 = "NO";
    defparam add_1077_17.INJECT1_1 = "NO";
    CCU2D add_1082_11 (.A0(d2[44]), .B0(n5211), .C0(n5212[8]), .D0(d1[44]), 
          .A1(d2[45]), .B1(n5211), .C1(n5212[9]), .D1(d1[45]), .CIN(n11718), 
          .COUT(n11719), .S0(d2_71__N_490[44]), .S1(d2_71__N_490[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1082_11.INIT0 = 16'h74b8;
    defparam add_1082_11.INIT1 = 16'h74b8;
    defparam add_1082_11.INJECT1_0 = "NO";
    defparam add_1082_11.INJECT1_1 = "NO";
    CCU2D add_1076_36 (.A0(MixerOutCos[11]), .B0(d1[70]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[71]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11791), .S0(n5060[34]), .S1(n5060[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1076_36.INIT0 = 16'h5666;
    defparam add_1076_36.INIT1 = 16'h5666;
    defparam add_1076_36.INJECT1_0 = "NO";
    defparam add_1076_36.INJECT1_1 = "NO";
    CCU2D add_1076_34 (.A0(MixerOutCos[11]), .B0(d1[68]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[69]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11790), .COUT(n11791), .S0(n5060[32]), 
          .S1(n5060[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1076_34.INIT0 = 16'h5666;
    defparam add_1076_34.INIT1 = 16'h5666;
    defparam add_1076_34.INJECT1_0 = "NO";
    defparam add_1076_34.INJECT1_1 = "NO";
    CCU2D add_1076_32 (.A0(MixerOutCos[11]), .B0(d1[66]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[67]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11789), .COUT(n11790), .S0(n5060[30]), 
          .S1(n5060[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1076_32.INIT0 = 16'h5666;
    defparam add_1076_32.INIT1 = 16'h5666;
    defparam add_1076_32.INJECT1_0 = "NO";
    defparam add_1076_32.INJECT1_1 = "NO";
    CCU2D add_1076_30 (.A0(MixerOutCos[11]), .B0(d1[64]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[65]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11788), .COUT(n11789), .S0(n5060[28]), 
          .S1(n5060[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1076_30.INIT0 = 16'h5666;
    defparam add_1076_30.INIT1 = 16'h5666;
    defparam add_1076_30.INJECT1_0 = "NO";
    defparam add_1076_30.INJECT1_1 = "NO";
    CCU2D add_1076_28 (.A0(MixerOutCos[11]), .B0(d1[62]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[63]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11787), .COUT(n11788), .S0(n5060[26]), 
          .S1(n5060[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1076_28.INIT0 = 16'h5666;
    defparam add_1076_28.INIT1 = 16'h5666;
    defparam add_1076_28.INJECT1_0 = "NO";
    defparam add_1076_28.INJECT1_1 = "NO";
    CCU2D add_1076_26 (.A0(MixerOutCos[11]), .B0(d1[60]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[61]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11786), .COUT(n11787), .S0(n5060[24]), 
          .S1(n5060[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1076_26.INIT0 = 16'h5666;
    defparam add_1076_26.INIT1 = 16'h5666;
    defparam add_1076_26.INJECT1_0 = "NO";
    defparam add_1076_26.INJECT1_1 = "NO";
    CCU2D add_1076_24 (.A0(MixerOutCos[11]), .B0(d1[58]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[59]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11785), .COUT(n11786), .S0(n5060[22]), 
          .S1(n5060[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1076_24.INIT0 = 16'h5666;
    defparam add_1076_24.INIT1 = 16'h5666;
    defparam add_1076_24.INJECT1_0 = "NO";
    defparam add_1076_24.INJECT1_1 = "NO";
    CCU2D add_1076_22 (.A0(MixerOutCos[11]), .B0(d1[56]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[57]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11784), .COUT(n11785), .S0(n5060[20]), 
          .S1(n5060[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1076_22.INIT0 = 16'h5666;
    defparam add_1076_22.INIT1 = 16'h5666;
    defparam add_1076_22.INJECT1_0 = "NO";
    defparam add_1076_22.INJECT1_1 = "NO";
    CCU2D add_1076_20 (.A0(MixerOutCos[11]), .B0(d1[54]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[55]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11783), .COUT(n11784), .S0(n5060[18]), 
          .S1(n5060[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1076_20.INIT0 = 16'h5666;
    defparam add_1076_20.INIT1 = 16'h5666;
    defparam add_1076_20.INJECT1_0 = "NO";
    defparam add_1076_20.INJECT1_1 = "NO";
    CCU2D add_1076_18 (.A0(MixerOutCos[11]), .B0(d1[52]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[53]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11782), .COUT(n11783), .S0(n5060[16]), 
          .S1(n5060[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1076_18.INIT0 = 16'h5666;
    defparam add_1076_18.INIT1 = 16'h5666;
    defparam add_1076_18.INJECT1_0 = "NO";
    defparam add_1076_18.INJECT1_1 = "NO";
    CCU2D add_1076_16 (.A0(MixerOutCos[11]), .B0(d1[50]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[51]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11781), .COUT(n11782), .S0(n5060[14]), 
          .S1(n5060[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1076_16.INIT0 = 16'h5666;
    defparam add_1076_16.INIT1 = 16'h5666;
    defparam add_1076_16.INJECT1_0 = "NO";
    defparam add_1076_16.INJECT1_1 = "NO";
    CCU2D add_1076_14 (.A0(MixerOutCos[11]), .B0(d1[48]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[49]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11780), .COUT(n11781), .S0(n5060[12]), 
          .S1(n5060[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1076_14.INIT0 = 16'h5666;
    defparam add_1076_14.INIT1 = 16'h5666;
    defparam add_1076_14.INJECT1_0 = "NO";
    defparam add_1076_14.INJECT1_1 = "NO";
    CCU2D add_1076_12 (.A0(MixerOutCos[11]), .B0(d1[46]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[47]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11779), .COUT(n11780), .S0(n5060[10]), 
          .S1(n5060[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1076_12.INIT0 = 16'h5666;
    defparam add_1076_12.INIT1 = 16'h5666;
    defparam add_1076_12.INJECT1_0 = "NO";
    defparam add_1076_12.INJECT1_1 = "NO";
    CCU2D add_1076_10 (.A0(MixerOutCos[11]), .B0(d1[44]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[45]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11778), .COUT(n11779), .S0(n5060[8]), 
          .S1(n5060[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1076_10.INIT0 = 16'h5666;
    defparam add_1076_10.INIT1 = 16'h5666;
    defparam add_1076_10.INJECT1_0 = "NO";
    defparam add_1076_10.INJECT1_1 = "NO";
    CCU2D add_1076_8 (.A0(MixerOutCos[11]), .B0(d1[42]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[43]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11777), .COUT(n11778), .S0(n5060[6]), 
          .S1(n5060[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1076_8.INIT0 = 16'h5666;
    defparam add_1076_8.INIT1 = 16'h5666;
    defparam add_1076_8.INJECT1_0 = "NO";
    defparam add_1076_8.INJECT1_1 = "NO";
    CCU2D add_1076_6 (.A0(MixerOutCos[11]), .B0(d1[40]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[41]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11776), .COUT(n11777), .S0(n5060[4]), 
          .S1(n5060[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1076_6.INIT0 = 16'h5666;
    defparam add_1076_6.INIT1 = 16'h5666;
    defparam add_1076_6.INJECT1_0 = "NO";
    defparam add_1076_6.INJECT1_1 = "NO";
    CCU2D add_1076_4 (.A0(MixerOutCos[11]), .B0(d1[38]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[39]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11775), .COUT(n11776), .S0(n5060[2]), 
          .S1(n5060[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1076_4.INIT0 = 16'h5666;
    defparam add_1076_4.INIT1 = 16'h5666;
    defparam add_1076_4.INJECT1_0 = "NO";
    defparam add_1076_4.INJECT1_1 = "NO";
    CCU2D add_1076_2 (.A0(MixerOutCos[11]), .B0(d1[36]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[37]), .C1(GND_net), 
          .D1(GND_net), .COUT(n11775), .S1(n5060[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1076_2.INIT0 = 16'h7000;
    defparam add_1076_2.INIT1 = 16'h5666;
    defparam add_1076_2.INJECT1_0 = "NO";
    defparam add_1076_2.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module AMDemodulator
//

module AMDemodulator (CIC1_out_clkSin, \CIC1_outSin[0] , CIC1_outCos, 
            \DataInReg_11__N_1856[0] , GND_net, \CIC1_outSin[1] , \CIC1_outSin[2] , 
            \CIC1_outSin[3] , \CIC1_outSin[4] , \CIC1_outSin[5] , MYLED_c_0, 
            MYLED_c_1, MYLED_c_2, MYLED_c_3, MYLED_c_4, MYLED_c_5, 
            \DataInReg_11__N_1856[1] , \DataInReg_11__N_1856[2] , \DataInReg_11__N_1856[3] , 
            \DataInReg_11__N_1856[4] , \DataInReg_11__N_1856[5] , \DataInReg_11__N_1856[6] , 
            \DataInReg_11__N_1856[7] , \DataInReg_11__N_1856[8] , \DemodOut[9] , 
            VCC_net) /* synthesis syn_module_defined=1 */ ;
    input CIC1_out_clkSin;
    input \CIC1_outSin[0] ;
    input [11:0]CIC1_outCos;
    output \DataInReg_11__N_1856[0] ;
    input GND_net;
    input \CIC1_outSin[1] ;
    input \CIC1_outSin[2] ;
    input \CIC1_outSin[3] ;
    input \CIC1_outSin[4] ;
    input \CIC1_outSin[5] ;
    input MYLED_c_0;
    input MYLED_c_1;
    input MYLED_c_2;
    input MYLED_c_3;
    input MYLED_c_4;
    input MYLED_c_5;
    output \DataInReg_11__N_1856[1] ;
    output \DataInReg_11__N_1856[2] ;
    output \DataInReg_11__N_1856[3] ;
    output \DataInReg_11__N_1856[4] ;
    output \DataInReg_11__N_1856[5] ;
    output \DataInReg_11__N_1856[6] ;
    output \DataInReg_11__N_1856[7] ;
    output \DataInReg_11__N_1856[8] ;
    output \DemodOut[9] ;
    input VCC_net;
    
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(85[6:21])
    wire [11:0]MultDataB;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(29[21:30])
    wire [11:0]MultDataC;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(33[21:30])
    wire [31:0]ISquare;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(24[14:21])
    wire [31:0]ISquare_31__N_1895;
    wire [15:0]d_out_d;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(20[21:28])
    wire [17:0]d_out_d_11__N_1894;
    wire [17:0]d_out_d_11__N_2335;
    wire [17:0]d_out_d_11__N_2353;
    wire [17:0]d_out_d_11__N_1892;
    wire [17:0]d_out_d_11__N_1872;
    
    wire d_out_d_11__N_1871, n12154;
    wire [17:0]d_out_d_11__N_1890;
    
    wire d_out_d_11__N_1889;
    wire [17:0]d_out_d_11__N_1888;
    
    wire d_out_d_11__N_1887;
    wire [17:0]d_out_d_11__N_1886;
    
    wire d_out_d_11__N_1885;
    wire [17:0]d_out_d_11__N_1884;
    
    wire d_out_d_11__N_1883;
    wire [17:0]d_out_d_11__N_1882;
    
    wire d_out_d_11__N_1881, n11503;
    wire [17:0]d_out_d_11__N_1874;
    
    wire d_out_d_11__N_1873;
    wire [17:0]d_out_d_11__N_1876;
    
    wire n11502, n11501, n11500, n11499, n11498;
    wire [17:0]d_out_d_11__N_1880;
    
    wire d_out_d_11__N_1879;
    wire [17:0]d_out_d_11__N_1878;
    
    wire d_out_d_11__N_1877;
    wire [23:0]MultResult1;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(30[22:33])
    wire [23:0]MultResult2;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(35[22:33])
    
    wire d_out_d_11__N_1875, n11492, n11491, n12158, n12157, n209, 
        n12156, n11490, n11489, n11488, n11487, d_out_d_11__N_1891, 
        n10951, n10950, n10949, n10948, n10947, n10946, n10945, 
        n10944, n10943, n10942, n10941, n10940, n10702, n10701, 
        n10700, n10699, n10698, n12152, n12151, n12150, n12149, 
        n12148, n12147, n12146, n12145, n11486, n12139, n12138, 
        n12137, n12136, n12135, n12134, n12133, n12132, n11485, 
        n11465, n11464, n11463, n11462, n11461, n11460, n11459, 
        n11458, n11457, n11361, n11360, n11359, n11358, n11357, 
        n11356, n11355, n11354, n11353, n12104, n12103, n12102, 
        n12101, n12100, n12099, n12098, n12097, n12096, n12090, 
        n12089, n12088, n12087, n12086, n12085, n12084, n12083, 
        n12082, n12076, n12075, n12074, n12073, n12072, n12071, 
        n12070, n12069, n12068, n12062, n12061, n12060, n12059, 
        n12058, n12057, n12056, n12055, n12054, n12048, n12047, 
        n12046, n12045, n12044, n12043, n12042;
    
    FD1S3AX MultDataB_i0 (.D(\CIC1_outSin[0] ), .CK(CIC1_out_clkSin), .Q(MultDataB[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i0.GSR = "ENABLED";
    FD1S3AX MultDataC_i0 (.D(CIC1_outCos[0]), .CK(CIC1_out_clkSin), .Q(MultDataC[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i0.GSR = "ENABLED";
    FD1S3AX ISquare_i1 (.D(ISquare_31__N_1895[0]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i1.GSR = "ENABLED";
    FD1S3AX d_out_i1 (.D(d_out_d[0]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i1.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i1 (.D(d_out_d_11__N_1894[17]), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i1.GSR = "ENABLED";
    LUT4 mux_82_i1_3_lut (.A(d_out_d_11__N_2335[17]), .B(d_out_d_11__N_2353[17]), 
         .C(d_out_d_11__N_1892[17]), .Z(d_out_d_11__N_1894[17])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam mux_82_i1_3_lut.init = 16'h3535;
    LUT4 d_out_d_11__I_0_1_lut (.A(d_out_d_11__N_1872[17]), .Z(d_out_d_11__N_1871)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_0_1_lut.init = 16'h5555;
    LUT4 i4673_2_lut (.A(ISquare[23]), .B(ISquare[22]), .Z(n12154)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i4673_2_lut.init = 16'h9999;
    LUT4 d_out_d_11__I_9_1_lut (.A(d_out_d_11__N_1890[17]), .Z(d_out_d_11__N_1889)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_9_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_8_1_lut (.A(d_out_d_11__N_1888[17]), .Z(d_out_d_11__N_1887)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_8_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_7_1_lut (.A(d_out_d_11__N_1886[17]), .Z(d_out_d_11__N_1885)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_7_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_6_1_lut (.A(d_out_d_11__N_1884[17]), .Z(d_out_d_11__N_1883)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_6_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_5_1_lut (.A(d_out_d_11__N_1882[17]), .Z(d_out_d_11__N_1881)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_5_1_lut.init = 16'h5555;
    CCU2D add_457_13 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1873), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1874[17]), .B1(d_out_d_11__N_1873), 
          .C1(GND_net), .D1(GND_net), .CIN(n11503), .S0(d_out_d_11__N_1876[9]), 
          .S1(d_out_d_11__N_1876[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_457_13.INIT0 = 16'h5666;
    defparam add_457_13.INIT1 = 16'h5666;
    defparam add_457_13.INJECT1_0 = "NO";
    defparam add_457_13.INJECT1_1 = "NO";
    CCU2D add_457_11 (.A0(d_out_d_11__N_1874[6]), .B0(d_out_d_11__N_1874[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1874[7]), .B1(d_out_d_11__N_1874[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11502), .COUT(n11503), .S0(d_out_d_11__N_1876[7]), 
          .S1(d_out_d_11__N_1876[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_457_11.INIT0 = 16'h5999;
    defparam add_457_11.INIT1 = 16'h5999;
    defparam add_457_11.INJECT1_0 = "NO";
    defparam add_457_11.INJECT1_1 = "NO";
    CCU2D add_457_9 (.A0(ISquare[31]), .B0(d_out_d_11__N_1874[17]), .C0(d_out_d_11__N_1874[4]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1874[17]), 
          .C1(d_out_d_11__N_1874[5]), .D1(GND_net), .CIN(n11501), .COUT(n11502), 
          .S0(d_out_d_11__N_1876[5]), .S1(d_out_d_11__N_1876[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_457_9.INIT0 = 16'h6969;
    defparam add_457_9.INIT1 = 16'h6969;
    defparam add_457_9.INJECT1_0 = "NO";
    defparam add_457_9.INJECT1_1 = "NO";
    CCU2D add_457_7 (.A0(d_out_d_11__N_1874[2]), .B0(d_out_d_11__N_1874[17]), 
          .C0(GND_net), .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1874[17]), 
          .C1(d_out_d_11__N_1874[3]), .D1(GND_net), .CIN(n11500), .COUT(n11501), 
          .S0(d_out_d_11__N_1876[3]), .S1(d_out_d_11__N_1876[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_457_7.INIT0 = 16'h5999;
    defparam add_457_7.INIT1 = 16'h6969;
    defparam add_457_7.INJECT1_0 = "NO";
    defparam add_457_7.INJECT1_1 = "NO";
    CCU2D add_457_5 (.A0(d_out_d_11__N_1874[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1872[17]), .B1(d_out_d_11__N_1874[17]), 
          .C1(d_out_d_11__N_1874[1]), .D1(GND_net), .CIN(n11499), .COUT(n11500), 
          .S0(d_out_d_11__N_1876[1]), .S1(d_out_d_11__N_1876[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_457_5.INIT0 = 16'h5aaa;
    defparam add_457_5.INIT1 = 16'h9696;
    defparam add_457_5.INJECT1_0 = "NO";
    defparam add_457_5.INJECT1_1 = "NO";
    CCU2D add_457_3 (.A0(ISquare[18]), .B0(d_out_d_11__N_1874[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11498), .COUT(n11499), .S1(d_out_d_11__N_1876[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_457_3.INIT0 = 16'h5666;
    defparam add_457_3.INIT1 = 16'h5555;
    defparam add_457_3.INJECT1_0 = "NO";
    defparam add_457_3.INJECT1_1 = "NO";
    LUT4 d_out_d_11__I_4_1_lut (.A(d_out_d_11__N_1880[17]), .Z(d_out_d_11__N_1879)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_4_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_3_1_lut (.A(d_out_d_11__N_1878[17]), .Z(d_out_d_11__N_1877)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_3_1_lut.init = 16'h5555;
    LUT4 i4606_2_lut (.A(MultResult1[0]), .B(MultResult2[0]), .Z(ISquare_31__N_1895[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4606_2_lut.init = 16'h6666;
    LUT4 d_out_d_11__I_2_1_lut (.A(d_out_d_11__N_1876[17]), .Z(d_out_d_11__N_1875)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_2_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_1_1_lut (.A(d_out_d_11__N_1874[17]), .Z(d_out_d_11__N_1873)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_1_1_lut.init = 16'h5555;
    FD1S3AX MultDataB_i1 (.D(\CIC1_outSin[1] ), .CK(CIC1_out_clkSin), .Q(MultDataB[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i1.GSR = "ENABLED";
    FD1S3AX MultDataB_i2 (.D(\CIC1_outSin[2] ), .CK(CIC1_out_clkSin), .Q(MultDataB[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i2.GSR = "ENABLED";
    FD1S3AX MultDataB_i3 (.D(\CIC1_outSin[3] ), .CK(CIC1_out_clkSin), .Q(MultDataB[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i3.GSR = "ENABLED";
    FD1S3AX MultDataB_i4 (.D(\CIC1_outSin[4] ), .CK(CIC1_out_clkSin), .Q(MultDataB[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i4.GSR = "ENABLED";
    FD1S3AX MultDataB_i5 (.D(\CIC1_outSin[5] ), .CK(CIC1_out_clkSin), .Q(MultDataB[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i5.GSR = "ENABLED";
    FD1S3AX MultDataB_i6 (.D(MYLED_c_0), .CK(CIC1_out_clkSin), .Q(MultDataB[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i6.GSR = "ENABLED";
    FD1S3AX MultDataB_i7 (.D(MYLED_c_1), .CK(CIC1_out_clkSin), .Q(MultDataB[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i7.GSR = "ENABLED";
    FD1S3AX MultDataB_i8 (.D(MYLED_c_2), .CK(CIC1_out_clkSin), .Q(MultDataB[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i8.GSR = "ENABLED";
    FD1S3AX MultDataB_i9 (.D(MYLED_c_3), .CK(CIC1_out_clkSin), .Q(MultDataB[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i9.GSR = "ENABLED";
    FD1S3AX MultDataB_i10 (.D(MYLED_c_4), .CK(CIC1_out_clkSin), .Q(MultDataB[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i10.GSR = "ENABLED";
    FD1S3AX MultDataB_i11 (.D(MYLED_c_5), .CK(CIC1_out_clkSin), .Q(MultDataB[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i11.GSR = "ENABLED";
    FD1S3AX MultDataC_i1 (.D(CIC1_outCos[1]), .CK(CIC1_out_clkSin), .Q(MultDataC[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i1.GSR = "ENABLED";
    FD1S3AX MultDataC_i2 (.D(CIC1_outCos[2]), .CK(CIC1_out_clkSin), .Q(MultDataC[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i2.GSR = "ENABLED";
    FD1S3AX MultDataC_i3 (.D(CIC1_outCos[3]), .CK(CIC1_out_clkSin), .Q(MultDataC[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i3.GSR = "ENABLED";
    FD1S3AX MultDataC_i4 (.D(CIC1_outCos[4]), .CK(CIC1_out_clkSin), .Q(MultDataC[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i4.GSR = "ENABLED";
    FD1S3AX MultDataC_i5 (.D(CIC1_outCos[5]), .CK(CIC1_out_clkSin), .Q(MultDataC[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i5.GSR = "ENABLED";
    FD1S3AX MultDataC_i6 (.D(CIC1_outCos[6]), .CK(CIC1_out_clkSin), .Q(MultDataC[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i6.GSR = "ENABLED";
    FD1S3AX MultDataC_i7 (.D(CIC1_outCos[7]), .CK(CIC1_out_clkSin), .Q(MultDataC[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i7.GSR = "ENABLED";
    FD1S3AX MultDataC_i8 (.D(CIC1_outCos[8]), .CK(CIC1_out_clkSin), .Q(MultDataC[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i8.GSR = "ENABLED";
    FD1S3AX MultDataC_i9 (.D(CIC1_outCos[9]), .CK(CIC1_out_clkSin), .Q(MultDataC[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i9.GSR = "ENABLED";
    FD1S3AX MultDataC_i10 (.D(CIC1_outCos[10]), .CK(CIC1_out_clkSin), .Q(MultDataC[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i10.GSR = "ENABLED";
    FD1S3AX MultDataC_i11 (.D(CIC1_outCos[11]), .CK(CIC1_out_clkSin), .Q(MultDataC[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i11.GSR = "ENABLED";
    FD1S3AX ISquare_i2 (.D(ISquare_31__N_1895[1]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i2.GSR = "ENABLED";
    FD1S3AX ISquare_i3 (.D(ISquare_31__N_1895[2]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i3.GSR = "ENABLED";
    FD1S3AX ISquare_i4 (.D(ISquare_31__N_1895[3]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i4.GSR = "ENABLED";
    FD1S3AX ISquare_i5 (.D(ISquare_31__N_1895[4]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i5.GSR = "ENABLED";
    FD1S3AX ISquare_i6 (.D(ISquare_31__N_1895[5]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i6.GSR = "ENABLED";
    FD1S3AX ISquare_i7 (.D(ISquare_31__N_1895[6]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i7.GSR = "ENABLED";
    FD1S3AX ISquare_i8 (.D(ISquare_31__N_1895[7]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i8.GSR = "ENABLED";
    FD1S3AX ISquare_i9 (.D(ISquare_31__N_1895[8]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i9.GSR = "ENABLED";
    FD1S3AX ISquare_i10 (.D(ISquare_31__N_1895[9]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i10.GSR = "ENABLED";
    FD1S3AX ISquare_i11 (.D(ISquare_31__N_1895[10]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i11.GSR = "ENABLED";
    FD1S3AX ISquare_i12 (.D(ISquare_31__N_1895[11]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i12.GSR = "ENABLED";
    FD1S3AX ISquare_i13 (.D(ISquare_31__N_1895[12]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i13.GSR = "ENABLED";
    FD1S3AX ISquare_i14 (.D(ISquare_31__N_1895[13]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i14.GSR = "ENABLED";
    FD1S3AX ISquare_i15 (.D(ISquare_31__N_1895[14]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i15.GSR = "ENABLED";
    FD1S3AX ISquare_i16 (.D(ISquare_31__N_1895[15]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i16.GSR = "ENABLED";
    FD1S3AX ISquare_i17 (.D(ISquare_31__N_1895[16]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i17.GSR = "ENABLED";
    FD1S3AX ISquare_i18 (.D(ISquare_31__N_1895[17]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i18.GSR = "ENABLED";
    FD1S3AX ISquare_i19 (.D(ISquare_31__N_1895[18]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i19.GSR = "ENABLED";
    FD1S3AX ISquare_i20 (.D(ISquare_31__N_1895[19]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i20.GSR = "ENABLED";
    FD1S3AX ISquare_i21 (.D(ISquare_31__N_1895[20]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i21.GSR = "ENABLED";
    FD1S3AX ISquare_i22 (.D(ISquare_31__N_1895[21]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i22.GSR = "ENABLED";
    FD1S3AX ISquare_i23 (.D(ISquare_31__N_1895[22]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i23.GSR = "ENABLED";
    FD1S3AX ISquare_i24 (.D(ISquare_31__N_1895[23]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i24.GSR = "ENABLED";
    FD1S3AX ISquare_i25 (.D(ISquare_31__N_1895[24]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i25.GSR = "ENABLED";
    FD1S3AX d_out_i2 (.D(d_out_d[1]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i2.GSR = "ENABLED";
    FD1S3AX d_out_i3 (.D(d_out_d[2]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i3.GSR = "ENABLED";
    FD1S3AX d_out_i4 (.D(d_out_d[3]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i4.GSR = "ENABLED";
    FD1S3AX d_out_i5 (.D(d_out_d[4]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i5.GSR = "ENABLED";
    FD1S3AX d_out_i6 (.D(d_out_d[5]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i6.GSR = "ENABLED";
    FD1S3AX d_out_i7 (.D(d_out_d[6]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i7.GSR = "ENABLED";
    FD1S3AX d_out_i8 (.D(d_out_d[7]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i8.GSR = "ENABLED";
    FD1S3AX d_out_i9 (.D(d_out_d[8]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i9.GSR = "ENABLED";
    FD1S3AX d_out_i10 (.D(d_out_d[9]), .CK(CIC1_out_clkSin), .Q(\DemodOut[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=212, LSE_RLINE=217 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i10.GSR = "ENABLED";
    CCU2D add_457_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1874[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n11498));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_457_1.INIT0 = 16'hF000;
    defparam add_457_1.INIT1 = 16'h0aaa;
    defparam add_457_1.INJECT1_0 = "NO";
    defparam add_457_1.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_18 (.A0(d_out_d_11__N_1892[14]), .B0(ISquare[31]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[15]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n11492), .S1(d_out_d_11__N_2335[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_18.INIT0 = 16'h5999;
    defparam sub_78_add_2_18.INIT1 = 16'h5555;
    defparam sub_78_add_2_18.INJECT1_0 = "NO";
    defparam sub_78_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_16 (.A0(d_out_d_11__N_1892[12]), .B0(ISquare[31]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[13]), .B1(ISquare[31]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11491), .COUT(n11492));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_16.INIT0 = 16'h5999;
    defparam sub_78_add_2_16.INIT1 = 16'h5999;
    defparam sub_78_add_2_16.INJECT1_0 = "NO";
    defparam sub_78_add_2_16.INJECT1_1 = "NO";
    CCU2D add_3130_8 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n12158), 
          .S0(d_out_d_11__N_1872[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_3130_8.INIT0 = 16'h0fff;
    defparam add_3130_8.INIT1 = 16'h0000;
    defparam add_3130_8.INJECT1_0 = "NO";
    defparam add_3130_8.INJECT1_1 = "NO";
    CCU2D add_3130_6 (.A0(n209), .B0(ISquare[31]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n12157), 
          .COUT(n12158), .S0(d_out_d_11__N_1872[4]), .S1(d_out_d_11__N_1872[5]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_3130_6.INIT0 = 16'h5666;
    defparam add_3130_6.INIT1 = 16'h0fff;
    defparam add_3130_6.INJECT1_0 = "NO";
    defparam add_3130_6.INJECT1_1 = "NO";
    CCU2D add_3130_4 (.A0(n209), .B0(ISquare[31]), .C0(GND_net), .D0(GND_net), 
          .A1(ISquare[31]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12156), .COUT(n12157), .S0(d_out_d_11__N_1872[2]), .S1(d_out_d_11__N_1872[3]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_3130_4.INIT0 = 16'h5666;
    defparam add_3130_4.INIT1 = 16'h0555;
    defparam add_3130_4.INJECT1_0 = "NO";
    defparam add_3130_4.INJECT1_1 = "NO";
    CCU2D add_3130_2 (.A0(ISquare[23]), .B0(ISquare[22]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n12156), .S1(d_out_d_11__N_1872[1]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_3130_2.INIT0 = 16'h1000;
    defparam add_3130_2.INIT1 = 16'h0fff;
    defparam add_3130_2.INJECT1_0 = "NO";
    defparam add_3130_2.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_14 (.A0(d_out_d_11__N_1892[10]), .B0(d_out_d_11__N_1872[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[11]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n11490), .COUT(n11491));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_14.INIT0 = 16'h5666;
    defparam sub_78_add_2_14.INIT1 = 16'h5555;
    defparam sub_78_add_2_14.INJECT1_0 = "NO";
    defparam sub_78_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_12 (.A0(d_out_d_11__N_1892[8]), .B0(d_out_d_11__N_1876[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[9]), .B1(d_out_d_11__N_1874[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11489), .COUT(n11490));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_12.INIT0 = 16'h5666;
    defparam sub_78_add_2_12.INIT1 = 16'h5666;
    defparam sub_78_add_2_12.INJECT1_0 = "NO";
    defparam sub_78_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_10 (.A0(d_out_d_11__N_1892[6]), .B0(d_out_d_11__N_1880[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[7]), .B1(d_out_d_11__N_1878[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11488), .COUT(n11489));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_10.INIT0 = 16'h5666;
    defparam sub_78_add_2_10.INIT1 = 16'h5666;
    defparam sub_78_add_2_10.INJECT1_0 = "NO";
    defparam sub_78_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_8 (.A0(d_out_d_11__N_1892[4]), .B0(d_out_d_11__N_1884[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[5]), .B1(d_out_d_11__N_1882[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11487), .COUT(n11488));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_8.INIT0 = 16'h5666;
    defparam sub_78_add_2_8.INIT1 = 16'h5666;
    defparam sub_78_add_2_8.INJECT1_0 = "NO";
    defparam sub_78_add_2_8.INJECT1_1 = "NO";
    FD1S3AX d_out_d__0_i2 (.D(d_out_d_11__N_1891), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[1]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i2.GSR = "ENABLED";
    CCU2D MultResult1_23__I_0_26 (.A0(MultResult1[23]), .B0(MultResult2[23]), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10951), .S0(ISquare_31__N_1895[24]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_26.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_26.INIT1 = 16'h0000;
    defparam MultResult1_23__I_0_26.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_26.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_24 (.A0(MultResult1[22]), .B0(MultResult2[22]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[23]), .B1(MultResult2[23]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10950), .COUT(n10951), .S0(ISquare_31__N_1895[22]), 
          .S1(ISquare_31__N_1895[23]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_24.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_24.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_24.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_24.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_22 (.A0(MultResult1[20]), .B0(MultResult2[20]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[21]), .B1(MultResult2[21]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10949), .COUT(n10950), .S0(ISquare_31__N_1895[20]), 
          .S1(ISquare_31__N_1895[21]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_22.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_22.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_22.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_22.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_20 (.A0(MultResult1[18]), .B0(MultResult2[18]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[19]), .B1(MultResult2[19]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10948), .COUT(n10949), .S0(ISquare_31__N_1895[18]), 
          .S1(ISquare_31__N_1895[19]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_20.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_20.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_20.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_20.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_18 (.A0(MultResult1[16]), .B0(MultResult2[16]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[17]), .B1(MultResult2[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10947), .COUT(n10948), .S0(ISquare_31__N_1895[16]), 
          .S1(ISquare_31__N_1895[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_18.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_18.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_18.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_18.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_16 (.A0(MultResult1[14]), .B0(MultResult2[14]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[15]), .B1(MultResult2[15]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10946), .COUT(n10947), .S0(ISquare_31__N_1895[14]), 
          .S1(ISquare_31__N_1895[15]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_16.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_16.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_16.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_16.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_14 (.A0(MultResult1[12]), .B0(MultResult2[12]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[13]), .B1(MultResult2[13]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10945), .COUT(n10946), .S0(ISquare_31__N_1895[12]), 
          .S1(ISquare_31__N_1895[13]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_14.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_14.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_14.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_14.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_12 (.A0(MultResult1[10]), .B0(MultResult2[10]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[11]), .B1(MultResult2[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10944), .COUT(n10945), .S0(ISquare_31__N_1895[10]), 
          .S1(ISquare_31__N_1895[11]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_12.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_12.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_12.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_12.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_10 (.A0(MultResult1[8]), .B0(MultResult2[8]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[9]), .B1(MultResult2[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10943), .COUT(n10944), .S0(ISquare_31__N_1895[8]), 
          .S1(ISquare_31__N_1895[9]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_10.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_10.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_10.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_10.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_8 (.A0(MultResult1[6]), .B0(MultResult2[6]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[7]), .B1(MultResult2[7]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10942), .COUT(n10943), .S0(ISquare_31__N_1895[6]), 
          .S1(ISquare_31__N_1895[7]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_8.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_8.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_8.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_8.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_6 (.A0(MultResult1[4]), .B0(MultResult2[4]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[5]), .B1(MultResult2[5]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10941), .COUT(n10942), .S0(ISquare_31__N_1895[4]), 
          .S1(ISquare_31__N_1895[5]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_6.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_6.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_6.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_6.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_4 (.A0(MultResult1[2]), .B0(MultResult2[2]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[3]), .B1(MultResult2[3]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10940), .COUT(n10941), .S0(ISquare_31__N_1895[2]), 
          .S1(ISquare_31__N_1895[3]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_4.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_4.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_4.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_4.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_2 (.A0(MultResult1[0]), .B0(MultResult2[0]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[1]), .B1(MultResult2[1]), 
          .C1(GND_net), .D1(GND_net), .COUT(n10940), .S1(ISquare_31__N_1895[1]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_2.INIT0 = 16'h7000;
    defparam MultResult1_23__I_0_2.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_2.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_2.INJECT1_1 = "NO";
    CCU2D add_517_11 (.A0(d_out_d_11__N_1872[17]), .B0(d_out_d_11__N_1871), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1872[17]), .B1(d_out_d_11__N_1871), 
          .C1(GND_net), .D1(GND_net), .CIN(n10702), .S0(d_out_d_11__N_1874[7]), 
          .S1(d_out_d_11__N_1874[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_517_11.INIT0 = 16'h5666;
    defparam add_517_11.INIT1 = 16'h5666;
    defparam add_517_11.INJECT1_0 = "NO";
    defparam add_517_11.INJECT1_1 = "NO";
    CCU2D add_517_9 (.A0(ISquare[31]), .B0(d_out_d_11__N_1872[17]), .C0(d_out_d_11__N_1872[4]), 
          .D0(GND_net), .A1(d_out_d_11__N_1872[5]), .B1(d_out_d_11__N_1872[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10701), .COUT(n10702), .S0(d_out_d_11__N_1874[5]), 
          .S1(d_out_d_11__N_1874[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_517_9.INIT0 = 16'h6969;
    defparam add_517_9.INIT1 = 16'h5999;
    defparam add_517_9.INJECT1_0 = "NO";
    defparam add_517_9.INJECT1_1 = "NO";
    CCU2D add_517_7 (.A0(ISquare[31]), .B0(d_out_d_11__N_1872[17]), .C0(d_out_d_11__N_1872[2]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1872[17]), 
          .C1(d_out_d_11__N_1872[3]), .D1(GND_net), .CIN(n10700), .COUT(n10701), 
          .S0(d_out_d_11__N_1874[3]), .S1(d_out_d_11__N_1874[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_517_7.INIT0 = 16'h6969;
    defparam add_517_7.INIT1 = 16'h6969;
    defparam add_517_7.INJECT1_0 = "NO";
    defparam add_517_7.INJECT1_1 = "NO";
    CCU2D add_517_5 (.A0(n12154), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1872[1]), .B1(d_out_d_11__N_1872[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10699), .COUT(n10700), .S0(d_out_d_11__N_1874[1]), 
          .S1(d_out_d_11__N_1874[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_517_5.INIT0 = 16'h5aaa;
    defparam add_517_5.INIT1 = 16'h5999;
    defparam add_517_5.INJECT1_0 = "NO";
    defparam add_517_5.INJECT1_1 = "NO";
    CCU2D add_517_3 (.A0(ISquare[20]), .B0(d_out_d_11__N_1872[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10698), .COUT(n10699), .S1(d_out_d_11__N_1874[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_517_3.INIT0 = 16'h5666;
    defparam add_517_3.INIT1 = 16'h5555;
    defparam add_517_3.INJECT1_0 = "NO";
    defparam add_517_3.INJECT1_1 = "NO";
    CCU2D add_517_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1872[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n10698));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_517_1.INIT0 = 16'hF000;
    defparam add_517_1.INIT1 = 16'h0aaa;
    defparam add_517_1.INJECT1_0 = "NO";
    defparam add_517_1.INJECT1_1 = "NO";
    FD1S3AX d_out_d__0_i3 (.D(d_out_d_11__N_1889), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i3.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i4 (.D(d_out_d_11__N_1887), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[3]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i4.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i5 (.D(d_out_d_11__N_1885), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i5.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i6 (.D(d_out_d_11__N_1883), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[5]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i6.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i7 (.D(d_out_d_11__N_1881), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i7.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i8 (.D(d_out_d_11__N_1879), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[7]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i8.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i9 (.D(d_out_d_11__N_1877), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i9.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i10 (.D(d_out_d_11__N_1875), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[9]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i10.GSR = "ENABLED";
    CCU2D add_417_17 (.A0(d_out_d_11__N_1878[17]), .B0(d_out_d_11__N_1877), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1878[17]), .B1(d_out_d_11__N_1877), 
          .C1(GND_net), .D1(GND_net), .CIN(n12152), .S0(d_out_d_11__N_1880[13]), 
          .S1(d_out_d_11__N_1880[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_417_17.INIT0 = 16'h5666;
    defparam add_417_17.INIT1 = 16'h5666;
    defparam add_417_17.INJECT1_0 = "NO";
    defparam add_417_17.INJECT1_1 = "NO";
    CCU2D add_417_15 (.A0(d_out_d_11__N_1878[10]), .B0(d_out_d_11__N_1878[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1878[11]), .B1(d_out_d_11__N_1878[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12151), .COUT(n12152), .S0(d_out_d_11__N_1880[11]), 
          .S1(d_out_d_11__N_1880[12]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_417_15.INIT0 = 16'h5999;
    defparam add_417_15.INIT1 = 16'h5999;
    defparam add_417_15.INJECT1_0 = "NO";
    defparam add_417_15.INJECT1_1 = "NO";
    CCU2D add_417_13 (.A0(d_out_d_11__N_1878[8]), .B0(d_out_d_11__N_1878[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1878[9]), .B1(d_out_d_11__N_1878[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12150), .COUT(n12151), .S0(d_out_d_11__N_1880[9]), 
          .S1(d_out_d_11__N_1880[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_417_13.INIT0 = 16'h5999;
    defparam add_417_13.INIT1 = 16'h5999;
    defparam add_417_13.INJECT1_0 = "NO";
    defparam add_417_13.INJECT1_1 = "NO";
    CCU2D add_417_11 (.A0(ISquare[31]), .B0(d_out_d_11__N_1878[17]), .C0(d_out_d_11__N_1878[6]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1878[17]), 
          .C1(d_out_d_11__N_1878[7]), .D1(GND_net), .CIN(n12149), .COUT(n12150), 
          .S0(d_out_d_11__N_1880[7]), .S1(d_out_d_11__N_1880[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_417_11.INIT0 = 16'h6969;
    defparam add_417_11.INIT1 = 16'h6969;
    defparam add_417_11.INJECT1_0 = "NO";
    defparam add_417_11.INJECT1_1 = "NO";
    CCU2D add_417_9 (.A0(d_out_d_11__N_1878[4]), .B0(d_out_d_11__N_1878[17]), 
          .C0(GND_net), .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1878[17]), 
          .C1(d_out_d_11__N_1878[5]), .D1(GND_net), .CIN(n12148), .COUT(n12149), 
          .S0(d_out_d_11__N_1880[5]), .S1(d_out_d_11__N_1880[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_417_9.INIT0 = 16'h5999;
    defparam add_417_9.INIT1 = 16'h6969;
    defparam add_417_9.INJECT1_0 = "NO";
    defparam add_417_9.INJECT1_1 = "NO";
    CCU2D add_417_7 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1878[17]), 
          .C0(d_out_d_11__N_1878[2]), .D0(GND_net), .A1(d_out_d_11__N_1872[17]), 
          .B1(d_out_d_11__N_1878[17]), .C1(d_out_d_11__N_1878[3]), .D1(GND_net), 
          .CIN(n12147), .COUT(n12148), .S0(d_out_d_11__N_1880[3]), .S1(d_out_d_11__N_1880[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_417_7.INIT0 = 16'h9696;
    defparam add_417_7.INIT1 = 16'h9696;
    defparam add_417_7.INJECT1_0 = "NO";
    defparam add_417_7.INJECT1_1 = "NO";
    CCU2D add_417_5 (.A0(d_out_d_11__N_1878[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1876[17]), .B1(d_out_d_11__N_1878[17]), 
          .C1(d_out_d_11__N_1878[1]), .D1(GND_net), .CIN(n12146), .COUT(n12147), 
          .S0(d_out_d_11__N_1880[1]), .S1(d_out_d_11__N_1880[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_417_5.INIT0 = 16'h5aaa;
    defparam add_417_5.INIT1 = 16'h9696;
    defparam add_417_5.INJECT1_0 = "NO";
    defparam add_417_5.INJECT1_1 = "NO";
    CCU2D add_417_3 (.A0(ISquare[14]), .B0(d_out_d_11__N_1878[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12145), .COUT(n12146), .S1(d_out_d_11__N_1880[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_417_3.INIT0 = 16'h5666;
    defparam add_417_3.INIT1 = 16'h5555;
    defparam add_417_3.INJECT1_0 = "NO";
    defparam add_417_3.INJECT1_1 = "NO";
    CCU2D add_417_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1878[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n12145));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_417_1.INIT0 = 16'hF000;
    defparam add_417_1.INIT1 = 16'h0aaa;
    defparam add_417_1.INJECT1_0 = "NO";
    defparam add_417_1.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_6 (.A0(d_out_d_11__N_1892[2]), .B0(d_out_d_11__N_1888[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[3]), .B1(d_out_d_11__N_1886[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11486), .COUT(n11487));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_6.INIT0 = 16'h5666;
    defparam sub_78_add_2_6.INIT1 = 16'h5666;
    defparam sub_78_add_2_6.INJECT1_0 = "NO";
    defparam sub_78_add_2_6.INJECT1_1 = "NO";
    CCU2D add_144_17 (.A0(d_out_d_11__N_1892[14]), .B0(ISquare[31]), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1892[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12139), .S1(d_out_d_11__N_2353[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_144_17.INIT0 = 16'h5666;
    defparam add_144_17.INIT1 = 16'h5aaa;
    defparam add_144_17.INJECT1_0 = "NO";
    defparam add_144_17.INJECT1_1 = "NO";
    CCU2D add_144_15 (.A0(d_out_d_11__N_1892[12]), .B0(ISquare[31]), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1892[13]), .B1(ISquare[31]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12138), .COUT(n12139));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_144_15.INIT0 = 16'h5666;
    defparam add_144_15.INIT1 = 16'h5666;
    defparam add_144_15.INJECT1_0 = "NO";
    defparam add_144_15.INJECT1_1 = "NO";
    CCU2D add_144_13 (.A0(d_out_d_11__N_1892[10]), .B0(d_out_d_11__N_1872[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[11]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12137), .COUT(n12138));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_144_13.INIT0 = 16'h5999;
    defparam add_144_13.INIT1 = 16'h5aaa;
    defparam add_144_13.INJECT1_0 = "NO";
    defparam add_144_13.INJECT1_1 = "NO";
    CCU2D add_144_11 (.A0(d_out_d_11__N_1892[8]), .B0(d_out_d_11__N_1876[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[9]), .B1(d_out_d_11__N_1874[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12136), .COUT(n12137));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_144_11.INIT0 = 16'h5999;
    defparam add_144_11.INIT1 = 16'h5999;
    defparam add_144_11.INJECT1_0 = "NO";
    defparam add_144_11.INJECT1_1 = "NO";
    CCU2D add_144_9 (.A0(d_out_d_11__N_1892[6]), .B0(d_out_d_11__N_1880[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[7]), .B1(d_out_d_11__N_1878[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12135), .COUT(n12136));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_144_9.INIT0 = 16'h5999;
    defparam add_144_9.INIT1 = 16'h5999;
    defparam add_144_9.INJECT1_0 = "NO";
    defparam add_144_9.INJECT1_1 = "NO";
    CCU2D add_144_7 (.A0(d_out_d_11__N_1892[4]), .B0(d_out_d_11__N_1884[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[5]), .B1(d_out_d_11__N_1882[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12134), .COUT(n12135));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_144_7.INIT0 = 16'h5999;
    defparam add_144_7.INIT1 = 16'h5999;
    defparam add_144_7.INJECT1_0 = "NO";
    defparam add_144_7.INJECT1_1 = "NO";
    CCU2D add_144_5 (.A0(d_out_d_11__N_1892[2]), .B0(d_out_d_11__N_1888[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[3]), .B1(d_out_d_11__N_1886[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12133), .COUT(n12134));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_144_5.INIT0 = 16'h5999;
    defparam add_144_5.INIT1 = 16'h5999;
    defparam add_144_5.INJECT1_0 = "NO";
    defparam add_144_5.INJECT1_1 = "NO";
    CCU2D add_144_3 (.A0(d_out_d_11__N_1892[0]), .B0(d_out_d_11__N_1892[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[1]), .B1(d_out_d_11__N_1890[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12132), .COUT(n12133));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_144_3.INIT0 = 16'h5999;
    defparam add_144_3.INIT1 = 16'h5999;
    defparam add_144_3.INJECT1_0 = "NO";
    defparam add_144_3.INJECT1_1 = "NO";
    CCU2D add_144_1 (.A0(ISquare[0]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(ISquare[1]), .B1(d_out_d_11__N_1892[17]), .C1(GND_net), 
          .D1(GND_net), .COUT(n12132));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_144_1.INIT0 = 16'h5000;
    defparam add_144_1.INIT1 = 16'h5666;
    defparam add_144_1.INJECT1_0 = "NO";
    defparam add_144_1.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_4 (.A0(d_out_d_11__N_1892[0]), .B0(d_out_d_11__N_1892[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[1]), .B1(d_out_d_11__N_1890[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11485), .COUT(n11486));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_4.INIT0 = 16'h5666;
    defparam sub_78_add_2_4.INIT1 = 16'h5666;
    defparam sub_78_add_2_4.INJECT1_0 = "NO";
    defparam sub_78_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_2 (.A0(ISquare[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[1]), .B1(d_out_d_11__N_1892[17]), 
          .C1(GND_net), .D1(GND_net), .COUT(n11485));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_2.INIT0 = 16'h5000;
    defparam sub_78_add_2_2.INIT1 = 16'h5999;
    defparam sub_78_add_2_2.INJECT1_0 = "NO";
    defparam sub_78_add_2_2.INJECT1_1 = "NO";
    CCU2D add_577_19 (.A0(d_out_d_11__N_1886[14]), .B0(d_out_d_11__N_1886[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1886[15]), .B1(d_out_d_11__N_1886[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11465), .S0(d_out_d_11__N_1888[15]), 
          .S1(d_out_d_11__N_1888[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_577_19.INIT0 = 16'h5999;
    defparam add_577_19.INIT1 = 16'h5999;
    defparam add_577_19.INJECT1_0 = "NO";
    defparam add_577_19.INJECT1_1 = "NO";
    CCU2D add_577_17 (.A0(d_out_d_11__N_1886[12]), .B0(d_out_d_11__N_1886[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1886[13]), .B1(d_out_d_11__N_1886[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11464), .COUT(n11465), .S0(d_out_d_11__N_1888[13]), 
          .S1(d_out_d_11__N_1888[14]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_577_17.INIT0 = 16'h5999;
    defparam add_577_17.INIT1 = 16'h5999;
    defparam add_577_17.INJECT1_0 = "NO";
    defparam add_577_17.INJECT1_1 = "NO";
    CCU2D add_577_15 (.A0(ISquare[31]), .B0(d_out_d_11__N_1886[17]), .C0(d_out_d_11__N_1886[10]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1886[17]), 
          .C1(d_out_d_11__N_1886[11]), .D1(GND_net), .CIN(n11463), .COUT(n11464), 
          .S0(d_out_d_11__N_1888[11]), .S1(d_out_d_11__N_1888[12]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_577_15.INIT0 = 16'h6969;
    defparam add_577_15.INIT1 = 16'h6969;
    defparam add_577_15.INJECT1_0 = "NO";
    defparam add_577_15.INJECT1_1 = "NO";
    CCU2D add_577_13 (.A0(d_out_d_11__N_1886[8]), .B0(d_out_d_11__N_1886[17]), 
          .C0(GND_net), .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1886[17]), 
          .C1(d_out_d_11__N_1886[9]), .D1(GND_net), .CIN(n11462), .COUT(n11463), 
          .S0(d_out_d_11__N_1888[9]), .S1(d_out_d_11__N_1888[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_577_13.INIT0 = 16'h5999;
    defparam add_577_13.INIT1 = 16'h6969;
    defparam add_577_13.INJECT1_0 = "NO";
    defparam add_577_13.INJECT1_1 = "NO";
    CCU2D add_577_11 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1886[17]), 
          .C0(d_out_d_11__N_1886[6]), .D0(GND_net), .A1(d_out_d_11__N_1872[17]), 
          .B1(d_out_d_11__N_1886[17]), .C1(d_out_d_11__N_1886[7]), .D1(GND_net), 
          .CIN(n11461), .COUT(n11462), .S0(d_out_d_11__N_1888[7]), .S1(d_out_d_11__N_1888[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_577_11.INIT0 = 16'h9696;
    defparam add_577_11.INIT1 = 16'h9696;
    defparam add_577_11.INJECT1_0 = "NO";
    defparam add_577_11.INJECT1_1 = "NO";
    CCU2D add_577_9 (.A0(d_out_d_11__N_1878[17]), .B0(d_out_d_11__N_1886[17]), 
          .C0(d_out_d_11__N_1886[4]), .D0(GND_net), .A1(d_out_d_11__N_1876[17]), 
          .B1(d_out_d_11__N_1886[17]), .C1(d_out_d_11__N_1886[5]), .D1(GND_net), 
          .CIN(n11460), .COUT(n11461), .S0(d_out_d_11__N_1888[5]), .S1(d_out_d_11__N_1888[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_577_9.INIT0 = 16'h9696;
    defparam add_577_9.INIT1 = 16'h9696;
    defparam add_577_9.INJECT1_0 = "NO";
    defparam add_577_9.INJECT1_1 = "NO";
    CCU2D add_577_7 (.A0(d_out_d_11__N_1882[17]), .B0(d_out_d_11__N_1886[17]), 
          .C0(d_out_d_11__N_1886[2]), .D0(GND_net), .A1(d_out_d_11__N_1880[17]), 
          .B1(d_out_d_11__N_1886[17]), .C1(d_out_d_11__N_1886[3]), .D1(GND_net), 
          .CIN(n11459), .COUT(n11460), .S0(d_out_d_11__N_1888[3]), .S1(d_out_d_11__N_1888[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_577_7.INIT0 = 16'h9696;
    defparam add_577_7.INIT1 = 16'h9696;
    defparam add_577_7.INJECT1_0 = "NO";
    defparam add_577_7.INJECT1_1 = "NO";
    CCU2D add_577_5 (.A0(d_out_d_11__N_1886[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1884[17]), .B1(d_out_d_11__N_1886[17]), 
          .C1(d_out_d_11__N_1886[1]), .D1(GND_net), .CIN(n11458), .COUT(n11459), 
          .S0(d_out_d_11__N_1888[1]), .S1(d_out_d_11__N_1888[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_577_5.INIT0 = 16'h5aaa;
    defparam add_577_5.INIT1 = 16'h9696;
    defparam add_577_5.INJECT1_0 = "NO";
    defparam add_577_5.INJECT1_1 = "NO";
    CCU2D add_577_3 (.A0(ISquare[6]), .B0(d_out_d_11__N_1886[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11457), .COUT(n11458), .S1(d_out_d_11__N_1888[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_577_3.INIT0 = 16'h5666;
    defparam add_577_3.INIT1 = 16'h5555;
    defparam add_577_3.INJECT1_0 = "NO";
    defparam add_577_3.INJECT1_1 = "NO";
    CCU2D add_577_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1886[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n11457));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_577_1.INIT0 = 16'hF000;
    defparam add_577_1.INIT1 = 16'h0aaa;
    defparam add_577_1.INJECT1_0 = "NO";
    defparam add_577_1.INJECT1_1 = "NO";
    CCU2D add_497_19 (.A0(d_out_d_11__N_1880[17]), .B0(d_out_d_11__N_1879), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1880[17]), .B1(d_out_d_11__N_1879), 
          .C1(GND_net), .D1(GND_net), .CIN(n11361), .S0(d_out_d_11__N_1882[15]), 
          .S1(d_out_d_11__N_1882[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_497_19.INIT0 = 16'h5666;
    defparam add_497_19.INIT1 = 16'h5666;
    defparam add_497_19.INJECT1_0 = "NO";
    defparam add_497_19.INJECT1_1 = "NO";
    CCU2D add_497_17 (.A0(d_out_d_11__N_1880[12]), .B0(d_out_d_11__N_1880[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1880[13]), .B1(d_out_d_11__N_1880[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11360), .COUT(n11361), .S0(d_out_d_11__N_1882[13]), 
          .S1(d_out_d_11__N_1882[14]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_497_17.INIT0 = 16'h5999;
    defparam add_497_17.INIT1 = 16'h5999;
    defparam add_497_17.INJECT1_0 = "NO";
    defparam add_497_17.INJECT1_1 = "NO";
    CCU2D add_497_15 (.A0(d_out_d_11__N_1880[10]), .B0(d_out_d_11__N_1880[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1880[11]), .B1(d_out_d_11__N_1880[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11359), .COUT(n11360), .S0(d_out_d_11__N_1882[11]), 
          .S1(d_out_d_11__N_1882[12]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_497_15.INIT0 = 16'h5999;
    defparam add_497_15.INIT1 = 16'h5999;
    defparam add_497_15.INJECT1_0 = "NO";
    defparam add_497_15.INJECT1_1 = "NO";
    CCU2D add_497_13 (.A0(ISquare[31]), .B0(d_out_d_11__N_1880[17]), .C0(d_out_d_11__N_1880[8]), 
          .D0(GND_net), .A1(d_out_d_11__N_1880[9]), .B1(d_out_d_11__N_1880[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11358), .COUT(n11359), .S0(d_out_d_11__N_1882[9]), 
          .S1(d_out_d_11__N_1882[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_497_13.INIT0 = 16'h6969;
    defparam add_497_13.INIT1 = 16'h5999;
    defparam add_497_13.INJECT1_0 = "NO";
    defparam add_497_13.INJECT1_1 = "NO";
    CCU2D add_497_11 (.A0(ISquare[31]), .B0(d_out_d_11__N_1880[17]), .C0(d_out_d_11__N_1880[6]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1880[17]), 
          .C1(d_out_d_11__N_1880[7]), .D1(GND_net), .CIN(n11357), .COUT(n11358), 
          .S0(d_out_d_11__N_1882[7]), .S1(d_out_d_11__N_1882[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_497_11.INIT0 = 16'h6969;
    defparam add_497_11.INIT1 = 16'h6969;
    defparam add_497_11.INJECT1_0 = "NO";
    defparam add_497_11.INJECT1_1 = "NO";
    CCU2D add_497_9 (.A0(d_out_d_11__N_1872[17]), .B0(d_out_d_11__N_1880[17]), 
          .C0(d_out_d_11__N_1880[4]), .D0(GND_net), .A1(d_out_d_11__N_1880[5]), 
          .B1(d_out_d_11__N_1880[17]), .C1(GND_net), .D1(GND_net), .CIN(n11356), 
          .COUT(n11357), .S0(d_out_d_11__N_1882[5]), .S1(d_out_d_11__N_1882[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_497_9.INIT0 = 16'h9696;
    defparam add_497_9.INIT1 = 16'h5999;
    defparam add_497_9.INJECT1_0 = "NO";
    defparam add_497_9.INJECT1_1 = "NO";
    CCU2D add_497_7 (.A0(d_out_d_11__N_1876[17]), .B0(d_out_d_11__N_1880[17]), 
          .C0(d_out_d_11__N_1880[2]), .D0(GND_net), .A1(d_out_d_11__N_1874[17]), 
          .B1(d_out_d_11__N_1880[17]), .C1(d_out_d_11__N_1880[3]), .D1(GND_net), 
          .CIN(n11355), .COUT(n11356), .S0(d_out_d_11__N_1882[3]), .S1(d_out_d_11__N_1882[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_497_7.INIT0 = 16'h9696;
    defparam add_497_7.INIT1 = 16'h9696;
    defparam add_497_7.INJECT1_0 = "NO";
    defparam add_497_7.INJECT1_1 = "NO";
    CCU2D add_497_5 (.A0(d_out_d_11__N_1880[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1878[17]), .B1(d_out_d_11__N_1880[17]), 
          .C1(d_out_d_11__N_1880[1]), .D1(GND_net), .CIN(n11354), .COUT(n11355), 
          .S0(d_out_d_11__N_1882[1]), .S1(d_out_d_11__N_1882[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_497_5.INIT0 = 16'h5aaa;
    defparam add_497_5.INIT1 = 16'h9696;
    defparam add_497_5.INJECT1_0 = "NO";
    defparam add_497_5.INJECT1_1 = "NO";
    CCU2D add_497_3 (.A0(ISquare[12]), .B0(d_out_d_11__N_1880[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11353), .COUT(n11354), .S1(d_out_d_11__N_1882[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_497_3.INIT0 = 16'h5666;
    defparam add_497_3.INIT1 = 16'h5555;
    defparam add_497_3.INJECT1_0 = "NO";
    defparam add_497_3.INJECT1_1 = "NO";
    CCU2D add_497_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1880[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n11353));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_497_1.INIT0 = 16'hF000;
    defparam add_497_1.INIT1 = 16'h0aaa;
    defparam add_497_1.INJECT1_0 = "NO";
    defparam add_497_1.INJECT1_1 = "NO";
    CCU2D add_617_19 (.A0(d_out_d_11__N_1884[14]), .B0(d_out_d_11__N_1884[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1884[15]), .B1(d_out_d_11__N_1884[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12104), .S0(d_out_d_11__N_1886[15]), 
          .S1(d_out_d_11__N_1886[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_617_19.INIT0 = 16'h5999;
    defparam add_617_19.INIT1 = 16'h5999;
    defparam add_617_19.INJECT1_0 = "NO";
    defparam add_617_19.INJECT1_1 = "NO";
    CCU2D add_617_17 (.A0(d_out_d_11__N_1884[12]), .B0(d_out_d_11__N_1884[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1884[13]), .B1(d_out_d_11__N_1884[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12103), .COUT(n12104), .S0(d_out_d_11__N_1886[13]), 
          .S1(d_out_d_11__N_1886[14]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_617_17.INIT0 = 16'h5999;
    defparam add_617_17.INIT1 = 16'h5999;
    defparam add_617_17.INJECT1_0 = "NO";
    defparam add_617_17.INJECT1_1 = "NO";
    CCU2D add_617_15 (.A0(ISquare[31]), .B0(d_out_d_11__N_1884[17]), .C0(d_out_d_11__N_1884[10]), 
          .D0(GND_net), .A1(d_out_d_11__N_1884[11]), .B1(d_out_d_11__N_1884[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12102), .COUT(n12103), .S0(d_out_d_11__N_1886[11]), 
          .S1(d_out_d_11__N_1886[12]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_617_15.INIT0 = 16'h6969;
    defparam add_617_15.INIT1 = 16'h5999;
    defparam add_617_15.INJECT1_0 = "NO";
    defparam add_617_15.INJECT1_1 = "NO";
    CCU2D add_617_13 (.A0(ISquare[31]), .B0(d_out_d_11__N_1884[17]), .C0(d_out_d_11__N_1884[8]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1884[17]), 
          .C1(d_out_d_11__N_1884[9]), .D1(GND_net), .CIN(n12101), .COUT(n12102), 
          .S0(d_out_d_11__N_1886[9]), .S1(d_out_d_11__N_1886[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_617_13.INIT0 = 16'h6969;
    defparam add_617_13.INIT1 = 16'h6969;
    defparam add_617_13.INJECT1_0 = "NO";
    defparam add_617_13.INJECT1_1 = "NO";
    CCU2D add_617_11 (.A0(d_out_d_11__N_1872[17]), .B0(d_out_d_11__N_1884[17]), 
          .C0(d_out_d_11__N_1884[6]), .D0(GND_net), .A1(d_out_d_11__N_1884[7]), 
          .B1(d_out_d_11__N_1884[17]), .C1(GND_net), .D1(GND_net), .CIN(n12100), 
          .COUT(n12101), .S0(d_out_d_11__N_1886[7]), .S1(d_out_d_11__N_1886[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_617_11.INIT0 = 16'h9696;
    defparam add_617_11.INIT1 = 16'h5999;
    defparam add_617_11.INJECT1_0 = "NO";
    defparam add_617_11.INJECT1_1 = "NO";
    CCU2D add_617_9 (.A0(d_out_d_11__N_1876[17]), .B0(d_out_d_11__N_1884[17]), 
          .C0(d_out_d_11__N_1884[4]), .D0(GND_net), .A1(d_out_d_11__N_1874[17]), 
          .B1(d_out_d_11__N_1884[17]), .C1(d_out_d_11__N_1884[5]), .D1(GND_net), 
          .CIN(n12099), .COUT(n12100), .S0(d_out_d_11__N_1886[5]), .S1(d_out_d_11__N_1886[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_617_9.INIT0 = 16'h9696;
    defparam add_617_9.INIT1 = 16'h9696;
    defparam add_617_9.INJECT1_0 = "NO";
    defparam add_617_9.INJECT1_1 = "NO";
    CCU2D add_617_7 (.A0(d_out_d_11__N_1880[17]), .B0(d_out_d_11__N_1884[17]), 
          .C0(d_out_d_11__N_1884[2]), .D0(GND_net), .A1(d_out_d_11__N_1878[17]), 
          .B1(d_out_d_11__N_1884[17]), .C1(d_out_d_11__N_1884[3]), .D1(GND_net), 
          .CIN(n12098), .COUT(n12099), .S0(d_out_d_11__N_1886[3]), .S1(d_out_d_11__N_1886[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_617_7.INIT0 = 16'h9696;
    defparam add_617_7.INIT1 = 16'h9696;
    defparam add_617_7.INJECT1_0 = "NO";
    defparam add_617_7.INJECT1_1 = "NO";
    CCU2D add_617_5 (.A0(d_out_d_11__N_1884[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1882[17]), .B1(d_out_d_11__N_1884[17]), 
          .C1(d_out_d_11__N_1884[1]), .D1(GND_net), .CIN(n12097), .COUT(n12098), 
          .S0(d_out_d_11__N_1886[1]), .S1(d_out_d_11__N_1886[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_617_5.INIT0 = 16'h5aaa;
    defparam add_617_5.INIT1 = 16'h9696;
    defparam add_617_5.INJECT1_0 = "NO";
    defparam add_617_5.INJECT1_1 = "NO";
    CCU2D add_617_3 (.A0(ISquare[8]), .B0(d_out_d_11__N_1884[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12096), .COUT(n12097), .S1(d_out_d_11__N_1886[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_617_3.INIT0 = 16'h5666;
    defparam add_617_3.INIT1 = 16'h5555;
    defparam add_617_3.INJECT1_0 = "NO";
    defparam add_617_3.INJECT1_1 = "NO";
    CCU2D add_617_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1884[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n12096));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_617_1.INIT0 = 16'hF000;
    defparam add_617_1.INIT1 = 16'h0aaa;
    defparam add_617_1.INJECT1_0 = "NO";
    defparam add_617_1.INJECT1_1 = "NO";
    CCU2D add_657_19 (.A0(d_out_d_11__N_1882[14]), .B0(d_out_d_11__N_1882[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1882[15]), .B1(d_out_d_11__N_1882[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12090), .S0(d_out_d_11__N_1884[15]), 
          .S1(d_out_d_11__N_1884[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_657_19.INIT0 = 16'h5999;
    defparam add_657_19.INIT1 = 16'h5999;
    defparam add_657_19.INJECT1_0 = "NO";
    defparam add_657_19.INJECT1_1 = "NO";
    CCU2D add_657_17 (.A0(d_out_d_11__N_1882[12]), .B0(d_out_d_11__N_1882[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1882[13]), .B1(d_out_d_11__N_1882[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12089), .COUT(n12090), .S0(d_out_d_11__N_1884[13]), 
          .S1(d_out_d_11__N_1884[14]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_657_17.INIT0 = 16'h5999;
    defparam add_657_17.INIT1 = 16'h5999;
    defparam add_657_17.INJECT1_0 = "NO";
    defparam add_657_17.INJECT1_1 = "NO";
    CCU2D add_657_15 (.A0(d_out_d_11__N_1882[10]), .B0(d_out_d_11__N_1882[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1882[11]), .B1(d_out_d_11__N_1882[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12088), .COUT(n12089), .S0(d_out_d_11__N_1884[11]), 
          .S1(d_out_d_11__N_1884[12]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_657_15.INIT0 = 16'h5999;
    defparam add_657_15.INIT1 = 16'h5999;
    defparam add_657_15.INJECT1_0 = "NO";
    defparam add_657_15.INJECT1_1 = "NO";
    CCU2D add_657_13 (.A0(ISquare[31]), .B0(d_out_d_11__N_1882[17]), .C0(d_out_d_11__N_1882[8]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1882[17]), 
          .C1(d_out_d_11__N_1882[9]), .D1(GND_net), .CIN(n12087), .COUT(n12088), 
          .S0(d_out_d_11__N_1884[9]), .S1(d_out_d_11__N_1884[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_657_13.INIT0 = 16'h6969;
    defparam add_657_13.INIT1 = 16'h6969;
    defparam add_657_13.INJECT1_0 = "NO";
    defparam add_657_13.INJECT1_1 = "NO";
    CCU2D add_657_11 (.A0(d_out_d_11__N_1882[6]), .B0(d_out_d_11__N_1882[17]), 
          .C0(GND_net), .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1882[17]), 
          .C1(d_out_d_11__N_1882[7]), .D1(GND_net), .CIN(n12086), .COUT(n12087), 
          .S0(d_out_d_11__N_1884[7]), .S1(d_out_d_11__N_1884[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_657_11.INIT0 = 16'h5999;
    defparam add_657_11.INIT1 = 16'h6969;
    defparam add_657_11.INJECT1_0 = "NO";
    defparam add_657_11.INJECT1_1 = "NO";
    CCU2D add_657_9 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1882[17]), 
          .C0(d_out_d_11__N_1882[4]), .D0(GND_net), .A1(d_out_d_11__N_1872[17]), 
          .B1(d_out_d_11__N_1882[17]), .C1(d_out_d_11__N_1882[5]), .D1(GND_net), 
          .CIN(n12085), .COUT(n12086), .S0(d_out_d_11__N_1884[5]), .S1(d_out_d_11__N_1884[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_657_9.INIT0 = 16'h9696;
    defparam add_657_9.INIT1 = 16'h9696;
    defparam add_657_9.INJECT1_0 = "NO";
    defparam add_657_9.INJECT1_1 = "NO";
    CCU2D add_657_7 (.A0(d_out_d_11__N_1878[17]), .B0(d_out_d_11__N_1882[17]), 
          .C0(d_out_d_11__N_1882[2]), .D0(GND_net), .A1(d_out_d_11__N_1876[17]), 
          .B1(d_out_d_11__N_1882[17]), .C1(d_out_d_11__N_1882[3]), .D1(GND_net), 
          .CIN(n12084), .COUT(n12085), .S0(d_out_d_11__N_1884[3]), .S1(d_out_d_11__N_1884[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_657_7.INIT0 = 16'h9696;
    defparam add_657_7.INIT1 = 16'h9696;
    defparam add_657_7.INJECT1_0 = "NO";
    defparam add_657_7.INJECT1_1 = "NO";
    CCU2D add_657_5 (.A0(d_out_d_11__N_1882[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1880[17]), .B1(d_out_d_11__N_1882[17]), 
          .C1(d_out_d_11__N_1882[1]), .D1(GND_net), .CIN(n12083), .COUT(n12084), 
          .S0(d_out_d_11__N_1884[1]), .S1(d_out_d_11__N_1884[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_657_5.INIT0 = 16'h5aaa;
    defparam add_657_5.INIT1 = 16'h9696;
    defparam add_657_5.INJECT1_0 = "NO";
    defparam add_657_5.INJECT1_1 = "NO";
    CCU2D add_657_3 (.A0(ISquare[10]), .B0(d_out_d_11__N_1882[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12082), .COUT(n12083), .S1(d_out_d_11__N_1884[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_657_3.INIT0 = 16'h5666;
    defparam add_657_3.INIT1 = 16'h5555;
    defparam add_657_3.INJECT1_0 = "NO";
    defparam add_657_3.INJECT1_1 = "NO";
    CCU2D add_657_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1882[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n12082));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_657_1.INIT0 = 16'hF000;
    defparam add_657_1.INIT1 = 16'h0aaa;
    defparam add_657_1.INJECT1_0 = "NO";
    defparam add_657_1.INJECT1_1 = "NO";
    CCU2D add_537_19 (.A0(d_out_d_11__N_1890[14]), .B0(d_out_d_11__N_1890[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1890[15]), .B1(d_out_d_11__N_1890[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12076), .S0(d_out_d_11__N_1892[15]), 
          .S1(d_out_d_11__N_1892[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_537_19.INIT0 = 16'h5999;
    defparam add_537_19.INIT1 = 16'h5999;
    defparam add_537_19.INJECT1_0 = "NO";
    defparam add_537_19.INJECT1_1 = "NO";
    CCU2D add_537_17 (.A0(ISquare[31]), .B0(d_out_d_11__N_1890[17]), .C0(d_out_d_11__N_1890[12]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1890[17]), 
          .C1(d_out_d_11__N_1890[13]), .D1(GND_net), .CIN(n12075), .COUT(n12076), 
          .S0(d_out_d_11__N_1892[13]), .S1(d_out_d_11__N_1892[14]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_537_17.INIT0 = 16'h6969;
    defparam add_537_17.INIT1 = 16'h6969;
    defparam add_537_17.INJECT1_0 = "NO";
    defparam add_537_17.INJECT1_1 = "NO";
    CCU2D add_537_15 (.A0(d_out_d_11__N_1890[10]), .B0(d_out_d_11__N_1890[17]), 
          .C0(GND_net), .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1890[17]), 
          .C1(d_out_d_11__N_1890[11]), .D1(GND_net), .CIN(n12074), .COUT(n12075), 
          .S0(d_out_d_11__N_1892[11]), .S1(d_out_d_11__N_1892[12]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_537_15.INIT0 = 16'h5999;
    defparam add_537_15.INIT1 = 16'h6969;
    defparam add_537_15.INJECT1_0 = "NO";
    defparam add_537_15.INJECT1_1 = "NO";
    CCU2D add_537_13 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(d_out_d_11__N_1890[8]), .D0(GND_net), .A1(d_out_d_11__N_1872[17]), 
          .B1(d_out_d_11__N_1890[17]), .C1(d_out_d_11__N_1890[9]), .D1(GND_net), 
          .CIN(n12073), .COUT(n12074), .S0(d_out_d_11__N_1892[9]), .S1(d_out_d_11__N_1892[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_537_13.INIT0 = 16'h9696;
    defparam add_537_13.INIT1 = 16'h9696;
    defparam add_537_13.INJECT1_0 = "NO";
    defparam add_537_13.INJECT1_1 = "NO";
    CCU2D add_537_11 (.A0(d_out_d_11__N_1878[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(d_out_d_11__N_1890[6]), .D0(GND_net), .A1(d_out_d_11__N_1876[17]), 
          .B1(d_out_d_11__N_1890[17]), .C1(d_out_d_11__N_1890[7]), .D1(GND_net), 
          .CIN(n12072), .COUT(n12073), .S0(d_out_d_11__N_1892[7]), .S1(d_out_d_11__N_1892[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_537_11.INIT0 = 16'h9696;
    defparam add_537_11.INIT1 = 16'h9696;
    defparam add_537_11.INJECT1_0 = "NO";
    defparam add_537_11.INJECT1_1 = "NO";
    CCU2D add_537_9 (.A0(d_out_d_11__N_1882[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(d_out_d_11__N_1890[4]), .D0(GND_net), .A1(d_out_d_11__N_1880[17]), 
          .B1(d_out_d_11__N_1890[17]), .C1(d_out_d_11__N_1890[5]), .D1(GND_net), 
          .CIN(n12071), .COUT(n12072), .S0(d_out_d_11__N_1892[5]), .S1(d_out_d_11__N_1892[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_537_9.INIT0 = 16'h9696;
    defparam add_537_9.INIT1 = 16'h9696;
    defparam add_537_9.INJECT1_0 = "NO";
    defparam add_537_9.INJECT1_1 = "NO";
    CCU2D add_537_7 (.A0(d_out_d_11__N_1886[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(d_out_d_11__N_1890[2]), .D0(GND_net), .A1(d_out_d_11__N_1884[17]), 
          .B1(d_out_d_11__N_1890[17]), .C1(d_out_d_11__N_1890[3]), .D1(GND_net), 
          .CIN(n12070), .COUT(n12071), .S0(d_out_d_11__N_1892[3]), .S1(d_out_d_11__N_1892[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_537_7.INIT0 = 16'h9696;
    defparam add_537_7.INIT1 = 16'h9696;
    defparam add_537_7.INJECT1_0 = "NO";
    defparam add_537_7.INJECT1_1 = "NO";
    CCU2D add_537_5 (.A0(d_out_d_11__N_1890[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1888[17]), .B1(d_out_d_11__N_1890[17]), 
          .C1(d_out_d_11__N_1890[1]), .D1(GND_net), .CIN(n12069), .COUT(n12070), 
          .S0(d_out_d_11__N_1892[1]), .S1(d_out_d_11__N_1892[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_537_5.INIT0 = 16'h5aaa;
    defparam add_537_5.INIT1 = 16'h9696;
    defparam add_537_5.INJECT1_0 = "NO";
    defparam add_537_5.INJECT1_1 = "NO";
    CCU2D add_537_3 (.A0(ISquare[2]), .B0(d_out_d_11__N_1890[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12068), .COUT(n12069), .S1(d_out_d_11__N_1892[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_537_3.INIT0 = 16'h5666;
    defparam add_537_3.INIT1 = 16'h5555;
    defparam add_537_3.INJECT1_0 = "NO";
    defparam add_537_3.INJECT1_1 = "NO";
    CCU2D add_537_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1890[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n12068));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_537_1.INIT0 = 16'hF000;
    defparam add_537_1.INIT1 = 16'h0aaa;
    defparam add_537_1.INJECT1_0 = "NO";
    defparam add_537_1.INJECT1_1 = "NO";
    CCU2D add_557_19 (.A0(d_out_d_11__N_1888[14]), .B0(d_out_d_11__N_1888[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1888[15]), .B1(d_out_d_11__N_1888[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12062), .S0(d_out_d_11__N_1890[15]), 
          .S1(d_out_d_11__N_1890[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_557_19.INIT0 = 16'h5999;
    defparam add_557_19.INIT1 = 16'h5999;
    defparam add_557_19.INJECT1_0 = "NO";
    defparam add_557_19.INJECT1_1 = "NO";
    CCU2D add_557_17 (.A0(ISquare[31]), .B0(d_out_d_11__N_1888[17]), .C0(d_out_d_11__N_1888[12]), 
          .D0(GND_net), .A1(d_out_d_11__N_1888[13]), .B1(d_out_d_11__N_1888[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12061), .COUT(n12062), .S0(d_out_d_11__N_1890[13]), 
          .S1(d_out_d_11__N_1890[14]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_557_17.INIT0 = 16'h6969;
    defparam add_557_17.INIT1 = 16'h5999;
    defparam add_557_17.INJECT1_0 = "NO";
    defparam add_557_17.INJECT1_1 = "NO";
    CCU2D add_557_15 (.A0(ISquare[31]), .B0(d_out_d_11__N_1888[17]), .C0(d_out_d_11__N_1888[10]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1888[17]), 
          .C1(d_out_d_11__N_1888[11]), .D1(GND_net), .CIN(n12060), .COUT(n12061), 
          .S0(d_out_d_11__N_1890[11]), .S1(d_out_d_11__N_1890[12]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_557_15.INIT0 = 16'h6969;
    defparam add_557_15.INIT1 = 16'h6969;
    defparam add_557_15.INJECT1_0 = "NO";
    defparam add_557_15.INJECT1_1 = "NO";
    CCU2D add_557_13 (.A0(d_out_d_11__N_1872[17]), .B0(d_out_d_11__N_1888[17]), 
          .C0(d_out_d_11__N_1888[8]), .D0(GND_net), .A1(d_out_d_11__N_1888[9]), 
          .B1(d_out_d_11__N_1888[17]), .C1(GND_net), .D1(GND_net), .CIN(n12059), 
          .COUT(n12060), .S0(d_out_d_11__N_1890[9]), .S1(d_out_d_11__N_1890[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_557_13.INIT0 = 16'h9696;
    defparam add_557_13.INIT1 = 16'h5999;
    defparam add_557_13.INJECT1_0 = "NO";
    defparam add_557_13.INJECT1_1 = "NO";
    CCU2D add_557_11 (.A0(d_out_d_11__N_1876[17]), .B0(d_out_d_11__N_1888[17]), 
          .C0(d_out_d_11__N_1888[6]), .D0(GND_net), .A1(d_out_d_11__N_1874[17]), 
          .B1(d_out_d_11__N_1888[17]), .C1(d_out_d_11__N_1888[7]), .D1(GND_net), 
          .CIN(n12058), .COUT(n12059), .S0(d_out_d_11__N_1890[7]), .S1(d_out_d_11__N_1890[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_557_11.INIT0 = 16'h9696;
    defparam add_557_11.INIT1 = 16'h9696;
    defparam add_557_11.INJECT1_0 = "NO";
    defparam add_557_11.INJECT1_1 = "NO";
    CCU2D add_557_9 (.A0(d_out_d_11__N_1880[17]), .B0(d_out_d_11__N_1888[17]), 
          .C0(d_out_d_11__N_1888[4]), .D0(GND_net), .A1(d_out_d_11__N_1878[17]), 
          .B1(d_out_d_11__N_1888[17]), .C1(d_out_d_11__N_1888[5]), .D1(GND_net), 
          .CIN(n12057), .COUT(n12058), .S0(d_out_d_11__N_1890[5]), .S1(d_out_d_11__N_1890[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_557_9.INIT0 = 16'h9696;
    defparam add_557_9.INIT1 = 16'h9696;
    defparam add_557_9.INJECT1_0 = "NO";
    defparam add_557_9.INJECT1_1 = "NO";
    CCU2D add_557_7 (.A0(d_out_d_11__N_1884[17]), .B0(d_out_d_11__N_1888[17]), 
          .C0(d_out_d_11__N_1888[2]), .D0(GND_net), .A1(d_out_d_11__N_1882[17]), 
          .B1(d_out_d_11__N_1888[17]), .C1(d_out_d_11__N_1888[3]), .D1(GND_net), 
          .CIN(n12056), .COUT(n12057), .S0(d_out_d_11__N_1890[3]), .S1(d_out_d_11__N_1890[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_557_7.INIT0 = 16'h9696;
    defparam add_557_7.INIT1 = 16'h9696;
    defparam add_557_7.INJECT1_0 = "NO";
    defparam add_557_7.INJECT1_1 = "NO";
    CCU2D add_557_5 (.A0(d_out_d_11__N_1888[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1886[17]), .B1(d_out_d_11__N_1888[17]), 
          .C1(d_out_d_11__N_1888[1]), .D1(GND_net), .CIN(n12055), .COUT(n12056), 
          .S0(d_out_d_11__N_1890[1]), .S1(d_out_d_11__N_1890[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_557_5.INIT0 = 16'h5aaa;
    defparam add_557_5.INIT1 = 16'h9696;
    defparam add_557_5.INJECT1_0 = "NO";
    defparam add_557_5.INJECT1_1 = "NO";
    CCU2D add_557_3 (.A0(ISquare[4]), .B0(d_out_d_11__N_1888[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12054), .COUT(n12055), .S1(d_out_d_11__N_1890[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_557_3.INIT0 = 16'h5666;
    defparam add_557_3.INIT1 = 16'h5555;
    defparam add_557_3.INJECT1_0 = "NO";
    defparam add_557_3.INJECT1_1 = "NO";
    LUT4 i1335_1_lut (.A(ISquare[31]), .Z(n209)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1335_1_lut.init = 16'h5555;
    CCU2D add_557_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1888[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n12054));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_557_1.INIT0 = 16'hF000;
    defparam add_557_1.INIT1 = 16'h0aaa;
    defparam add_557_1.INJECT1_0 = "NO";
    defparam add_557_1.INJECT1_1 = "NO";
    CCU2D add_437_15 (.A0(d_out_d_11__N_1876[17]), .B0(d_out_d_11__N_1875), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1876[17]), .B1(d_out_d_11__N_1875), 
          .C1(GND_net), .D1(GND_net), .CIN(n12048), .S0(d_out_d_11__N_1878[11]), 
          .S1(d_out_d_11__N_1878[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_437_15.INIT0 = 16'h5666;
    defparam add_437_15.INIT1 = 16'h5666;
    defparam add_437_15.INJECT1_0 = "NO";
    defparam add_437_15.INJECT1_1 = "NO";
    CCU2D add_437_13 (.A0(d_out_d_11__N_1876[8]), .B0(d_out_d_11__N_1876[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1876[9]), .B1(d_out_d_11__N_1876[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12047), .COUT(n12048), .S0(d_out_d_11__N_1878[9]), 
          .S1(d_out_d_11__N_1878[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_437_13.INIT0 = 16'h5999;
    defparam add_437_13.INIT1 = 16'h5999;
    defparam add_437_13.INJECT1_0 = "NO";
    defparam add_437_13.INJECT1_1 = "NO";
    CCU2D add_437_11 (.A0(ISquare[31]), .B0(d_out_d_11__N_1876[17]), .C0(d_out_d_11__N_1876[6]), 
          .D0(GND_net), .A1(d_out_d_11__N_1876[7]), .B1(d_out_d_11__N_1876[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12046), .COUT(n12047), .S0(d_out_d_11__N_1878[7]), 
          .S1(d_out_d_11__N_1878[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_437_11.INIT0 = 16'h6969;
    defparam add_437_11.INIT1 = 16'h5999;
    defparam add_437_11.INJECT1_0 = "NO";
    defparam add_437_11.INJECT1_1 = "NO";
    CCU2D add_437_9 (.A0(ISquare[31]), .B0(d_out_d_11__N_1876[17]), .C0(d_out_d_11__N_1876[4]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1876[17]), 
          .C1(d_out_d_11__N_1876[5]), .D1(GND_net), .CIN(n12045), .COUT(n12046), 
          .S0(d_out_d_11__N_1878[5]), .S1(d_out_d_11__N_1878[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_437_9.INIT0 = 16'h6969;
    defparam add_437_9.INIT1 = 16'h6969;
    defparam add_437_9.INJECT1_0 = "NO";
    defparam add_437_9.INJECT1_1 = "NO";
    CCU2D add_437_7 (.A0(d_out_d_11__N_1872[17]), .B0(d_out_d_11__N_1876[17]), 
          .C0(d_out_d_11__N_1876[2]), .D0(GND_net), .A1(d_out_d_11__N_1876[3]), 
          .B1(d_out_d_11__N_1876[17]), .C1(GND_net), .D1(GND_net), .CIN(n12044), 
          .COUT(n12045), .S0(d_out_d_11__N_1878[3]), .S1(d_out_d_11__N_1878[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_437_7.INIT0 = 16'h9696;
    defparam add_437_7.INIT1 = 16'h5999;
    defparam add_437_7.INJECT1_0 = "NO";
    defparam add_437_7.INJECT1_1 = "NO";
    CCU2D add_437_5 (.A0(d_out_d_11__N_1876[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1874[17]), .B1(d_out_d_11__N_1876[17]), 
          .C1(d_out_d_11__N_1876[1]), .D1(GND_net), .CIN(n12043), .COUT(n12044), 
          .S0(d_out_d_11__N_1878[1]), .S1(d_out_d_11__N_1878[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_437_5.INIT0 = 16'h5aaa;
    defparam add_437_5.INIT1 = 16'h9696;
    defparam add_437_5.INJECT1_0 = "NO";
    defparam add_437_5.INJECT1_1 = "NO";
    LUT4 d_out_d_11__I_10_1_lut (.A(d_out_d_11__N_1892[17]), .Z(d_out_d_11__N_1891)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_10_1_lut.init = 16'h5555;
    CCU2D add_437_3 (.A0(ISquare[16]), .B0(d_out_d_11__N_1876[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12042), .COUT(n12043), .S1(d_out_d_11__N_1878[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_437_3.INIT0 = 16'h5666;
    defparam add_437_3.INIT1 = 16'h5555;
    defparam add_437_3.INJECT1_0 = "NO";
    defparam add_437_3.INJECT1_1 = "NO";
    CCU2D add_437_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1876[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n12042));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_437_1.INIT0 = 16'hF000;
    defparam add_437_1.INIT1 = 16'h0aaa;
    defparam add_437_1.INJECT1_0 = "NO";
    defparam add_437_1.INJECT1_1 = "NO";
    Multiplier Multiplier2 (.CIC1_out_clkSin(CIC1_out_clkSin), .VCC_net(VCC_net), 
            .GND_net(GND_net), .MultDataC({MultDataC}), .MultResult2({MultResult2})) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    Multiplier_U0 Multiplier1 (.CIC1_out_clkSin(CIC1_out_clkSin), .VCC_net(VCC_net), 
            .GND_net(GND_net), .MultDataB({MultDataB}), .MultResult1({MultResult1})) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    
endmodule
//
// Verilog Description of module Multiplier
//

module Multiplier (CIC1_out_clkSin, VCC_net, GND_net, MultDataC, MultResult2) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input CIC1_out_clkSin;
    input VCC_net;
    input GND_net;
    input [11:0]MultDataC;
    output [23:0]MultResult2;
    
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(85[6:21])
    
    wire Multiplier_0_mult_0_5_n1, regb_b_1, rega_a_11, Multiplier_0_pp_1_2, 
        regb_b_2, regb_b_0, Multiplier_0_mult_2_5_n1, regb_b_3, Multiplier_0_pp_2_4, 
        regb_b_4, Multiplier_0_mult_4_5_n1, regb_b_5, Multiplier_0_pp_3_6, 
        regb_b_6, Multiplier_0_mult_6_5_n1, regb_b_7, Multiplier_0_pp_4_8, 
        regb_b_8, Multiplier_0_mult_8_5_n1, regb_b_9, Multiplier_0_pp_5_10, 
        regb_b_10, Multiplier_0_mult_10_0_n0, regb_b_11, Multiplier_0_mult_10_1_n1, 
        rega_a_3, rega_a_2, Multiplier_0_mult_10_1_n0, Multiplier_0_mult_10_2_n1, 
        rega_a_5, rega_a_4, Multiplier_0_mult_10_2_n0, Multiplier_0_mult_10_3_n1, 
        rega_a_7, rega_a_6, Multiplier_0_mult_10_3_n0, Multiplier_0_mult_10_4_n1, 
        rega_a_9, rega_a_8, Multiplier_0_mult_10_4_n0, Multiplier_0_mult_10_5_n2, 
        rega_a_10, Multiplier_0_mult_10_5_n0, rega_a_1, rego_o_0, rego_o_1, 
        rego_o_2, rego_o_3, rego_o_4, rego_o_5, rego_o_6, rego_o_7, 
        rego_o_8, rego_o_9, rego_o_10, rego_o_11, rego_o_12, rego_o_13, 
        rego_o_14, rego_o_15, rego_o_16, rego_o_17, rego_o_18, rego_o_19, 
        rego_o_20, rego_o_21, rego_o_22, rego_o_23, Multiplier_0_pp_0_0, 
        Multiplier_0_pp_0_1, s_Multiplier_0_0_2, s_Multiplier_0_0_3, s_Multiplier_0_0_4, 
        f_s_Multiplier_0_0_4, s_Multiplier_0_0_5, f_s_Multiplier_0_0_5, 
        s_Multiplier_0_0_6, f_s_Multiplier_0_0_6, s_Multiplier_0_0_7, 
        f_s_Multiplier_0_0_7, s_Multiplier_0_0_8, f_s_Multiplier_0_0_8, 
        s_Multiplier_0_0_9, f_s_Multiplier_0_0_9, s_Multiplier_0_0_10, 
        f_s_Multiplier_0_0_10, s_Multiplier_0_0_11, f_s_Multiplier_0_0_11, 
        s_Multiplier_0_0_12, f_s_Multiplier_0_0_12, s_Multiplier_0_0_13, 
        f_s_Multiplier_0_0_13, s_Multiplier_0_0_14, f_s_Multiplier_0_0_14, 
        s_Multiplier_0_0_15, f_s_Multiplier_0_0_15, s_Multiplier_0_0_16, 
        f_s_Multiplier_0_0_16, s_Multiplier_0_0_17, f_s_Multiplier_0_0_17, 
        f_Multiplier_0_pp_2_4, f_Multiplier_0_pp_2_5, Multiplier_0_pp_2_5, 
        s_Multiplier_0_1_6, f_s_Multiplier_0_1_6, s_Multiplier_0_1_7, 
        f_s_Multiplier_0_1_7, s_Multiplier_0_1_8, f_s_Multiplier_0_1_8, 
        s_Multiplier_0_1_9, f_s_Multiplier_0_1_9, s_Multiplier_0_1_10, 
        f_s_Multiplier_0_1_10, s_Multiplier_0_1_11, f_s_Multiplier_0_1_11, 
        s_Multiplier_0_1_12, f_s_Multiplier_0_1_12, s_Multiplier_0_1_13, 
        f_s_Multiplier_0_1_13, s_Multiplier_0_1_14, f_s_Multiplier_0_1_14, 
        s_Multiplier_0_1_15, f_s_Multiplier_0_1_15, s_Multiplier_0_1_16, 
        f_s_Multiplier_0_1_16, s_Multiplier_0_1_17, f_s_Multiplier_0_1_17, 
        s_Multiplier_0_1_18, f_s_Multiplier_0_1_18, s_Multiplier_0_1_19, 
        f_s_Multiplier_0_1_19, s_Multiplier_0_1_20, f_s_Multiplier_0_1_20, 
        s_Multiplier_0_1_21, f_s_Multiplier_0_1_21, f_Multiplier_0_pp_4_8, 
        f_Multiplier_0_pp_4_9, Multiplier_0_pp_4_9, s_Multiplier_0_2_10, 
        f_s_Multiplier_0_2_10, s_Multiplier_0_2_11, f_s_Multiplier_0_2_11, 
        s_Multiplier_0_2_12, f_s_Multiplier_0_2_12, s_Multiplier_0_2_13, 
        f_s_Multiplier_0_2_13, s_Multiplier_0_2_14, f_s_Multiplier_0_2_14, 
        s_Multiplier_0_2_15, f_s_Multiplier_0_2_15, s_Multiplier_0_2_16, 
        f_s_Multiplier_0_2_16, s_Multiplier_0_2_17, f_s_Multiplier_0_2_17, 
        s_Multiplier_0_2_18, f_s_Multiplier_0_2_18, s_Multiplier_0_2_19, 
        f_s_Multiplier_0_2_19, s_Multiplier_0_2_20, f_s_Multiplier_0_2_20, 
        s_Multiplier_0_2_21, f_s_Multiplier_0_2_21, s_Multiplier_0_2_22, 
        f_s_Multiplier_0_2_22, s_Multiplier_0_2_23, f_s_Multiplier_0_2_23, 
        Multiplier_0_cin_lr_0, Multiplier_0_pp_0_13, mfco, Multiplier_0_cin_lr_2, 
        Multiplier_0_pp_1_15, mfco_1, Multiplier_0_cin_lr_4, Multiplier_0_pp_2_17, 
        mfco_2, Multiplier_0_cin_lr_6, Multiplier_0_pp_3_19, mfco_3, 
        Multiplier_0_cin_lr_8, Multiplier_0_pp_4_21, mfco_4, Multiplier_0_cin_lr_10, 
        Multiplier_0_pp_5_23, mfco_5, co_Multiplier_0_0_1, Multiplier_0_pp_0_2, 
        co_Multiplier_0_0_2, Multiplier_0_pp_0_4, Multiplier_0_pp_0_3, 
        Multiplier_0_pp_1_4, Multiplier_0_pp_1_3, co_Multiplier_0_0_3, 
        Multiplier_0_pp_0_6, Multiplier_0_pp_0_5, Multiplier_0_pp_1_6, 
        Multiplier_0_pp_1_5, co_Multiplier_0_0_4, Multiplier_0_pp_0_8, 
        Multiplier_0_pp_0_7, Multiplier_0_pp_1_8, Multiplier_0_pp_1_7, 
        co_Multiplier_0_0_5, Multiplier_0_pp_0_10, Multiplier_0_pp_0_9, 
        Multiplier_0_pp_1_10, Multiplier_0_pp_1_9, co_Multiplier_0_0_6, 
        Multiplier_0_pp_0_12, Multiplier_0_pp_0_11, Multiplier_0_pp_1_12, 
        Multiplier_0_pp_1_11, co_Multiplier_0_0_7, Multiplier_0_pp_1_14, 
        Multiplier_0_pp_1_13, co_Multiplier_0_0_8, co_Multiplier_0_1_1, 
        Multiplier_0_pp_2_6, co_Multiplier_0_1_2, Multiplier_0_pp_2_8, 
        Multiplier_0_pp_2_7, Multiplier_0_pp_3_8, Multiplier_0_pp_3_7, 
        co_Multiplier_0_1_3, Multiplier_0_pp_2_10, Multiplier_0_pp_2_9, 
        Multiplier_0_pp_3_10, Multiplier_0_pp_3_9, co_Multiplier_0_1_4, 
        Multiplier_0_pp_2_12, Multiplier_0_pp_2_11, Multiplier_0_pp_3_12, 
        Multiplier_0_pp_3_11, co_Multiplier_0_1_5, Multiplier_0_pp_2_14, 
        Multiplier_0_pp_2_13, Multiplier_0_pp_3_14, Multiplier_0_pp_3_13, 
        co_Multiplier_0_1_6, Multiplier_0_pp_2_16, Multiplier_0_pp_2_15, 
        Multiplier_0_pp_3_16, Multiplier_0_pp_3_15, co_Multiplier_0_1_7, 
        Multiplier_0_pp_3_18, Multiplier_0_pp_3_17, co_Multiplier_0_1_8, 
        co_Multiplier_0_2_1, Multiplier_0_pp_4_10, co_Multiplier_0_2_2, 
        Multiplier_0_pp_4_12, Multiplier_0_pp_4_11, Multiplier_0_pp_5_12, 
        Multiplier_0_pp_5_11, co_Multiplier_0_2_3, Multiplier_0_pp_4_14, 
        Multiplier_0_pp_4_13, Multiplier_0_pp_5_14, Multiplier_0_pp_5_13, 
        co_Multiplier_0_2_4, Multiplier_0_pp_4_16, Multiplier_0_pp_4_15, 
        Multiplier_0_pp_5_16, Multiplier_0_pp_5_15, co_Multiplier_0_2_5, 
        Multiplier_0_pp_4_18, Multiplier_0_pp_4_17, Multiplier_0_pp_5_18, 
        Multiplier_0_pp_5_17, co_Multiplier_0_2_6, Multiplier_0_pp_4_20, 
        Multiplier_0_pp_4_19, Multiplier_0_pp_5_20, Multiplier_0_pp_5_19, 
        co_Multiplier_0_2_7, Multiplier_0_pp_5_22, Multiplier_0_pp_5_21, 
        co_Multiplier_0_3_1, co_Multiplier_0_3_2, co_Multiplier_0_3_3, 
        s_Multiplier_0_3_8, co_Multiplier_0_3_4, s_Multiplier_0_3_9, s_Multiplier_0_3_10, 
        co_Multiplier_0_3_5, s_Multiplier_0_3_11, s_Multiplier_0_3_12, 
        co_Multiplier_0_3_6, s_Multiplier_0_3_13, s_Multiplier_0_3_14, 
        co_Multiplier_0_3_7, s_Multiplier_0_3_15, s_Multiplier_0_3_16, 
        co_Multiplier_0_3_8, s_Multiplier_0_3_17, s_Multiplier_0_3_18, 
        co_Multiplier_0_3_9, s_Multiplier_0_3_19, s_Multiplier_0_3_20, 
        co_Multiplier_0_3_10, s_Multiplier_0_3_21, s_Multiplier_0_3_22, 
        s_Multiplier_0_3_23, co_t_Multiplier_0_4_1, co_t_Multiplier_0_4_2, 
        co_t_Multiplier_0_4_3, co_t_Multiplier_0_4_4, co_t_Multiplier_0_4_5, 
        co_t_Multiplier_0_4_6, co_t_Multiplier_0_4_7, co_t_Multiplier_0_4_8, 
        mco, mco_1, mco_2, mco_3, mco_4, Multiplier_0_mult_0_5_n2, 
        mco_5, mco_6, mco_7, mco_8, mco_9, Multiplier_0_mult_2_5_n2, 
        mco_10, mco_11, mco_12, mco_13, mco_14, Multiplier_0_mult_4_5_n2, 
        mco_15, mco_16, mco_17, mco_18, mco_19, Multiplier_0_mult_6_5_n2, 
        mco_20, mco_21, mco_22, mco_23, mco_24, Multiplier_0_mult_8_5_n2, 
        Multiplier_0_mult_10_0_n1, mco_25, mco_26, mco_27, mco_28, 
        mco_29;
    
    ND2 ND2_t25 (.A(rega_a_11), .B(regb_b_1), .Z(Multiplier_0_mult_0_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    AND2 AND2_t24 (.A(regb_b_0), .B(regb_b_2), .Z(Multiplier_0_pp_1_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(382[10:72])
    ND2 ND2_t22 (.A(rega_a_11), .B(regb_b_3), .Z(Multiplier_0_mult_2_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    AND2 AND2_t21 (.A(regb_b_0), .B(regb_b_4), .Z(Multiplier_0_pp_2_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(388[10:72])
    ND2 ND2_t19 (.A(rega_a_11), .B(regb_b_5), .Z(Multiplier_0_mult_4_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    AND2 AND2_t18 (.A(regb_b_0), .B(regb_b_6), .Z(Multiplier_0_pp_3_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(394[10:72])
    ND2 ND2_t16 (.A(rega_a_11), .B(regb_b_7), .Z(Multiplier_0_mult_6_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    AND2 AND2_t15 (.A(regb_b_0), .B(regb_b_8), .Z(Multiplier_0_pp_4_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(400[10:72])
    ND2 ND2_t13 (.A(rega_a_11), .B(regb_b_9), .Z(Multiplier_0_mult_8_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    AND2 AND2_t12 (.A(regb_b_0), .B(regb_b_10), .Z(Multiplier_0_pp_5_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(406[10:74])
    ND2 ND2_t10 (.A(regb_b_0), .B(regb_b_11), .Z(Multiplier_0_mult_10_0_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t9 (.A(rega_a_3), .B(regb_b_11), .Z(Multiplier_0_mult_10_1_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t8 (.A(rega_a_2), .B(regb_b_11), .Z(Multiplier_0_mult_10_1_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t7 (.A(rega_a_5), .B(regb_b_11), .Z(Multiplier_0_mult_10_2_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t6 (.A(rega_a_4), .B(regb_b_11), .Z(Multiplier_0_mult_10_2_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t5 (.A(rega_a_7), .B(regb_b_11), .Z(Multiplier_0_mult_10_3_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t4 (.A(rega_a_6), .B(regb_b_11), .Z(Multiplier_0_mult_10_3_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t3 (.A(rega_a_9), .B(regb_b_11), .Z(Multiplier_0_mult_10_4_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t2 (.A(rega_a_8), .B(regb_b_11), .Z(Multiplier_0_mult_10_4_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t1 (.A(rega_a_11), .B(regb_b_10), .Z(Multiplier_0_mult_10_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t0 (.A(rega_a_10), .B(regb_b_11), .Z(Multiplier_0_mult_10_5_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FD1P3DX FF_98 (.D(MultDataC[1]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(435[13:82])
    defparam FF_98.GSR = "ENABLED";
    FD1P3DX FF_97 (.D(MultDataC[2]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(438[13:82])
    defparam FF_97.GSR = "ENABLED";
    FD1P3DX FF_96 (.D(MultDataC[3]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(441[13:82])
    defparam FF_96.GSR = "ENABLED";
    FD1P3DX FF_95 (.D(MultDataC[4]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(444[13:82])
    defparam FF_95.GSR = "ENABLED";
    FD1P3DX FF_94 (.D(MultDataC[5]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(447[13:82])
    defparam FF_94.GSR = "ENABLED";
    FD1P3DX FF_93 (.D(MultDataC[6]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(450[13:82])
    defparam FF_93.GSR = "ENABLED";
    FD1P3DX FF_92 (.D(MultDataC[7]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(453[13:82])
    defparam FF_92.GSR = "ENABLED";
    FD1P3DX FF_91 (.D(MultDataC[8]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(456[13:82])
    defparam FF_91.GSR = "ENABLED";
    FD1P3DX FF_90 (.D(MultDataC[9]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(459[13:82])
    defparam FF_90.GSR = "ENABLED";
    FD1P3DX FF_89 (.D(MultDataC[10]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(462[13:84])
    defparam FF_89.GSR = "ENABLED";
    FD1P3DX FF_88 (.D(MultDataC[11]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(465[13:84])
    defparam FF_88.GSR = "ENABLED";
    FD1P3DX FF_87 (.D(MultDataC[0]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_0)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(468[13:82])
    defparam FF_87.GSR = "ENABLED";
    FD1P3DX FF_86 (.D(MultDataC[1]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(471[13:82])
    defparam FF_86.GSR = "ENABLED";
    FD1P3DX FF_85 (.D(MultDataC[2]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(474[13:82])
    defparam FF_85.GSR = "ENABLED";
    FD1P3DX FF_84 (.D(MultDataC[3]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(477[13:82])
    defparam FF_84.GSR = "ENABLED";
    FD1P3DX FF_83 (.D(MultDataC[4]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(480[13:82])
    defparam FF_83.GSR = "ENABLED";
    FD1P3DX FF_82 (.D(MultDataC[5]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(483[13:82])
    defparam FF_82.GSR = "ENABLED";
    FD1P3DX FF_81 (.D(MultDataC[6]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(486[13:82])
    defparam FF_81.GSR = "ENABLED";
    FD1P3DX FF_80 (.D(MultDataC[7]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(489[13:82])
    defparam FF_80.GSR = "ENABLED";
    FD1P3DX FF_79 (.D(MultDataC[8]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(492[13:82])
    defparam FF_79.GSR = "ENABLED";
    FD1P3DX FF_78 (.D(MultDataC[9]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(495[13:82])
    defparam FF_78.GSR = "ENABLED";
    FD1P3DX FF_77 (.D(MultDataC[10]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(498[13:84])
    defparam FF_77.GSR = "ENABLED";
    FD1P3DX FF_76 (.D(MultDataC[11]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(501[13:84])
    defparam FF_76.GSR = "ENABLED";
    FD1P3DX FF_75 (.D(rego_o_0), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[0])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(504[13:83])
    defparam FF_75.GSR = "ENABLED";
    FD1P3DX FF_74 (.D(rego_o_1), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[1])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(507[13:83])
    defparam FF_74.GSR = "ENABLED";
    FD1P3DX FF_73 (.D(rego_o_2), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[2])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(510[13:83])
    defparam FF_73.GSR = "ENABLED";
    FD1P3DX FF_72 (.D(rego_o_3), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[3])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(513[13:83])
    defparam FF_72.GSR = "ENABLED";
    FD1P3DX FF_71 (.D(rego_o_4), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[4])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(516[13:83])
    defparam FF_71.GSR = "ENABLED";
    FD1P3DX FF_70 (.D(rego_o_5), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[5])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(519[13:83])
    defparam FF_70.GSR = "ENABLED";
    FD1P3DX FF_69 (.D(rego_o_6), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[6])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(522[13:83])
    defparam FF_69.GSR = "ENABLED";
    FD1P3DX FF_68 (.D(rego_o_7), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[7])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(525[13:83])
    defparam FF_68.GSR = "ENABLED";
    FD1P3DX FF_67 (.D(rego_o_8), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[8])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(528[13:83])
    defparam FF_67.GSR = "ENABLED";
    FD1P3DX FF_66 (.D(rego_o_9), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[9])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(531[13:83])
    defparam FF_66.GSR = "ENABLED";
    FD1P3DX FF_65 (.D(rego_o_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[10])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(534[13:85])
    defparam FF_65.GSR = "ENABLED";
    FD1P3DX FF_64 (.D(rego_o_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[11])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(537[13:85])
    defparam FF_64.GSR = "ENABLED";
    FD1P3DX FF_63 (.D(rego_o_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[12])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(540[13:85])
    defparam FF_63.GSR = "ENABLED";
    FD1P3DX FF_62 (.D(rego_o_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[13])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(543[13:85])
    defparam FF_62.GSR = "ENABLED";
    FD1P3DX FF_61 (.D(rego_o_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[14])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(546[13:85])
    defparam FF_61.GSR = "ENABLED";
    FD1P3DX FF_60 (.D(rego_o_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[15])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(549[13:85])
    defparam FF_60.GSR = "ENABLED";
    FD1P3DX FF_59 (.D(rego_o_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[16])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(552[13:85])
    defparam FF_59.GSR = "ENABLED";
    FD1P3DX FF_58 (.D(rego_o_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[17])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(555[13:85])
    defparam FF_58.GSR = "ENABLED";
    FD1P3DX FF_57 (.D(rego_o_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[18])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(558[13:85])
    defparam FF_57.GSR = "ENABLED";
    FD1P3DX FF_56 (.D(rego_o_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[19])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(561[13:85])
    defparam FF_56.GSR = "ENABLED";
    FD1P3DX FF_55 (.D(rego_o_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[20])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(564[13:85])
    defparam FF_55.GSR = "ENABLED";
    FD1P3DX FF_54 (.D(rego_o_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[21])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(567[13:85])
    defparam FF_54.GSR = "ENABLED";
    FD1P3DX FF_53 (.D(rego_o_22), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[22])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(570[13:85])
    defparam FF_53.GSR = "ENABLED";
    FD1P3DX FF_52 (.D(rego_o_23), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[23])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(573[13:85])
    defparam FF_52.GSR = "ENABLED";
    FD1P3DX FF_51 (.D(Multiplier_0_pp_0_0), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_0)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(576[13] 577[35])
    defparam FF_51.GSR = "ENABLED";
    FD1P3DX FF_50 (.D(Multiplier_0_pp_0_1), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(580[13] 581[35])
    defparam FF_50.GSR = "ENABLED";
    FD1P3DX FF_49 (.D(s_Multiplier_0_0_2), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(584[13] 585[34])
    defparam FF_49.GSR = "ENABLED";
    FD1P3DX FF_48 (.D(s_Multiplier_0_0_3), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(588[13] 589[34])
    defparam FF_48.GSR = "ENABLED";
    FD1P3DX FF_47 (.D(s_Multiplier_0_0_4), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(592[13] 593[34])
    defparam FF_47.GSR = "ENABLED";
    FD1P3DX FF_46 (.D(s_Multiplier_0_0_5), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(596[13] 597[34])
    defparam FF_46.GSR = "ENABLED";
    FD1P3DX FF_45 (.D(s_Multiplier_0_0_6), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(600[13] 601[34])
    defparam FF_45.GSR = "ENABLED";
    FD1P3DX FF_44 (.D(s_Multiplier_0_0_7), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(604[13] 605[34])
    defparam FF_44.GSR = "ENABLED";
    FD1P3DX FF_43 (.D(s_Multiplier_0_0_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(608[13] 609[34])
    defparam FF_43.GSR = "ENABLED";
    FD1P3DX FF_42 (.D(s_Multiplier_0_0_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(612[13] 613[34])
    defparam FF_42.GSR = "ENABLED";
    FD1P3DX FF_41 (.D(s_Multiplier_0_0_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(616[13] 617[35])
    defparam FF_41.GSR = "ENABLED";
    FD1P3DX FF_40 (.D(s_Multiplier_0_0_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(620[13] 621[35])
    defparam FF_40.GSR = "ENABLED";
    FD1P3DX FF_39 (.D(s_Multiplier_0_0_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(624[13] 625[35])
    defparam FF_39.GSR = "ENABLED";
    FD1P3DX FF_38 (.D(s_Multiplier_0_0_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(628[13] 629[35])
    defparam FF_38.GSR = "ENABLED";
    FD1P3DX FF_37 (.D(s_Multiplier_0_0_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(632[13] 633[35])
    defparam FF_37.GSR = "ENABLED";
    FD1P3DX FF_36 (.D(s_Multiplier_0_0_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(636[13] 637[35])
    defparam FF_36.GSR = "ENABLED";
    FD1P3DX FF_35 (.D(s_Multiplier_0_0_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(640[13] 641[35])
    defparam FF_35.GSR = "ENABLED";
    FD1P3DX FF_34 (.D(s_Multiplier_0_0_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(644[13] 645[35])
    defparam FF_34.GSR = "ENABLED";
    FD1P3DX FF_33 (.D(Multiplier_0_pp_2_4), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_2_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(648[13] 649[35])
    defparam FF_33.GSR = "ENABLED";
    FD1P3DX FF_32 (.D(Multiplier_0_pp_2_5), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_2_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(652[13] 653[35])
    defparam FF_32.GSR = "ENABLED";
    FD1P3DX FF_31 (.D(s_Multiplier_0_1_6), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(656[13] 657[34])
    defparam FF_31.GSR = "ENABLED";
    FD1P3DX FF_30 (.D(s_Multiplier_0_1_7), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(660[13] 661[34])
    defparam FF_30.GSR = "ENABLED";
    FD1P3DX FF_29 (.D(s_Multiplier_0_1_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(664[13] 665[34])
    defparam FF_29.GSR = "ENABLED";
    FD1P3DX FF_28 (.D(s_Multiplier_0_1_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(668[13] 669[34])
    defparam FF_28.GSR = "ENABLED";
    FD1P3DX FF_27 (.D(s_Multiplier_0_1_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(672[13] 673[35])
    defparam FF_27.GSR = "ENABLED";
    FD1P3DX FF_26 (.D(s_Multiplier_0_1_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(676[13] 677[35])
    defparam FF_26.GSR = "ENABLED";
    FD1P3DX FF_25 (.D(s_Multiplier_0_1_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(680[13] 681[35])
    defparam FF_25.GSR = "ENABLED";
    FD1P3DX FF_24 (.D(s_Multiplier_0_1_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(684[13] 685[35])
    defparam FF_24.GSR = "ENABLED";
    FD1P3DX FF_23 (.D(s_Multiplier_0_1_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(688[13] 689[35])
    defparam FF_23.GSR = "ENABLED";
    FD1P3DX FF_22 (.D(s_Multiplier_0_1_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(692[13] 693[35])
    defparam FF_22.GSR = "ENABLED";
    FD1P3DX FF_21 (.D(s_Multiplier_0_1_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(696[13] 697[35])
    defparam FF_21.GSR = "ENABLED";
    FD1P3DX FF_20 (.D(s_Multiplier_0_1_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(700[13] 701[35])
    defparam FF_20.GSR = "ENABLED";
    FD1P3DX FF_19 (.D(s_Multiplier_0_1_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(704[13] 705[35])
    defparam FF_19.GSR = "ENABLED";
    FD1P3DX FF_18 (.D(s_Multiplier_0_1_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(708[13] 709[35])
    defparam FF_18.GSR = "ENABLED";
    FD1P3DX FF_17 (.D(s_Multiplier_0_1_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(712[13] 713[35])
    defparam FF_17.GSR = "ENABLED";
    FD1P3DX FF_16 (.D(s_Multiplier_0_1_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(716[13] 717[35])
    defparam FF_16.GSR = "ENABLED";
    FD1P3DX FF_15 (.D(Multiplier_0_pp_4_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_4_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(720[13] 721[35])
    defparam FF_15.GSR = "ENABLED";
    FD1P3DX FF_14 (.D(Multiplier_0_pp_4_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_4_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(724[13] 725[35])
    defparam FF_14.GSR = "ENABLED";
    FD1P3DX FF_13 (.D(s_Multiplier_0_2_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(728[13] 729[35])
    defparam FF_13.GSR = "ENABLED";
    FD1P3DX FF_12 (.D(s_Multiplier_0_2_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(732[13] 733[35])
    defparam FF_12.GSR = "ENABLED";
    FD1P3DX FF_11 (.D(s_Multiplier_0_2_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(736[13] 737[35])
    defparam FF_11.GSR = "ENABLED";
    FD1P3DX FF_10 (.D(s_Multiplier_0_2_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(740[13] 741[35])
    defparam FF_10.GSR = "ENABLED";
    FD1P3DX FF_9 (.D(s_Multiplier_0_2_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(744[13] 745[35])
    defparam FF_9.GSR = "ENABLED";
    FD1P3DX FF_8 (.D(s_Multiplier_0_2_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(748[13] 749[35])
    defparam FF_8.GSR = "ENABLED";
    FD1P3DX FF_7 (.D(s_Multiplier_0_2_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(752[13] 753[35])
    defparam FF_7.GSR = "ENABLED";
    FD1P3DX FF_6 (.D(s_Multiplier_0_2_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(756[13] 757[35])
    defparam FF_6.GSR = "ENABLED";
    FD1P3DX FF_5 (.D(s_Multiplier_0_2_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(760[13] 761[35])
    defparam FF_5.GSR = "ENABLED";
    FD1P3DX FF_4 (.D(s_Multiplier_0_2_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(764[13] 765[35])
    defparam FF_4.GSR = "ENABLED";
    FD1P3DX FF_3 (.D(s_Multiplier_0_2_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(768[13] 769[35])
    defparam FF_3.GSR = "ENABLED";
    FD1P3DX FF_2 (.D(s_Multiplier_0_2_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(772[13] 773[35])
    defparam FF_2.GSR = "ENABLED";
    FD1P3DX FF_1 (.D(s_Multiplier_0_2_22), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_22)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(776[13] 777[35])
    defparam FF_1.GSR = "ENABLED";
    FD1P3DX FF_0 (.D(s_Multiplier_0_2_23), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_23)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(780[13] 781[35])
    defparam FF_0.GSR = "ENABLED";
    FADD2B Multiplier_0_cin_lr_add_0 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_Cadd_0_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco), .S0(Multiplier_0_pp_0_13)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_cin_lr_add_2 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_Cadd_2_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_1), .S0(Multiplier_0_pp_1_15)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_cin_lr_add_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_Cadd_4_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_2), .S0(Multiplier_0_pp_2_17)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_cin_lr_add_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_Cadd_6_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_3), .S0(Multiplier_0_pp_3_19)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_cin_lr_add_8 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_Cadd_8_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_4), .S0(Multiplier_0_pp_4_21)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_cin_lr_add_10 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_Cadd_10_6 (.A0(VCC_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_5), .S0(Multiplier_0_pp_5_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_Multiplier_0_0_1 (.A0(GND_net), .A1(Multiplier_0_pp_0_2), 
           .B0(GND_net), .B1(Multiplier_0_pp_1_2), .CI(GND_net), .COUT(co_Multiplier_0_0_1), 
           .S1(s_Multiplier_0_0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_0_2 (.A0(Multiplier_0_pp_0_3), .A1(Multiplier_0_pp_0_4), 
           .B0(Multiplier_0_pp_1_3), .B1(Multiplier_0_pp_1_4), .CI(co_Multiplier_0_0_1), 
           .COUT(co_Multiplier_0_0_2), .S0(s_Multiplier_0_0_3), .S1(s_Multiplier_0_0_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_0_3 (.A0(Multiplier_0_pp_0_5), .A1(Multiplier_0_pp_0_6), 
           .B0(Multiplier_0_pp_1_5), .B1(Multiplier_0_pp_1_6), .CI(co_Multiplier_0_0_2), 
           .COUT(co_Multiplier_0_0_3), .S0(s_Multiplier_0_0_5), .S1(s_Multiplier_0_0_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_0_4 (.A0(Multiplier_0_pp_0_7), .A1(Multiplier_0_pp_0_8), 
           .B0(Multiplier_0_pp_1_7), .B1(Multiplier_0_pp_1_8), .CI(co_Multiplier_0_0_3), 
           .COUT(co_Multiplier_0_0_4), .S0(s_Multiplier_0_0_7), .S1(s_Multiplier_0_0_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_0_5 (.A0(Multiplier_0_pp_0_9), .A1(Multiplier_0_pp_0_10), 
           .B0(Multiplier_0_pp_1_9), .B1(Multiplier_0_pp_1_10), .CI(co_Multiplier_0_0_4), 
           .COUT(co_Multiplier_0_0_5), .S0(s_Multiplier_0_0_9), .S1(s_Multiplier_0_0_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_0_6 (.A0(Multiplier_0_pp_0_11), .A1(Multiplier_0_pp_0_12), 
           .B0(Multiplier_0_pp_1_11), .B1(Multiplier_0_pp_1_12), .CI(co_Multiplier_0_0_5), 
           .COUT(co_Multiplier_0_0_6), .S0(s_Multiplier_0_0_11), .S1(s_Multiplier_0_0_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_0_7 (.A0(Multiplier_0_pp_0_13), .A1(GND_net), 
           .B0(Multiplier_0_pp_1_13), .B1(Multiplier_0_pp_1_14), .CI(co_Multiplier_0_0_6), 
           .COUT(co_Multiplier_0_0_7), .S0(s_Multiplier_0_0_13), .S1(s_Multiplier_0_0_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_0_8 (.A0(GND_net), .A1(GND_net), .B0(Multiplier_0_pp_1_15), 
           .B1(GND_net), .CI(co_Multiplier_0_0_7), .COUT(co_Multiplier_0_0_8), 
           .S0(s_Multiplier_0_0_15), .S1(s_Multiplier_0_0_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_Multiplier_0_0_9 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_Multiplier_0_0_8), .S0(s_Multiplier_0_0_17)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_Multiplier_0_1_1 (.A0(GND_net), .A1(Multiplier_0_pp_2_6), 
           .B0(GND_net), .B1(Multiplier_0_pp_3_6), .CI(GND_net), .COUT(co_Multiplier_0_1_1), 
           .S1(s_Multiplier_0_1_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_1_2 (.A0(Multiplier_0_pp_2_7), .A1(Multiplier_0_pp_2_8), 
           .B0(Multiplier_0_pp_3_7), .B1(Multiplier_0_pp_3_8), .CI(co_Multiplier_0_1_1), 
           .COUT(co_Multiplier_0_1_2), .S0(s_Multiplier_0_1_7), .S1(s_Multiplier_0_1_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_1_3 (.A0(Multiplier_0_pp_2_9), .A1(Multiplier_0_pp_2_10), 
           .B0(Multiplier_0_pp_3_9), .B1(Multiplier_0_pp_3_10), .CI(co_Multiplier_0_1_2), 
           .COUT(co_Multiplier_0_1_3), .S0(s_Multiplier_0_1_9), .S1(s_Multiplier_0_1_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_1_4 (.A0(Multiplier_0_pp_2_11), .A1(Multiplier_0_pp_2_12), 
           .B0(Multiplier_0_pp_3_11), .B1(Multiplier_0_pp_3_12), .CI(co_Multiplier_0_1_3), 
           .COUT(co_Multiplier_0_1_4), .S0(s_Multiplier_0_1_11), .S1(s_Multiplier_0_1_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_1_5 (.A0(Multiplier_0_pp_2_13), .A1(Multiplier_0_pp_2_14), 
           .B0(Multiplier_0_pp_3_13), .B1(Multiplier_0_pp_3_14), .CI(co_Multiplier_0_1_4), 
           .COUT(co_Multiplier_0_1_5), .S0(s_Multiplier_0_1_13), .S1(s_Multiplier_0_1_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_1_6 (.A0(Multiplier_0_pp_2_15), .A1(Multiplier_0_pp_2_16), 
           .B0(Multiplier_0_pp_3_15), .B1(Multiplier_0_pp_3_16), .CI(co_Multiplier_0_1_5), 
           .COUT(co_Multiplier_0_1_6), .S0(s_Multiplier_0_1_15), .S1(s_Multiplier_0_1_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_1_7 (.A0(Multiplier_0_pp_2_17), .A1(GND_net), 
           .B0(Multiplier_0_pp_3_17), .B1(Multiplier_0_pp_3_18), .CI(co_Multiplier_0_1_6), 
           .COUT(co_Multiplier_0_1_7), .S0(s_Multiplier_0_1_17), .S1(s_Multiplier_0_1_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_1_8 (.A0(GND_net), .A1(GND_net), .B0(Multiplier_0_pp_3_19), 
           .B1(GND_net), .CI(co_Multiplier_0_1_7), .COUT(co_Multiplier_0_1_8), 
           .S0(s_Multiplier_0_1_19), .S1(s_Multiplier_0_1_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_Multiplier_0_1_9 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_Multiplier_0_1_8), .S0(s_Multiplier_0_1_21)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_Multiplier_0_2_1 (.A0(GND_net), .A1(Multiplier_0_pp_4_10), 
           .B0(GND_net), .B1(Multiplier_0_pp_5_10), .CI(GND_net), .COUT(co_Multiplier_0_2_1), 
           .S1(s_Multiplier_0_2_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_2_2 (.A0(Multiplier_0_pp_4_11), .A1(Multiplier_0_pp_4_12), 
           .B0(Multiplier_0_pp_5_11), .B1(Multiplier_0_pp_5_12), .CI(co_Multiplier_0_2_1), 
           .COUT(co_Multiplier_0_2_2), .S0(s_Multiplier_0_2_11), .S1(s_Multiplier_0_2_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_2_3 (.A0(Multiplier_0_pp_4_13), .A1(Multiplier_0_pp_4_14), 
           .B0(Multiplier_0_pp_5_13), .B1(Multiplier_0_pp_5_14), .CI(co_Multiplier_0_2_2), 
           .COUT(co_Multiplier_0_2_3), .S0(s_Multiplier_0_2_13), .S1(s_Multiplier_0_2_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_2_4 (.A0(Multiplier_0_pp_4_15), .A1(Multiplier_0_pp_4_16), 
           .B0(Multiplier_0_pp_5_15), .B1(Multiplier_0_pp_5_16), .CI(co_Multiplier_0_2_3), 
           .COUT(co_Multiplier_0_2_4), .S0(s_Multiplier_0_2_15), .S1(s_Multiplier_0_2_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_2_5 (.A0(Multiplier_0_pp_4_17), .A1(Multiplier_0_pp_4_18), 
           .B0(Multiplier_0_pp_5_17), .B1(Multiplier_0_pp_5_18), .CI(co_Multiplier_0_2_4), 
           .COUT(co_Multiplier_0_2_5), .S0(s_Multiplier_0_2_17), .S1(s_Multiplier_0_2_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_2_6 (.A0(Multiplier_0_pp_4_19), .A1(Multiplier_0_pp_4_20), 
           .B0(Multiplier_0_pp_5_19), .B1(Multiplier_0_pp_5_20), .CI(co_Multiplier_0_2_5), 
           .COUT(co_Multiplier_0_2_6), .S0(s_Multiplier_0_2_19), .S1(s_Multiplier_0_2_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_2_7 (.A0(Multiplier_0_pp_4_21), .A1(GND_net), 
           .B0(Multiplier_0_pp_5_21), .B1(Multiplier_0_pp_5_22), .CI(co_Multiplier_0_2_6), 
           .COUT(co_Multiplier_0_2_7), .S0(s_Multiplier_0_2_21), .S1(s_Multiplier_0_2_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_2_8 (.A0(GND_net), .A1(GND_net), .B0(Multiplier_0_pp_5_23), 
           .B1(GND_net), .CI(co_Multiplier_0_2_7), .S0(s_Multiplier_0_2_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_Multiplier_0_3_1 (.A0(GND_net), .A1(f_s_Multiplier_0_0_4), 
           .B0(GND_net), .B1(f_Multiplier_0_pp_2_4), .CI(GND_net), .COUT(co_Multiplier_0_3_1), 
           .S1(rego_o_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_2 (.A0(f_s_Multiplier_0_0_5), .A1(f_s_Multiplier_0_0_6), 
           .B0(f_Multiplier_0_pp_2_5), .B1(f_s_Multiplier_0_1_6), .CI(co_Multiplier_0_3_1), 
           .COUT(co_Multiplier_0_3_2), .S0(rego_o_5), .S1(rego_o_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_3 (.A0(f_s_Multiplier_0_0_7), .A1(f_s_Multiplier_0_0_8), 
           .B0(f_s_Multiplier_0_1_7), .B1(f_s_Multiplier_0_1_8), .CI(co_Multiplier_0_3_2), 
           .COUT(co_Multiplier_0_3_3), .S0(rego_o_7), .S1(s_Multiplier_0_3_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_4 (.A0(f_s_Multiplier_0_0_9), .A1(f_s_Multiplier_0_0_10), 
           .B0(f_s_Multiplier_0_1_9), .B1(f_s_Multiplier_0_1_10), .CI(co_Multiplier_0_3_3), 
           .COUT(co_Multiplier_0_3_4), .S0(s_Multiplier_0_3_9), .S1(s_Multiplier_0_3_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_5 (.A0(f_s_Multiplier_0_0_11), .A1(f_s_Multiplier_0_0_12), 
           .B0(f_s_Multiplier_0_1_11), .B1(f_s_Multiplier_0_1_12), .CI(co_Multiplier_0_3_4), 
           .COUT(co_Multiplier_0_3_5), .S0(s_Multiplier_0_3_11), .S1(s_Multiplier_0_3_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_6 (.A0(f_s_Multiplier_0_0_13), .A1(f_s_Multiplier_0_0_14), 
           .B0(f_s_Multiplier_0_1_13), .B1(f_s_Multiplier_0_1_14), .CI(co_Multiplier_0_3_5), 
           .COUT(co_Multiplier_0_3_6), .S0(s_Multiplier_0_3_13), .S1(s_Multiplier_0_3_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_7 (.A0(f_s_Multiplier_0_0_15), .A1(f_s_Multiplier_0_0_16), 
           .B0(f_s_Multiplier_0_1_15), .B1(f_s_Multiplier_0_1_16), .CI(co_Multiplier_0_3_6), 
           .COUT(co_Multiplier_0_3_7), .S0(s_Multiplier_0_3_15), .S1(s_Multiplier_0_3_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_8 (.A0(f_s_Multiplier_0_0_17), .A1(GND_net), 
           .B0(f_s_Multiplier_0_1_17), .B1(f_s_Multiplier_0_1_18), .CI(co_Multiplier_0_3_7), 
           .COUT(co_Multiplier_0_3_8), .S0(s_Multiplier_0_3_17), .S1(s_Multiplier_0_3_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_9 (.A0(GND_net), .A1(GND_net), .B0(f_s_Multiplier_0_1_19), 
           .B1(f_s_Multiplier_0_1_20), .CI(co_Multiplier_0_3_8), .COUT(co_Multiplier_0_3_9), 
           .S0(s_Multiplier_0_3_19), .S1(s_Multiplier_0_3_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_10 (.A0(GND_net), .A1(GND_net), .B0(f_s_Multiplier_0_1_21), 
           .B1(GND_net), .CI(co_Multiplier_0_3_9), .COUT(co_Multiplier_0_3_10), 
           .S0(s_Multiplier_0_3_21), .S1(s_Multiplier_0_3_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_Multiplier_0_3_11 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_Multiplier_0_3_10), .S0(s_Multiplier_0_3_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_t_Multiplier_0_4_1 (.A0(GND_net), .A1(s_Multiplier_0_3_8), 
           .B0(GND_net), .B1(f_Multiplier_0_pp_4_8), .CI(GND_net), .COUT(co_t_Multiplier_0_4_1), 
           .S1(rego_o_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_2 (.A0(s_Multiplier_0_3_9), .A1(s_Multiplier_0_3_10), 
           .B0(f_Multiplier_0_pp_4_9), .B1(f_s_Multiplier_0_2_10), .CI(co_t_Multiplier_0_4_1), 
           .COUT(co_t_Multiplier_0_4_2), .S0(rego_o_9), .S1(rego_o_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_3 (.A0(s_Multiplier_0_3_11), .A1(s_Multiplier_0_3_12), 
           .B0(f_s_Multiplier_0_2_11), .B1(f_s_Multiplier_0_2_12), .CI(co_t_Multiplier_0_4_2), 
           .COUT(co_t_Multiplier_0_4_3), .S0(rego_o_11), .S1(rego_o_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_4 (.A0(s_Multiplier_0_3_13), .A1(s_Multiplier_0_3_14), 
           .B0(f_s_Multiplier_0_2_13), .B1(f_s_Multiplier_0_2_14), .CI(co_t_Multiplier_0_4_3), 
           .COUT(co_t_Multiplier_0_4_4), .S0(rego_o_13), .S1(rego_o_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_5 (.A0(s_Multiplier_0_3_15), .A1(s_Multiplier_0_3_16), 
           .B0(f_s_Multiplier_0_2_15), .B1(f_s_Multiplier_0_2_16), .CI(co_t_Multiplier_0_4_4), 
           .COUT(co_t_Multiplier_0_4_5), .S0(rego_o_15), .S1(rego_o_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_6 (.A0(s_Multiplier_0_3_17), .A1(s_Multiplier_0_3_18), 
           .B0(f_s_Multiplier_0_2_17), .B1(f_s_Multiplier_0_2_18), .CI(co_t_Multiplier_0_4_5), 
           .COUT(co_t_Multiplier_0_4_6), .S0(rego_o_17), .S1(rego_o_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_7 (.A0(s_Multiplier_0_3_19), .A1(s_Multiplier_0_3_20), 
           .B0(f_s_Multiplier_0_2_19), .B1(f_s_Multiplier_0_2_20), .CI(co_t_Multiplier_0_4_6), 
           .COUT(co_t_Multiplier_0_4_7), .S0(rego_o_19), .S1(rego_o_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_8 (.A0(s_Multiplier_0_3_21), .A1(s_Multiplier_0_3_22), 
           .B0(f_s_Multiplier_0_2_21), .B1(f_s_Multiplier_0_2_22), .CI(co_t_Multiplier_0_4_7), 
           .COUT(co_t_Multiplier_0_4_8), .S0(rego_o_21), .S1(rego_o_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_9 (.A0(s_Multiplier_0_3_23), .A1(GND_net), 
           .B0(f_s_Multiplier_0_2_23), .B1(GND_net), .CI(co_t_Multiplier_0_4_8), 
           .S0(rego_o_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_0_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(Multiplier_0_cin_lr_0), .CO(mco), .P0(Multiplier_0_pp_0_1), 
          .P1(Multiplier_0_pp_0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_0_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco), .CO(mco_1), .P0(Multiplier_0_pp_0_3), 
          .P1(Multiplier_0_pp_0_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_0_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco_1), .CO(mco_2), .P0(Multiplier_0_pp_0_5), 
          .P1(Multiplier_0_pp_0_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_0_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco_2), .CO(mco_3), .P0(Multiplier_0_pp_0_7), 
          .P1(Multiplier_0_pp_0_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_0_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco_3), .CO(mco_4), .P0(Multiplier_0_pp_0_9), 
          .P1(Multiplier_0_pp_0_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_0_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_0_5_n2), 
          .A2(Multiplier_0_mult_0_5_n1), .A3(VCC_net), .B0(regb_b_1), 
          .B1(VCC_net), .B2(VCC_net), .B3(VCC_net), .CI(mco_4), .CO(mfco), 
          .P0(Multiplier_0_pp_0_11), .P1(Multiplier_0_pp_0_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_2_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(Multiplier_0_cin_lr_2), .CO(mco_5), .P0(Multiplier_0_pp_1_3), 
          .P1(Multiplier_0_pp_1_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_2_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_5), .CO(mco_6), .P0(Multiplier_0_pp_1_5), 
          .P1(Multiplier_0_pp_1_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_2_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_6), .CO(mco_7), .P0(Multiplier_0_pp_1_7), 
          .P1(Multiplier_0_pp_1_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_2_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_7), .CO(mco_8), .P0(Multiplier_0_pp_1_9), 
          .P1(Multiplier_0_pp_1_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_2_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_8), .CO(mco_9), .P0(Multiplier_0_pp_1_11), 
          .P1(Multiplier_0_pp_1_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_2_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_2_5_n2), 
          .A2(Multiplier_0_mult_2_5_n1), .A3(GND_net), .B0(regb_b_3), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_2), .CI(mco_9), .CO(mfco_1), 
          .P0(Multiplier_0_pp_1_13), .P1(Multiplier_0_pp_1_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_4_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(Multiplier_0_cin_lr_4), .CO(mco_10), .P0(Multiplier_0_pp_2_5), 
          .P1(Multiplier_0_pp_2_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_4_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_10), .CO(mco_11), .P0(Multiplier_0_pp_2_7), 
          .P1(Multiplier_0_pp_2_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_4_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_11), .CO(mco_12), .P0(Multiplier_0_pp_2_9), 
          .P1(Multiplier_0_pp_2_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_4_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_12), .CO(mco_13), .P0(Multiplier_0_pp_2_11), 
          .P1(Multiplier_0_pp_2_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_4_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_13), .CO(mco_14), .P0(Multiplier_0_pp_2_13), 
          .P1(Multiplier_0_pp_2_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_4_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_4_5_n2), 
          .A2(Multiplier_0_mult_4_5_n1), .A3(GND_net), .B0(regb_b_5), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_4), .CI(mco_14), .CO(mfco_2), 
          .P0(Multiplier_0_pp_2_15), .P1(Multiplier_0_pp_2_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_6_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(Multiplier_0_cin_lr_6), .CO(mco_15), .P0(Multiplier_0_pp_3_7), 
          .P1(Multiplier_0_pp_3_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_6_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_15), .CO(mco_16), .P0(Multiplier_0_pp_3_9), 
          .P1(Multiplier_0_pp_3_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_6_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_16), .CO(mco_17), .P0(Multiplier_0_pp_3_11), 
          .P1(Multiplier_0_pp_3_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_6_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_17), .CO(mco_18), .P0(Multiplier_0_pp_3_13), 
          .P1(Multiplier_0_pp_3_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_6_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_18), .CO(mco_19), .P0(Multiplier_0_pp_3_15), 
          .P1(Multiplier_0_pp_3_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_6_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_6_5_n2), 
          .A2(Multiplier_0_mult_6_5_n1), .A3(GND_net), .B0(regb_b_7), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_6), .CI(mco_19), .CO(mfco_3), 
          .P0(Multiplier_0_pp_3_17), .P1(Multiplier_0_pp_3_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_8_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(Multiplier_0_cin_lr_8), .CO(mco_20), .P0(Multiplier_0_pp_4_9), 
          .P1(Multiplier_0_pp_4_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_8_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_20), .CO(mco_21), .P0(Multiplier_0_pp_4_11), 
          .P1(Multiplier_0_pp_4_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_8_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_21), .CO(mco_22), .P0(Multiplier_0_pp_4_13), 
          .P1(Multiplier_0_pp_4_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_8_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_22), .CO(mco_23), .P0(Multiplier_0_pp_4_15), 
          .P1(Multiplier_0_pp_4_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_8_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_23), .CO(mco_24), .P0(Multiplier_0_pp_4_17), 
          .P1(Multiplier_0_pp_4_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_8_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_8_5_n2), 
          .A2(Multiplier_0_mult_8_5_n1), .A3(GND_net), .B0(regb_b_9), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_8), .CI(mco_24), .CO(mfco_4), 
          .P0(Multiplier_0_pp_4_19), .P1(Multiplier_0_pp_4_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_10_0 (.A0(Multiplier_0_mult_10_0_n0), .A1(rega_a_1), 
          .A2(Multiplier_0_mult_10_0_n1), .A3(rega_a_2), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(Multiplier_0_cin_lr_10), 
          .CO(mco_25), .P0(Multiplier_0_pp_5_11), .P1(Multiplier_0_pp_5_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_10_1 (.A0(Multiplier_0_mult_10_1_n0), .A1(rega_a_3), 
          .A2(Multiplier_0_mult_10_1_n1), .A3(rega_a_4), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_25), 
          .CO(mco_26), .P0(Multiplier_0_pp_5_13), .P1(Multiplier_0_pp_5_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_10_2 (.A0(Multiplier_0_mult_10_2_n0), .A1(rega_a_5), 
          .A2(Multiplier_0_mult_10_2_n1), .A3(rega_a_6), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_26), 
          .CO(mco_27), .P0(Multiplier_0_pp_5_15), .P1(Multiplier_0_pp_5_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_10_3 (.A0(Multiplier_0_mult_10_3_n0), .A1(rega_a_7), 
          .A2(Multiplier_0_mult_10_3_n1), .A3(rega_a_8), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_27), 
          .CO(mco_28), .P0(Multiplier_0_pp_5_17), .P1(Multiplier_0_pp_5_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_10_4 (.A0(Multiplier_0_mult_10_4_n0), .A1(rega_a_9), 
          .A2(Multiplier_0_mult_10_4_n1), .A3(rega_a_10), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_28), 
          .CO(mco_29), .P0(Multiplier_0_pp_5_19), .P1(Multiplier_0_pp_5_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_10_5 (.A0(Multiplier_0_mult_10_5_n0), .A1(Multiplier_0_mult_10_5_n2), 
          .A2(rega_a_11), .A3(GND_net), .B0(VCC_net), .B1(VCC_net), 
          .B2(regb_b_11), .B3(regb_b_10), .CI(mco_29), .CO(mfco_5), 
          .P0(Multiplier_0_pp_5_21), .P1(Multiplier_0_pp_5_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    AND2 AND2_t27 (.A(regb_b_0), .B(regb_b_0), .Z(Multiplier_0_pp_0_0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(376[10:72])
    ND2 ND2_t26 (.A(rega_a_11), .B(regb_b_0), .Z(Multiplier_0_mult_0_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t23 (.A(rega_a_11), .B(regb_b_2), .Z(Multiplier_0_mult_2_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t20 (.A(rega_a_11), .B(regb_b_4), .Z(Multiplier_0_mult_4_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t17 (.A(rega_a_11), .B(regb_b_6), .Z(Multiplier_0_mult_6_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t14 (.A(rega_a_11), .B(regb_b_8), .Z(Multiplier_0_mult_8_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t11 (.A(rega_a_1), .B(regb_b_11), .Z(Multiplier_0_mult_10_0_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    
endmodule
//
// Verilog Description of module Multiplier_U0
//

module Multiplier_U0 (CIC1_out_clkSin, VCC_net, GND_net, MultDataB, 
            MultResult1) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input CIC1_out_clkSin;
    input VCC_net;
    input GND_net;
    input [11:0]MultDataB;
    output [23:0]MultResult1;
    
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(85[6:21])
    
    wire Multiplier_0_mult_0_5_n1, regb_b_1, rega_a_11, Multiplier_0_pp_1_2, 
        regb_b_2, regb_b_0, Multiplier_0_mult_2_5_n1, regb_b_3, Multiplier_0_pp_2_4, 
        regb_b_4, Multiplier_0_mult_4_5_n1, regb_b_5, Multiplier_0_pp_3_6, 
        regb_b_6, Multiplier_0_mult_6_5_n1, regb_b_7, Multiplier_0_pp_4_8, 
        regb_b_8, Multiplier_0_mult_8_5_n1, regb_b_9, Multiplier_0_pp_5_10, 
        regb_b_10, Multiplier_0_mult_10_0_n0, regb_b_11, Multiplier_0_mult_10_1_n1, 
        rega_a_3, rega_a_2, Multiplier_0_mult_10_1_n0, Multiplier_0_mult_10_2_n1, 
        rega_a_5, rega_a_4, Multiplier_0_mult_10_2_n0, Multiplier_0_mult_10_3_n1, 
        rega_a_7, rega_a_6, Multiplier_0_mult_10_3_n0, Multiplier_0_mult_10_4_n1, 
        rega_a_9, rega_a_8, Multiplier_0_mult_10_4_n0, Multiplier_0_mult_10_5_n2, 
        rega_a_10, Multiplier_0_mult_10_5_n0, rega_a_1, rego_o_0, rego_o_1, 
        rego_o_2, rego_o_3, rego_o_4, rego_o_5, rego_o_6, rego_o_7, 
        rego_o_8, rego_o_9, rego_o_10, rego_o_11, rego_o_12, rego_o_13, 
        rego_o_14, rego_o_15, rego_o_16, rego_o_17, rego_o_18, rego_o_19, 
        rego_o_20, rego_o_21, rego_o_22, rego_o_23, Multiplier_0_pp_0_0, 
        Multiplier_0_pp_0_1, s_Multiplier_0_0_2, s_Multiplier_0_0_3, s_Multiplier_0_0_4, 
        f_s_Multiplier_0_0_4, s_Multiplier_0_0_5, f_s_Multiplier_0_0_5, 
        s_Multiplier_0_0_6, f_s_Multiplier_0_0_6, s_Multiplier_0_0_7, 
        f_s_Multiplier_0_0_7, s_Multiplier_0_0_8, f_s_Multiplier_0_0_8, 
        s_Multiplier_0_0_9, f_s_Multiplier_0_0_9, s_Multiplier_0_0_10, 
        f_s_Multiplier_0_0_10, s_Multiplier_0_0_11, f_s_Multiplier_0_0_11, 
        s_Multiplier_0_0_12, f_s_Multiplier_0_0_12, s_Multiplier_0_0_13, 
        f_s_Multiplier_0_0_13, s_Multiplier_0_0_14, f_s_Multiplier_0_0_14, 
        s_Multiplier_0_0_15, f_s_Multiplier_0_0_15, s_Multiplier_0_0_16, 
        f_s_Multiplier_0_0_16, s_Multiplier_0_0_17, f_s_Multiplier_0_0_17, 
        f_Multiplier_0_pp_2_4, f_Multiplier_0_pp_2_5, Multiplier_0_pp_2_5, 
        s_Multiplier_0_1_6, f_s_Multiplier_0_1_6, s_Multiplier_0_1_7, 
        f_s_Multiplier_0_1_7, s_Multiplier_0_1_8, f_s_Multiplier_0_1_8, 
        s_Multiplier_0_1_9, f_s_Multiplier_0_1_9, s_Multiplier_0_1_10, 
        f_s_Multiplier_0_1_10, s_Multiplier_0_1_11, f_s_Multiplier_0_1_11, 
        s_Multiplier_0_1_12, f_s_Multiplier_0_1_12, s_Multiplier_0_1_13, 
        f_s_Multiplier_0_1_13, s_Multiplier_0_1_14, f_s_Multiplier_0_1_14, 
        s_Multiplier_0_1_15, f_s_Multiplier_0_1_15, s_Multiplier_0_1_16, 
        f_s_Multiplier_0_1_16, s_Multiplier_0_1_17, f_s_Multiplier_0_1_17, 
        s_Multiplier_0_1_18, f_s_Multiplier_0_1_18, s_Multiplier_0_1_19, 
        f_s_Multiplier_0_1_19, s_Multiplier_0_1_20, f_s_Multiplier_0_1_20, 
        s_Multiplier_0_1_21, f_s_Multiplier_0_1_21, f_Multiplier_0_pp_4_8, 
        f_Multiplier_0_pp_4_9, Multiplier_0_pp_4_9, s_Multiplier_0_2_10, 
        f_s_Multiplier_0_2_10, s_Multiplier_0_2_11, f_s_Multiplier_0_2_11, 
        s_Multiplier_0_2_12, f_s_Multiplier_0_2_12, s_Multiplier_0_2_13, 
        f_s_Multiplier_0_2_13, s_Multiplier_0_2_14, f_s_Multiplier_0_2_14, 
        s_Multiplier_0_2_15, f_s_Multiplier_0_2_15, s_Multiplier_0_2_16, 
        f_s_Multiplier_0_2_16, s_Multiplier_0_2_17, f_s_Multiplier_0_2_17, 
        s_Multiplier_0_2_18, f_s_Multiplier_0_2_18, s_Multiplier_0_2_19, 
        f_s_Multiplier_0_2_19, s_Multiplier_0_2_20, f_s_Multiplier_0_2_20, 
        s_Multiplier_0_2_21, f_s_Multiplier_0_2_21, s_Multiplier_0_2_22, 
        f_s_Multiplier_0_2_22, s_Multiplier_0_2_23, f_s_Multiplier_0_2_23, 
        Multiplier_0_cin_lr_0, Multiplier_0_pp_0_13, mfco, Multiplier_0_cin_lr_2, 
        Multiplier_0_pp_1_15, mfco_1, Multiplier_0_cin_lr_4, Multiplier_0_pp_2_17, 
        mfco_2, Multiplier_0_cin_lr_6, Multiplier_0_pp_3_19, mfco_3, 
        Multiplier_0_cin_lr_8, Multiplier_0_pp_4_21, mfco_4, Multiplier_0_cin_lr_10, 
        Multiplier_0_pp_5_23, mfco_5, co_Multiplier_0_0_1, Multiplier_0_pp_0_2, 
        co_Multiplier_0_0_2, Multiplier_0_pp_0_4, Multiplier_0_pp_0_3, 
        Multiplier_0_pp_1_4, Multiplier_0_pp_1_3, co_Multiplier_0_0_3, 
        Multiplier_0_pp_0_6, Multiplier_0_pp_0_5, Multiplier_0_pp_1_6, 
        Multiplier_0_pp_1_5, co_Multiplier_0_0_4, Multiplier_0_pp_0_8, 
        Multiplier_0_pp_0_7, Multiplier_0_pp_1_8, Multiplier_0_pp_1_7, 
        co_Multiplier_0_0_5, Multiplier_0_pp_0_10, Multiplier_0_pp_0_9, 
        Multiplier_0_pp_1_10, Multiplier_0_pp_1_9, co_Multiplier_0_0_6, 
        Multiplier_0_pp_0_12, Multiplier_0_pp_0_11, Multiplier_0_pp_1_12, 
        Multiplier_0_pp_1_11, co_Multiplier_0_0_7, Multiplier_0_pp_1_14, 
        Multiplier_0_pp_1_13, co_Multiplier_0_0_8, co_Multiplier_0_1_1, 
        Multiplier_0_pp_2_6, co_Multiplier_0_1_2, Multiplier_0_pp_2_8, 
        Multiplier_0_pp_2_7, Multiplier_0_pp_3_8, Multiplier_0_pp_3_7, 
        co_Multiplier_0_1_3, Multiplier_0_pp_2_10, Multiplier_0_pp_2_9, 
        Multiplier_0_pp_3_10, Multiplier_0_pp_3_9, co_Multiplier_0_1_4, 
        Multiplier_0_pp_2_12, Multiplier_0_pp_2_11, Multiplier_0_pp_3_12, 
        Multiplier_0_pp_3_11, co_Multiplier_0_1_5, Multiplier_0_pp_2_14, 
        Multiplier_0_pp_2_13, Multiplier_0_pp_3_14, Multiplier_0_pp_3_13, 
        co_Multiplier_0_1_6, Multiplier_0_pp_2_16, Multiplier_0_pp_2_15, 
        Multiplier_0_pp_3_16, Multiplier_0_pp_3_15, co_Multiplier_0_1_7, 
        Multiplier_0_pp_3_18, Multiplier_0_pp_3_17, co_Multiplier_0_1_8, 
        co_Multiplier_0_2_1, Multiplier_0_pp_4_10, co_Multiplier_0_2_2, 
        Multiplier_0_pp_4_12, Multiplier_0_pp_4_11, Multiplier_0_pp_5_12, 
        Multiplier_0_pp_5_11, co_Multiplier_0_2_3, Multiplier_0_pp_4_14, 
        Multiplier_0_pp_4_13, Multiplier_0_pp_5_14, Multiplier_0_pp_5_13, 
        co_Multiplier_0_2_4, Multiplier_0_pp_4_16, Multiplier_0_pp_4_15, 
        Multiplier_0_pp_5_16, Multiplier_0_pp_5_15, co_Multiplier_0_2_5, 
        Multiplier_0_pp_4_18, Multiplier_0_pp_4_17, Multiplier_0_pp_5_18, 
        Multiplier_0_pp_5_17, co_Multiplier_0_2_6, Multiplier_0_pp_4_20, 
        Multiplier_0_pp_4_19, Multiplier_0_pp_5_20, Multiplier_0_pp_5_19, 
        co_Multiplier_0_2_7, Multiplier_0_pp_5_22, Multiplier_0_pp_5_21, 
        co_Multiplier_0_3_1, co_Multiplier_0_3_2, co_Multiplier_0_3_3, 
        s_Multiplier_0_3_8, co_Multiplier_0_3_4, s_Multiplier_0_3_9, s_Multiplier_0_3_10, 
        co_Multiplier_0_3_5, s_Multiplier_0_3_11, s_Multiplier_0_3_12, 
        co_Multiplier_0_3_6, s_Multiplier_0_3_13, s_Multiplier_0_3_14, 
        co_Multiplier_0_3_7, s_Multiplier_0_3_15, s_Multiplier_0_3_16, 
        co_Multiplier_0_3_8, s_Multiplier_0_3_17, s_Multiplier_0_3_18, 
        co_Multiplier_0_3_9, s_Multiplier_0_3_19, s_Multiplier_0_3_20, 
        co_Multiplier_0_3_10, s_Multiplier_0_3_21, s_Multiplier_0_3_22, 
        s_Multiplier_0_3_23, co_t_Multiplier_0_4_1, co_t_Multiplier_0_4_2, 
        co_t_Multiplier_0_4_3, co_t_Multiplier_0_4_4, co_t_Multiplier_0_4_5, 
        co_t_Multiplier_0_4_6, co_t_Multiplier_0_4_7, co_t_Multiplier_0_4_8, 
        mco, mco_1, mco_2, mco_3, mco_4, Multiplier_0_mult_0_5_n2, 
        mco_5, mco_6, mco_7, mco_8, mco_9, Multiplier_0_mult_2_5_n2, 
        mco_10, mco_11, mco_12, mco_13, mco_14, Multiplier_0_mult_4_5_n2, 
        mco_15, mco_16, mco_17, mco_18, mco_19, Multiplier_0_mult_6_5_n2, 
        mco_20, mco_21, mco_22, mco_23, mco_24, Multiplier_0_mult_8_5_n2, 
        Multiplier_0_mult_10_0_n1, mco_25, mco_26, mco_27, mco_28, 
        mco_29;
    
    ND2 ND2_t25 (.A(rega_a_11), .B(regb_b_1), .Z(Multiplier_0_mult_0_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    AND2 AND2_t24 (.A(regb_b_0), .B(regb_b_2), .Z(Multiplier_0_pp_1_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(382[10:72])
    ND2 ND2_t22 (.A(rega_a_11), .B(regb_b_3), .Z(Multiplier_0_mult_2_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    AND2 AND2_t21 (.A(regb_b_0), .B(regb_b_4), .Z(Multiplier_0_pp_2_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(388[10:72])
    ND2 ND2_t19 (.A(rega_a_11), .B(regb_b_5), .Z(Multiplier_0_mult_4_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    AND2 AND2_t18 (.A(regb_b_0), .B(regb_b_6), .Z(Multiplier_0_pp_3_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(394[10:72])
    ND2 ND2_t16 (.A(rega_a_11), .B(regb_b_7), .Z(Multiplier_0_mult_6_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    AND2 AND2_t15 (.A(regb_b_0), .B(regb_b_8), .Z(Multiplier_0_pp_4_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(400[10:72])
    ND2 ND2_t13 (.A(rega_a_11), .B(regb_b_9), .Z(Multiplier_0_mult_8_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    AND2 AND2_t12 (.A(regb_b_0), .B(regb_b_10), .Z(Multiplier_0_pp_5_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(406[10:74])
    ND2 ND2_t10 (.A(regb_b_0), .B(regb_b_11), .Z(Multiplier_0_mult_10_0_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t9 (.A(rega_a_3), .B(regb_b_11), .Z(Multiplier_0_mult_10_1_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t8 (.A(rega_a_2), .B(regb_b_11), .Z(Multiplier_0_mult_10_1_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t7 (.A(rega_a_5), .B(regb_b_11), .Z(Multiplier_0_mult_10_2_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t6 (.A(rega_a_4), .B(regb_b_11), .Z(Multiplier_0_mult_10_2_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t5 (.A(rega_a_7), .B(regb_b_11), .Z(Multiplier_0_mult_10_3_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t4 (.A(rega_a_6), .B(regb_b_11), .Z(Multiplier_0_mult_10_3_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t3 (.A(rega_a_9), .B(regb_b_11), .Z(Multiplier_0_mult_10_4_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t2 (.A(rega_a_8), .B(regb_b_11), .Z(Multiplier_0_mult_10_4_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t1 (.A(rega_a_11), .B(regb_b_10), .Z(Multiplier_0_mult_10_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t0 (.A(rega_a_10), .B(regb_b_11), .Z(Multiplier_0_mult_10_5_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FD1P3DX FF_98 (.D(MultDataB[1]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(435[13:82])
    defparam FF_98.GSR = "ENABLED";
    FD1P3DX FF_97 (.D(MultDataB[2]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(438[13:82])
    defparam FF_97.GSR = "ENABLED";
    FD1P3DX FF_96 (.D(MultDataB[3]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(441[13:82])
    defparam FF_96.GSR = "ENABLED";
    FD1P3DX FF_95 (.D(MultDataB[4]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(444[13:82])
    defparam FF_95.GSR = "ENABLED";
    FD1P3DX FF_94 (.D(MultDataB[5]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(447[13:82])
    defparam FF_94.GSR = "ENABLED";
    FD1P3DX FF_93 (.D(MultDataB[6]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(450[13:82])
    defparam FF_93.GSR = "ENABLED";
    FD1P3DX FF_92 (.D(MultDataB[7]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(453[13:82])
    defparam FF_92.GSR = "ENABLED";
    FD1P3DX FF_91 (.D(MultDataB[8]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(456[13:82])
    defparam FF_91.GSR = "ENABLED";
    FD1P3DX FF_90 (.D(MultDataB[9]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(459[13:82])
    defparam FF_90.GSR = "ENABLED";
    FD1P3DX FF_89 (.D(MultDataB[10]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(462[13:84])
    defparam FF_89.GSR = "ENABLED";
    FD1P3DX FF_88 (.D(MultDataB[11]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(465[13:84])
    defparam FF_88.GSR = "ENABLED";
    FD1P3DX FF_87 (.D(MultDataB[0]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_0)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(468[13:82])
    defparam FF_87.GSR = "ENABLED";
    FD1P3DX FF_86 (.D(MultDataB[1]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(471[13:82])
    defparam FF_86.GSR = "ENABLED";
    FD1P3DX FF_85 (.D(MultDataB[2]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(474[13:82])
    defparam FF_85.GSR = "ENABLED";
    FD1P3DX FF_84 (.D(MultDataB[3]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(477[13:82])
    defparam FF_84.GSR = "ENABLED";
    FD1P3DX FF_83 (.D(MultDataB[4]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(480[13:82])
    defparam FF_83.GSR = "ENABLED";
    FD1P3DX FF_82 (.D(MultDataB[5]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(483[13:82])
    defparam FF_82.GSR = "ENABLED";
    FD1P3DX FF_81 (.D(MultDataB[6]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(486[13:82])
    defparam FF_81.GSR = "ENABLED";
    FD1P3DX FF_80 (.D(MultDataB[7]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(489[13:82])
    defparam FF_80.GSR = "ENABLED";
    FD1P3DX FF_79 (.D(MultDataB[8]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(492[13:82])
    defparam FF_79.GSR = "ENABLED";
    FD1P3DX FF_78 (.D(MultDataB[9]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(495[13:82])
    defparam FF_78.GSR = "ENABLED";
    FD1P3DX FF_77 (.D(MultDataB[10]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(498[13:84])
    defparam FF_77.GSR = "ENABLED";
    FD1P3DX FF_76 (.D(MultDataB[11]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(501[13:84])
    defparam FF_76.GSR = "ENABLED";
    FD1P3DX FF_75 (.D(rego_o_0), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[0])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(504[13:83])
    defparam FF_75.GSR = "ENABLED";
    FD1P3DX FF_74 (.D(rego_o_1), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[1])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(507[13:83])
    defparam FF_74.GSR = "ENABLED";
    FD1P3DX FF_73 (.D(rego_o_2), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[2])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(510[13:83])
    defparam FF_73.GSR = "ENABLED";
    FD1P3DX FF_72 (.D(rego_o_3), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[3])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(513[13:83])
    defparam FF_72.GSR = "ENABLED";
    FD1P3DX FF_71 (.D(rego_o_4), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[4])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(516[13:83])
    defparam FF_71.GSR = "ENABLED";
    FD1P3DX FF_70 (.D(rego_o_5), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[5])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(519[13:83])
    defparam FF_70.GSR = "ENABLED";
    FD1P3DX FF_69 (.D(rego_o_6), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[6])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(522[13:83])
    defparam FF_69.GSR = "ENABLED";
    FD1P3DX FF_68 (.D(rego_o_7), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[7])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(525[13:83])
    defparam FF_68.GSR = "ENABLED";
    FD1P3DX FF_67 (.D(rego_o_8), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[8])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(528[13:83])
    defparam FF_67.GSR = "ENABLED";
    FD1P3DX FF_66 (.D(rego_o_9), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[9])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(531[13:83])
    defparam FF_66.GSR = "ENABLED";
    FD1P3DX FF_65 (.D(rego_o_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[10])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(534[13:85])
    defparam FF_65.GSR = "ENABLED";
    FD1P3DX FF_64 (.D(rego_o_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[11])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(537[13:85])
    defparam FF_64.GSR = "ENABLED";
    FD1P3DX FF_63 (.D(rego_o_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[12])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(540[13:85])
    defparam FF_63.GSR = "ENABLED";
    FD1P3DX FF_62 (.D(rego_o_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[13])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(543[13:85])
    defparam FF_62.GSR = "ENABLED";
    FD1P3DX FF_61 (.D(rego_o_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[14])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(546[13:85])
    defparam FF_61.GSR = "ENABLED";
    FD1P3DX FF_60 (.D(rego_o_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[15])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(549[13:85])
    defparam FF_60.GSR = "ENABLED";
    FD1P3DX FF_59 (.D(rego_o_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[16])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(552[13:85])
    defparam FF_59.GSR = "ENABLED";
    FD1P3DX FF_58 (.D(rego_o_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[17])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(555[13:85])
    defparam FF_58.GSR = "ENABLED";
    FD1P3DX FF_57 (.D(rego_o_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[18])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(558[13:85])
    defparam FF_57.GSR = "ENABLED";
    FD1P3DX FF_56 (.D(rego_o_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[19])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(561[13:85])
    defparam FF_56.GSR = "ENABLED";
    FD1P3DX FF_55 (.D(rego_o_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[20])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(564[13:85])
    defparam FF_55.GSR = "ENABLED";
    FD1P3DX FF_54 (.D(rego_o_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[21])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(567[13:85])
    defparam FF_54.GSR = "ENABLED";
    FD1P3DX FF_53 (.D(rego_o_22), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[22])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(570[13:85])
    defparam FF_53.GSR = "ENABLED";
    FD1P3DX FF_52 (.D(rego_o_23), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[23])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(573[13:85])
    defparam FF_52.GSR = "ENABLED";
    FD1P3DX FF_51 (.D(Multiplier_0_pp_0_0), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_0)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(576[13] 577[35])
    defparam FF_51.GSR = "ENABLED";
    FD1P3DX FF_50 (.D(Multiplier_0_pp_0_1), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(580[13] 581[35])
    defparam FF_50.GSR = "ENABLED";
    FD1P3DX FF_49 (.D(s_Multiplier_0_0_2), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(584[13] 585[34])
    defparam FF_49.GSR = "ENABLED";
    FD1P3DX FF_48 (.D(s_Multiplier_0_0_3), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(588[13] 589[34])
    defparam FF_48.GSR = "ENABLED";
    FD1P3DX FF_47 (.D(s_Multiplier_0_0_4), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(592[13] 593[34])
    defparam FF_47.GSR = "ENABLED";
    FD1P3DX FF_46 (.D(s_Multiplier_0_0_5), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(596[13] 597[34])
    defparam FF_46.GSR = "ENABLED";
    FD1P3DX FF_45 (.D(s_Multiplier_0_0_6), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(600[13] 601[34])
    defparam FF_45.GSR = "ENABLED";
    FD1P3DX FF_44 (.D(s_Multiplier_0_0_7), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(604[13] 605[34])
    defparam FF_44.GSR = "ENABLED";
    FD1P3DX FF_43 (.D(s_Multiplier_0_0_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(608[13] 609[34])
    defparam FF_43.GSR = "ENABLED";
    FD1P3DX FF_42 (.D(s_Multiplier_0_0_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(612[13] 613[34])
    defparam FF_42.GSR = "ENABLED";
    FD1P3DX FF_41 (.D(s_Multiplier_0_0_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(616[13] 617[35])
    defparam FF_41.GSR = "ENABLED";
    FD1P3DX FF_40 (.D(s_Multiplier_0_0_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(620[13] 621[35])
    defparam FF_40.GSR = "ENABLED";
    FD1P3DX FF_39 (.D(s_Multiplier_0_0_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(624[13] 625[35])
    defparam FF_39.GSR = "ENABLED";
    FD1P3DX FF_38 (.D(s_Multiplier_0_0_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(628[13] 629[35])
    defparam FF_38.GSR = "ENABLED";
    FD1P3DX FF_37 (.D(s_Multiplier_0_0_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(632[13] 633[35])
    defparam FF_37.GSR = "ENABLED";
    FD1P3DX FF_36 (.D(s_Multiplier_0_0_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(636[13] 637[35])
    defparam FF_36.GSR = "ENABLED";
    FD1P3DX FF_35 (.D(s_Multiplier_0_0_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(640[13] 641[35])
    defparam FF_35.GSR = "ENABLED";
    FD1P3DX FF_34 (.D(s_Multiplier_0_0_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(644[13] 645[35])
    defparam FF_34.GSR = "ENABLED";
    FD1P3DX FF_33 (.D(Multiplier_0_pp_2_4), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_2_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(648[13] 649[35])
    defparam FF_33.GSR = "ENABLED";
    FD1P3DX FF_32 (.D(Multiplier_0_pp_2_5), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_2_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(652[13] 653[35])
    defparam FF_32.GSR = "ENABLED";
    FD1P3DX FF_31 (.D(s_Multiplier_0_1_6), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(656[13] 657[34])
    defparam FF_31.GSR = "ENABLED";
    FD1P3DX FF_30 (.D(s_Multiplier_0_1_7), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(660[13] 661[34])
    defparam FF_30.GSR = "ENABLED";
    FD1P3DX FF_29 (.D(s_Multiplier_0_1_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(664[13] 665[34])
    defparam FF_29.GSR = "ENABLED";
    FD1P3DX FF_28 (.D(s_Multiplier_0_1_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(668[13] 669[34])
    defparam FF_28.GSR = "ENABLED";
    FD1P3DX FF_27 (.D(s_Multiplier_0_1_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(672[13] 673[35])
    defparam FF_27.GSR = "ENABLED";
    FD1P3DX FF_26 (.D(s_Multiplier_0_1_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(676[13] 677[35])
    defparam FF_26.GSR = "ENABLED";
    FD1P3DX FF_25 (.D(s_Multiplier_0_1_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(680[13] 681[35])
    defparam FF_25.GSR = "ENABLED";
    FD1P3DX FF_24 (.D(s_Multiplier_0_1_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(684[13] 685[35])
    defparam FF_24.GSR = "ENABLED";
    FD1P3DX FF_23 (.D(s_Multiplier_0_1_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(688[13] 689[35])
    defparam FF_23.GSR = "ENABLED";
    FD1P3DX FF_22 (.D(s_Multiplier_0_1_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(692[13] 693[35])
    defparam FF_22.GSR = "ENABLED";
    FD1P3DX FF_21 (.D(s_Multiplier_0_1_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(696[13] 697[35])
    defparam FF_21.GSR = "ENABLED";
    FD1P3DX FF_20 (.D(s_Multiplier_0_1_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(700[13] 701[35])
    defparam FF_20.GSR = "ENABLED";
    FD1P3DX FF_19 (.D(s_Multiplier_0_1_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(704[13] 705[35])
    defparam FF_19.GSR = "ENABLED";
    FD1P3DX FF_18 (.D(s_Multiplier_0_1_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(708[13] 709[35])
    defparam FF_18.GSR = "ENABLED";
    FD1P3DX FF_17 (.D(s_Multiplier_0_1_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(712[13] 713[35])
    defparam FF_17.GSR = "ENABLED";
    FD1P3DX FF_16 (.D(s_Multiplier_0_1_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(716[13] 717[35])
    defparam FF_16.GSR = "ENABLED";
    FD1P3DX FF_15 (.D(Multiplier_0_pp_4_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_4_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(720[13] 721[35])
    defparam FF_15.GSR = "ENABLED";
    FD1P3DX FF_14 (.D(Multiplier_0_pp_4_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_4_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(724[13] 725[35])
    defparam FF_14.GSR = "ENABLED";
    FD1P3DX FF_13 (.D(s_Multiplier_0_2_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(728[13] 729[35])
    defparam FF_13.GSR = "ENABLED";
    FD1P3DX FF_12 (.D(s_Multiplier_0_2_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(732[13] 733[35])
    defparam FF_12.GSR = "ENABLED";
    FD1P3DX FF_11 (.D(s_Multiplier_0_2_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(736[13] 737[35])
    defparam FF_11.GSR = "ENABLED";
    FD1P3DX FF_10 (.D(s_Multiplier_0_2_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(740[13] 741[35])
    defparam FF_10.GSR = "ENABLED";
    FD1P3DX FF_9 (.D(s_Multiplier_0_2_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(744[13] 745[35])
    defparam FF_9.GSR = "ENABLED";
    FD1P3DX FF_8 (.D(s_Multiplier_0_2_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(748[13] 749[35])
    defparam FF_8.GSR = "ENABLED";
    FD1P3DX FF_7 (.D(s_Multiplier_0_2_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(752[13] 753[35])
    defparam FF_7.GSR = "ENABLED";
    FD1P3DX FF_6 (.D(s_Multiplier_0_2_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(756[13] 757[35])
    defparam FF_6.GSR = "ENABLED";
    FD1P3DX FF_5 (.D(s_Multiplier_0_2_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(760[13] 761[35])
    defparam FF_5.GSR = "ENABLED";
    FD1P3DX FF_4 (.D(s_Multiplier_0_2_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(764[13] 765[35])
    defparam FF_4.GSR = "ENABLED";
    FD1P3DX FF_3 (.D(s_Multiplier_0_2_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(768[13] 769[35])
    defparam FF_3.GSR = "ENABLED";
    FD1P3DX FF_2 (.D(s_Multiplier_0_2_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(772[13] 773[35])
    defparam FF_2.GSR = "ENABLED";
    FD1P3DX FF_1 (.D(s_Multiplier_0_2_22), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_22)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(776[13] 777[35])
    defparam FF_1.GSR = "ENABLED";
    FD1P3DX FF_0 (.D(s_Multiplier_0_2_23), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_23)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(780[13] 781[35])
    defparam FF_0.GSR = "ENABLED";
    FADD2B Multiplier_0_cin_lr_add_0 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_Cadd_0_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco), .S0(Multiplier_0_pp_0_13)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_cin_lr_add_2 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_Cadd_2_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_1), .S0(Multiplier_0_pp_1_15)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_cin_lr_add_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_Cadd_4_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_2), .S0(Multiplier_0_pp_2_17)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_cin_lr_add_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_Cadd_6_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_3), .S0(Multiplier_0_pp_3_19)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_cin_lr_add_8 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_Cadd_8_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_4), .S0(Multiplier_0_pp_4_21)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_cin_lr_add_10 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_Cadd_10_6 (.A0(VCC_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_5), .S0(Multiplier_0_pp_5_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_Multiplier_0_0_1 (.A0(GND_net), .A1(Multiplier_0_pp_0_2), 
           .B0(GND_net), .B1(Multiplier_0_pp_1_2), .CI(GND_net), .COUT(co_Multiplier_0_0_1), 
           .S1(s_Multiplier_0_0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_0_2 (.A0(Multiplier_0_pp_0_3), .A1(Multiplier_0_pp_0_4), 
           .B0(Multiplier_0_pp_1_3), .B1(Multiplier_0_pp_1_4), .CI(co_Multiplier_0_0_1), 
           .COUT(co_Multiplier_0_0_2), .S0(s_Multiplier_0_0_3), .S1(s_Multiplier_0_0_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_0_3 (.A0(Multiplier_0_pp_0_5), .A1(Multiplier_0_pp_0_6), 
           .B0(Multiplier_0_pp_1_5), .B1(Multiplier_0_pp_1_6), .CI(co_Multiplier_0_0_2), 
           .COUT(co_Multiplier_0_0_3), .S0(s_Multiplier_0_0_5), .S1(s_Multiplier_0_0_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_0_4 (.A0(Multiplier_0_pp_0_7), .A1(Multiplier_0_pp_0_8), 
           .B0(Multiplier_0_pp_1_7), .B1(Multiplier_0_pp_1_8), .CI(co_Multiplier_0_0_3), 
           .COUT(co_Multiplier_0_0_4), .S0(s_Multiplier_0_0_7), .S1(s_Multiplier_0_0_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_0_5 (.A0(Multiplier_0_pp_0_9), .A1(Multiplier_0_pp_0_10), 
           .B0(Multiplier_0_pp_1_9), .B1(Multiplier_0_pp_1_10), .CI(co_Multiplier_0_0_4), 
           .COUT(co_Multiplier_0_0_5), .S0(s_Multiplier_0_0_9), .S1(s_Multiplier_0_0_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_0_6 (.A0(Multiplier_0_pp_0_11), .A1(Multiplier_0_pp_0_12), 
           .B0(Multiplier_0_pp_1_11), .B1(Multiplier_0_pp_1_12), .CI(co_Multiplier_0_0_5), 
           .COUT(co_Multiplier_0_0_6), .S0(s_Multiplier_0_0_11), .S1(s_Multiplier_0_0_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_0_7 (.A0(Multiplier_0_pp_0_13), .A1(GND_net), 
           .B0(Multiplier_0_pp_1_13), .B1(Multiplier_0_pp_1_14), .CI(co_Multiplier_0_0_6), 
           .COUT(co_Multiplier_0_0_7), .S0(s_Multiplier_0_0_13), .S1(s_Multiplier_0_0_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_0_8 (.A0(GND_net), .A1(GND_net), .B0(Multiplier_0_pp_1_15), 
           .B1(GND_net), .CI(co_Multiplier_0_0_7), .COUT(co_Multiplier_0_0_8), 
           .S0(s_Multiplier_0_0_15), .S1(s_Multiplier_0_0_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_Multiplier_0_0_9 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_Multiplier_0_0_8), .S0(s_Multiplier_0_0_17)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_Multiplier_0_1_1 (.A0(GND_net), .A1(Multiplier_0_pp_2_6), 
           .B0(GND_net), .B1(Multiplier_0_pp_3_6), .CI(GND_net), .COUT(co_Multiplier_0_1_1), 
           .S1(s_Multiplier_0_1_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_1_2 (.A0(Multiplier_0_pp_2_7), .A1(Multiplier_0_pp_2_8), 
           .B0(Multiplier_0_pp_3_7), .B1(Multiplier_0_pp_3_8), .CI(co_Multiplier_0_1_1), 
           .COUT(co_Multiplier_0_1_2), .S0(s_Multiplier_0_1_7), .S1(s_Multiplier_0_1_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_1_3 (.A0(Multiplier_0_pp_2_9), .A1(Multiplier_0_pp_2_10), 
           .B0(Multiplier_0_pp_3_9), .B1(Multiplier_0_pp_3_10), .CI(co_Multiplier_0_1_2), 
           .COUT(co_Multiplier_0_1_3), .S0(s_Multiplier_0_1_9), .S1(s_Multiplier_0_1_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_1_4 (.A0(Multiplier_0_pp_2_11), .A1(Multiplier_0_pp_2_12), 
           .B0(Multiplier_0_pp_3_11), .B1(Multiplier_0_pp_3_12), .CI(co_Multiplier_0_1_3), 
           .COUT(co_Multiplier_0_1_4), .S0(s_Multiplier_0_1_11), .S1(s_Multiplier_0_1_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_1_5 (.A0(Multiplier_0_pp_2_13), .A1(Multiplier_0_pp_2_14), 
           .B0(Multiplier_0_pp_3_13), .B1(Multiplier_0_pp_3_14), .CI(co_Multiplier_0_1_4), 
           .COUT(co_Multiplier_0_1_5), .S0(s_Multiplier_0_1_13), .S1(s_Multiplier_0_1_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_1_6 (.A0(Multiplier_0_pp_2_15), .A1(Multiplier_0_pp_2_16), 
           .B0(Multiplier_0_pp_3_15), .B1(Multiplier_0_pp_3_16), .CI(co_Multiplier_0_1_5), 
           .COUT(co_Multiplier_0_1_6), .S0(s_Multiplier_0_1_15), .S1(s_Multiplier_0_1_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_1_7 (.A0(Multiplier_0_pp_2_17), .A1(GND_net), 
           .B0(Multiplier_0_pp_3_17), .B1(Multiplier_0_pp_3_18), .CI(co_Multiplier_0_1_6), 
           .COUT(co_Multiplier_0_1_7), .S0(s_Multiplier_0_1_17), .S1(s_Multiplier_0_1_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_1_8 (.A0(GND_net), .A1(GND_net), .B0(Multiplier_0_pp_3_19), 
           .B1(GND_net), .CI(co_Multiplier_0_1_7), .COUT(co_Multiplier_0_1_8), 
           .S0(s_Multiplier_0_1_19), .S1(s_Multiplier_0_1_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_Multiplier_0_1_9 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_Multiplier_0_1_8), .S0(s_Multiplier_0_1_21)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_Multiplier_0_2_1 (.A0(GND_net), .A1(Multiplier_0_pp_4_10), 
           .B0(GND_net), .B1(Multiplier_0_pp_5_10), .CI(GND_net), .COUT(co_Multiplier_0_2_1), 
           .S1(s_Multiplier_0_2_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_2_2 (.A0(Multiplier_0_pp_4_11), .A1(Multiplier_0_pp_4_12), 
           .B0(Multiplier_0_pp_5_11), .B1(Multiplier_0_pp_5_12), .CI(co_Multiplier_0_2_1), 
           .COUT(co_Multiplier_0_2_2), .S0(s_Multiplier_0_2_11), .S1(s_Multiplier_0_2_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_2_3 (.A0(Multiplier_0_pp_4_13), .A1(Multiplier_0_pp_4_14), 
           .B0(Multiplier_0_pp_5_13), .B1(Multiplier_0_pp_5_14), .CI(co_Multiplier_0_2_2), 
           .COUT(co_Multiplier_0_2_3), .S0(s_Multiplier_0_2_13), .S1(s_Multiplier_0_2_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_2_4 (.A0(Multiplier_0_pp_4_15), .A1(Multiplier_0_pp_4_16), 
           .B0(Multiplier_0_pp_5_15), .B1(Multiplier_0_pp_5_16), .CI(co_Multiplier_0_2_3), 
           .COUT(co_Multiplier_0_2_4), .S0(s_Multiplier_0_2_15), .S1(s_Multiplier_0_2_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_2_5 (.A0(Multiplier_0_pp_4_17), .A1(Multiplier_0_pp_4_18), 
           .B0(Multiplier_0_pp_5_17), .B1(Multiplier_0_pp_5_18), .CI(co_Multiplier_0_2_4), 
           .COUT(co_Multiplier_0_2_5), .S0(s_Multiplier_0_2_17), .S1(s_Multiplier_0_2_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_2_6 (.A0(Multiplier_0_pp_4_19), .A1(Multiplier_0_pp_4_20), 
           .B0(Multiplier_0_pp_5_19), .B1(Multiplier_0_pp_5_20), .CI(co_Multiplier_0_2_5), 
           .COUT(co_Multiplier_0_2_6), .S0(s_Multiplier_0_2_19), .S1(s_Multiplier_0_2_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_2_7 (.A0(Multiplier_0_pp_4_21), .A1(GND_net), 
           .B0(Multiplier_0_pp_5_21), .B1(Multiplier_0_pp_5_22), .CI(co_Multiplier_0_2_6), 
           .COUT(co_Multiplier_0_2_7), .S0(s_Multiplier_0_2_21), .S1(s_Multiplier_0_2_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_2_8 (.A0(GND_net), .A1(GND_net), .B0(Multiplier_0_pp_5_23), 
           .B1(GND_net), .CI(co_Multiplier_0_2_7), .S0(s_Multiplier_0_2_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_Multiplier_0_3_1 (.A0(GND_net), .A1(f_s_Multiplier_0_0_4), 
           .B0(GND_net), .B1(f_Multiplier_0_pp_2_4), .CI(GND_net), .COUT(co_Multiplier_0_3_1), 
           .S1(rego_o_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_2 (.A0(f_s_Multiplier_0_0_5), .A1(f_s_Multiplier_0_0_6), 
           .B0(f_Multiplier_0_pp_2_5), .B1(f_s_Multiplier_0_1_6), .CI(co_Multiplier_0_3_1), 
           .COUT(co_Multiplier_0_3_2), .S0(rego_o_5), .S1(rego_o_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_3 (.A0(f_s_Multiplier_0_0_7), .A1(f_s_Multiplier_0_0_8), 
           .B0(f_s_Multiplier_0_1_7), .B1(f_s_Multiplier_0_1_8), .CI(co_Multiplier_0_3_2), 
           .COUT(co_Multiplier_0_3_3), .S0(rego_o_7), .S1(s_Multiplier_0_3_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_4 (.A0(f_s_Multiplier_0_0_9), .A1(f_s_Multiplier_0_0_10), 
           .B0(f_s_Multiplier_0_1_9), .B1(f_s_Multiplier_0_1_10), .CI(co_Multiplier_0_3_3), 
           .COUT(co_Multiplier_0_3_4), .S0(s_Multiplier_0_3_9), .S1(s_Multiplier_0_3_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_5 (.A0(f_s_Multiplier_0_0_11), .A1(f_s_Multiplier_0_0_12), 
           .B0(f_s_Multiplier_0_1_11), .B1(f_s_Multiplier_0_1_12), .CI(co_Multiplier_0_3_4), 
           .COUT(co_Multiplier_0_3_5), .S0(s_Multiplier_0_3_11), .S1(s_Multiplier_0_3_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_6 (.A0(f_s_Multiplier_0_0_13), .A1(f_s_Multiplier_0_0_14), 
           .B0(f_s_Multiplier_0_1_13), .B1(f_s_Multiplier_0_1_14), .CI(co_Multiplier_0_3_5), 
           .COUT(co_Multiplier_0_3_6), .S0(s_Multiplier_0_3_13), .S1(s_Multiplier_0_3_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_7 (.A0(f_s_Multiplier_0_0_15), .A1(f_s_Multiplier_0_0_16), 
           .B0(f_s_Multiplier_0_1_15), .B1(f_s_Multiplier_0_1_16), .CI(co_Multiplier_0_3_6), 
           .COUT(co_Multiplier_0_3_7), .S0(s_Multiplier_0_3_15), .S1(s_Multiplier_0_3_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_8 (.A0(f_s_Multiplier_0_0_17), .A1(GND_net), 
           .B0(f_s_Multiplier_0_1_17), .B1(f_s_Multiplier_0_1_18), .CI(co_Multiplier_0_3_7), 
           .COUT(co_Multiplier_0_3_8), .S0(s_Multiplier_0_3_17), .S1(s_Multiplier_0_3_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_9 (.A0(GND_net), .A1(GND_net), .B0(f_s_Multiplier_0_1_19), 
           .B1(f_s_Multiplier_0_1_20), .CI(co_Multiplier_0_3_8), .COUT(co_Multiplier_0_3_9), 
           .S0(s_Multiplier_0_3_19), .S1(s_Multiplier_0_3_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_10 (.A0(GND_net), .A1(GND_net), .B0(f_s_Multiplier_0_1_21), 
           .B1(GND_net), .CI(co_Multiplier_0_3_9), .COUT(co_Multiplier_0_3_10), 
           .S0(s_Multiplier_0_3_21), .S1(s_Multiplier_0_3_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_Multiplier_0_3_11 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_Multiplier_0_3_10), .S0(s_Multiplier_0_3_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_t_Multiplier_0_4_1 (.A0(GND_net), .A1(s_Multiplier_0_3_8), 
           .B0(GND_net), .B1(f_Multiplier_0_pp_4_8), .CI(GND_net), .COUT(co_t_Multiplier_0_4_1), 
           .S1(rego_o_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_2 (.A0(s_Multiplier_0_3_9), .A1(s_Multiplier_0_3_10), 
           .B0(f_Multiplier_0_pp_4_9), .B1(f_s_Multiplier_0_2_10), .CI(co_t_Multiplier_0_4_1), 
           .COUT(co_t_Multiplier_0_4_2), .S0(rego_o_9), .S1(rego_o_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_3 (.A0(s_Multiplier_0_3_11), .A1(s_Multiplier_0_3_12), 
           .B0(f_s_Multiplier_0_2_11), .B1(f_s_Multiplier_0_2_12), .CI(co_t_Multiplier_0_4_2), 
           .COUT(co_t_Multiplier_0_4_3), .S0(rego_o_11), .S1(rego_o_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_4 (.A0(s_Multiplier_0_3_13), .A1(s_Multiplier_0_3_14), 
           .B0(f_s_Multiplier_0_2_13), .B1(f_s_Multiplier_0_2_14), .CI(co_t_Multiplier_0_4_3), 
           .COUT(co_t_Multiplier_0_4_4), .S0(rego_o_13), .S1(rego_o_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_5 (.A0(s_Multiplier_0_3_15), .A1(s_Multiplier_0_3_16), 
           .B0(f_s_Multiplier_0_2_15), .B1(f_s_Multiplier_0_2_16), .CI(co_t_Multiplier_0_4_4), 
           .COUT(co_t_Multiplier_0_4_5), .S0(rego_o_15), .S1(rego_o_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_6 (.A0(s_Multiplier_0_3_17), .A1(s_Multiplier_0_3_18), 
           .B0(f_s_Multiplier_0_2_17), .B1(f_s_Multiplier_0_2_18), .CI(co_t_Multiplier_0_4_5), 
           .COUT(co_t_Multiplier_0_4_6), .S0(rego_o_17), .S1(rego_o_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_7 (.A0(s_Multiplier_0_3_19), .A1(s_Multiplier_0_3_20), 
           .B0(f_s_Multiplier_0_2_19), .B1(f_s_Multiplier_0_2_20), .CI(co_t_Multiplier_0_4_6), 
           .COUT(co_t_Multiplier_0_4_7), .S0(rego_o_19), .S1(rego_o_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_8 (.A0(s_Multiplier_0_3_21), .A1(s_Multiplier_0_3_22), 
           .B0(f_s_Multiplier_0_2_21), .B1(f_s_Multiplier_0_2_22), .CI(co_t_Multiplier_0_4_7), 
           .COUT(co_t_Multiplier_0_4_8), .S0(rego_o_21), .S1(rego_o_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_9 (.A0(s_Multiplier_0_3_23), .A1(GND_net), 
           .B0(f_s_Multiplier_0_2_23), .B1(GND_net), .CI(co_t_Multiplier_0_4_8), 
           .S0(rego_o_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_0_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(Multiplier_0_cin_lr_0), .CO(mco), .P0(Multiplier_0_pp_0_1), 
          .P1(Multiplier_0_pp_0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_0_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco), .CO(mco_1), .P0(Multiplier_0_pp_0_3), 
          .P1(Multiplier_0_pp_0_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_0_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco_1), .CO(mco_2), .P0(Multiplier_0_pp_0_5), 
          .P1(Multiplier_0_pp_0_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_0_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco_2), .CO(mco_3), .P0(Multiplier_0_pp_0_7), 
          .P1(Multiplier_0_pp_0_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_0_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco_3), .CO(mco_4), .P0(Multiplier_0_pp_0_9), 
          .P1(Multiplier_0_pp_0_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_0_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_0_5_n2), 
          .A2(Multiplier_0_mult_0_5_n1), .A3(VCC_net), .B0(regb_b_1), 
          .B1(VCC_net), .B2(VCC_net), .B3(VCC_net), .CI(mco_4), .CO(mfco), 
          .P0(Multiplier_0_pp_0_11), .P1(Multiplier_0_pp_0_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_2_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(Multiplier_0_cin_lr_2), .CO(mco_5), .P0(Multiplier_0_pp_1_3), 
          .P1(Multiplier_0_pp_1_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_2_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_5), .CO(mco_6), .P0(Multiplier_0_pp_1_5), 
          .P1(Multiplier_0_pp_1_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_2_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_6), .CO(mco_7), .P0(Multiplier_0_pp_1_7), 
          .P1(Multiplier_0_pp_1_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_2_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_7), .CO(mco_8), .P0(Multiplier_0_pp_1_9), 
          .P1(Multiplier_0_pp_1_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_2_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_8), .CO(mco_9), .P0(Multiplier_0_pp_1_11), 
          .P1(Multiplier_0_pp_1_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_2_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_2_5_n2), 
          .A2(Multiplier_0_mult_2_5_n1), .A3(GND_net), .B0(regb_b_3), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_2), .CI(mco_9), .CO(mfco_1), 
          .P0(Multiplier_0_pp_1_13), .P1(Multiplier_0_pp_1_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_4_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(Multiplier_0_cin_lr_4), .CO(mco_10), .P0(Multiplier_0_pp_2_5), 
          .P1(Multiplier_0_pp_2_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_4_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_10), .CO(mco_11), .P0(Multiplier_0_pp_2_7), 
          .P1(Multiplier_0_pp_2_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_4_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_11), .CO(mco_12), .P0(Multiplier_0_pp_2_9), 
          .P1(Multiplier_0_pp_2_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_4_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_12), .CO(mco_13), .P0(Multiplier_0_pp_2_11), 
          .P1(Multiplier_0_pp_2_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_4_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_13), .CO(mco_14), .P0(Multiplier_0_pp_2_13), 
          .P1(Multiplier_0_pp_2_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_4_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_4_5_n2), 
          .A2(Multiplier_0_mult_4_5_n1), .A3(GND_net), .B0(regb_b_5), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_4), .CI(mco_14), .CO(mfco_2), 
          .P0(Multiplier_0_pp_2_15), .P1(Multiplier_0_pp_2_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_6_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(Multiplier_0_cin_lr_6), .CO(mco_15), .P0(Multiplier_0_pp_3_7), 
          .P1(Multiplier_0_pp_3_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_6_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_15), .CO(mco_16), .P0(Multiplier_0_pp_3_9), 
          .P1(Multiplier_0_pp_3_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_6_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_16), .CO(mco_17), .P0(Multiplier_0_pp_3_11), 
          .P1(Multiplier_0_pp_3_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_6_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_17), .CO(mco_18), .P0(Multiplier_0_pp_3_13), 
          .P1(Multiplier_0_pp_3_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_6_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_18), .CO(mco_19), .P0(Multiplier_0_pp_3_15), 
          .P1(Multiplier_0_pp_3_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_6_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_6_5_n2), 
          .A2(Multiplier_0_mult_6_5_n1), .A3(GND_net), .B0(regb_b_7), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_6), .CI(mco_19), .CO(mfco_3), 
          .P0(Multiplier_0_pp_3_17), .P1(Multiplier_0_pp_3_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_8_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(Multiplier_0_cin_lr_8), .CO(mco_20), .P0(Multiplier_0_pp_4_9), 
          .P1(Multiplier_0_pp_4_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_8_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_20), .CO(mco_21), .P0(Multiplier_0_pp_4_11), 
          .P1(Multiplier_0_pp_4_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_8_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_21), .CO(mco_22), .P0(Multiplier_0_pp_4_13), 
          .P1(Multiplier_0_pp_4_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_8_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_22), .CO(mco_23), .P0(Multiplier_0_pp_4_15), 
          .P1(Multiplier_0_pp_4_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_8_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_23), .CO(mco_24), .P0(Multiplier_0_pp_4_17), 
          .P1(Multiplier_0_pp_4_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_8_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_8_5_n2), 
          .A2(Multiplier_0_mult_8_5_n1), .A3(GND_net), .B0(regb_b_9), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_8), .CI(mco_24), .CO(mfco_4), 
          .P0(Multiplier_0_pp_4_19), .P1(Multiplier_0_pp_4_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_10_0 (.A0(Multiplier_0_mult_10_0_n0), .A1(rega_a_1), 
          .A2(Multiplier_0_mult_10_0_n1), .A3(rega_a_2), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(Multiplier_0_cin_lr_10), 
          .CO(mco_25), .P0(Multiplier_0_pp_5_11), .P1(Multiplier_0_pp_5_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_10_1 (.A0(Multiplier_0_mult_10_1_n0), .A1(rega_a_3), 
          .A2(Multiplier_0_mult_10_1_n1), .A3(rega_a_4), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_25), 
          .CO(mco_26), .P0(Multiplier_0_pp_5_13), .P1(Multiplier_0_pp_5_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_10_2 (.A0(Multiplier_0_mult_10_2_n0), .A1(rega_a_5), 
          .A2(Multiplier_0_mult_10_2_n1), .A3(rega_a_6), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_26), 
          .CO(mco_27), .P0(Multiplier_0_pp_5_15), .P1(Multiplier_0_pp_5_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_10_3 (.A0(Multiplier_0_mult_10_3_n0), .A1(rega_a_7), 
          .A2(Multiplier_0_mult_10_3_n1), .A3(rega_a_8), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_27), 
          .CO(mco_28), .P0(Multiplier_0_pp_5_17), .P1(Multiplier_0_pp_5_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_10_4 (.A0(Multiplier_0_mult_10_4_n0), .A1(rega_a_9), 
          .A2(Multiplier_0_mult_10_4_n1), .A3(rega_a_10), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_28), 
          .CO(mco_29), .P0(Multiplier_0_pp_5_19), .P1(Multiplier_0_pp_5_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_10_5 (.A0(Multiplier_0_mult_10_5_n0), .A1(Multiplier_0_mult_10_5_n2), 
          .A2(rega_a_11), .A3(GND_net), .B0(VCC_net), .B1(VCC_net), 
          .B2(regb_b_11), .B3(regb_b_10), .CI(mco_29), .CO(mfco_5), 
          .P0(Multiplier_0_pp_5_21), .P1(Multiplier_0_pp_5_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t26 (.A(rega_a_11), .B(regb_b_0), .Z(Multiplier_0_mult_0_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    AND2 AND2_t27 (.A(regb_b_0), .B(regb_b_0), .Z(Multiplier_0_pp_0_0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(376[10:72])
    ND2 ND2_t23 (.A(rega_a_11), .B(regb_b_2), .Z(Multiplier_0_mult_2_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t20 (.A(rega_a_11), .B(regb_b_4), .Z(Multiplier_0_mult_4_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t17 (.A(rega_a_11), .B(regb_b_6), .Z(Multiplier_0_mult_6_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t14 (.A(rega_a_11), .B(regb_b_8), .Z(Multiplier_0_mult_8_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t11 (.A(rega_a_1), .B(regb_b_11), .Z(Multiplier_0_mult_10_0_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    
endmodule
