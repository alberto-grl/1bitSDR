// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.10.2.115
// Netlist written on Mon Nov 26 21:33:53 2018
//
// Verilog Description of module Mixer
//

module Mixer (clk, RFIn, sin_in, cos_in, MixerOutSin, MixerOutCos) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/fpgasdr/mixer.v(2[8:13])
    input clk;   // c:/users/user/lattice/fpgasdr/mixer.v(11[7:10])
    input RFIn;   // c:/users/user/lattice/fpgasdr/mixer.v(14[7:11])
    input [1:0]sin_in;   // c:/users/user/lattice/fpgasdr/mixer.v(12[13:19])
    input [1:0]cos_in;   // c:/users/user/lattice/fpgasdr/mixer.v(13[13:19])
    output [63:0]MixerOutSin;   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    output [63:0]MixerOutCos;   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    
    wire clk_c /* synthesis is_clock=1, SET_AS_NETWORK=clk_c */ ;   // c:/users/user/lattice/fpgasdr/mixer.v(11[7:10])
    
    wire GND_net, RFIn_c, MixerOutSin_c_0, RFInR1, VCC_net;
    
    VHI i16 (.Z(VCC_net));
    FD1S3AX RFInR1_6 (.D(RFIn_c), .CK(clk_c), .Q(RFInR1));   // c:/users/user/lattice/fpgasdr/mixer.v(20[8] 24[7])
    defparam RFInR1_6.GSR = "ENABLED";
    TSALL TSALL_INST (.TSALL(GND_net));
    OB MixerOutSin_pad_63 (.I(GND_net), .O(MixerOutSin[63]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_62 (.I(GND_net), .O(MixerOutSin[62]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_61 (.I(GND_net), .O(MixerOutSin[61]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_60 (.I(GND_net), .O(MixerOutSin[60]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_59 (.I(GND_net), .O(MixerOutSin[59]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_58 (.I(GND_net), .O(MixerOutSin[58]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_57 (.I(GND_net), .O(MixerOutSin[57]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_56 (.I(GND_net), .O(MixerOutSin[56]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_55 (.I(GND_net), .O(MixerOutSin[55]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_54 (.I(GND_net), .O(MixerOutSin[54]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_53 (.I(GND_net), .O(MixerOutSin[53]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_52 (.I(GND_net), .O(MixerOutSin[52]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_51 (.I(GND_net), .O(MixerOutSin[51]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_50 (.I(GND_net), .O(MixerOutSin[50]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_49 (.I(GND_net), .O(MixerOutSin[49]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_48 (.I(GND_net), .O(MixerOutSin[48]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_47 (.I(GND_net), .O(MixerOutSin[47]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_46 (.I(GND_net), .O(MixerOutSin[46]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_45 (.I(GND_net), .O(MixerOutSin[45]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_44 (.I(GND_net), .O(MixerOutSin[44]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_43 (.I(GND_net), .O(MixerOutSin[43]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_42 (.I(GND_net), .O(MixerOutSin[42]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_41 (.I(GND_net), .O(MixerOutSin[41]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_40 (.I(GND_net), .O(MixerOutSin[40]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_39 (.I(GND_net), .O(MixerOutSin[39]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_38 (.I(GND_net), .O(MixerOutSin[38]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_37 (.I(GND_net), .O(MixerOutSin[37]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_36 (.I(GND_net), .O(MixerOutSin[36]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_35 (.I(GND_net), .O(MixerOutSin[35]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_34 (.I(GND_net), .O(MixerOutSin[34]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_33 (.I(GND_net), .O(MixerOutSin[33]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_32 (.I(GND_net), .O(MixerOutSin[32]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_31 (.I(GND_net), .O(MixerOutSin[31]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_30 (.I(GND_net), .O(MixerOutSin[30]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_29 (.I(GND_net), .O(MixerOutSin[29]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_28 (.I(GND_net), .O(MixerOutSin[28]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_27 (.I(GND_net), .O(MixerOutSin[27]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_26 (.I(GND_net), .O(MixerOutSin[26]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_25 (.I(GND_net), .O(MixerOutSin[25]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_24 (.I(GND_net), .O(MixerOutSin[24]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_23 (.I(GND_net), .O(MixerOutSin[23]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_22 (.I(GND_net), .O(MixerOutSin[22]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_21 (.I(GND_net), .O(MixerOutSin[21]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_20 (.I(GND_net), .O(MixerOutSin[20]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_19 (.I(GND_net), .O(MixerOutSin[19]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_18 (.I(GND_net), .O(MixerOutSin[18]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_17 (.I(GND_net), .O(MixerOutSin[17]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_16 (.I(GND_net), .O(MixerOutSin[16]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_15 (.I(GND_net), .O(MixerOutSin[15]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_14 (.I(GND_net), .O(MixerOutSin[14]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_13 (.I(GND_net), .O(MixerOutSin[13]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_12 (.I(GND_net), .O(MixerOutSin[12]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_11 (.I(GND_net), .O(MixerOutSin[11]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_10 (.I(GND_net), .O(MixerOutSin[10]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_9 (.I(GND_net), .O(MixerOutSin[9]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_8 (.I(GND_net), .O(MixerOutSin[8]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_7 (.I(GND_net), .O(MixerOutSin[7]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_6 (.I(GND_net), .O(MixerOutSin[6]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_5 (.I(GND_net), .O(MixerOutSin[5]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_4 (.I(GND_net), .O(MixerOutSin[4]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_3 (.I(GND_net), .O(MixerOutSin[3]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_2 (.I(GND_net), .O(MixerOutSin[2]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_1 (.I(GND_net), .O(MixerOutSin[1]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutSin_pad_0 (.I(MixerOutSin_c_0), .O(MixerOutSin[0]));   // c:/users/user/lattice/fpgasdr/mixer.v(15[15:26])
    OB MixerOutCos_pad_63 (.I(GND_net), .O(MixerOutCos[63]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_62 (.I(GND_net), .O(MixerOutCos[62]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_61 (.I(GND_net), .O(MixerOutCos[61]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_60 (.I(GND_net), .O(MixerOutCos[60]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_59 (.I(GND_net), .O(MixerOutCos[59]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_58 (.I(GND_net), .O(MixerOutCos[58]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_57 (.I(GND_net), .O(MixerOutCos[57]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_56 (.I(GND_net), .O(MixerOutCos[56]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_55 (.I(GND_net), .O(MixerOutCos[55]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_54 (.I(GND_net), .O(MixerOutCos[54]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_53 (.I(GND_net), .O(MixerOutCos[53]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_52 (.I(GND_net), .O(MixerOutCos[52]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_51 (.I(GND_net), .O(MixerOutCos[51]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_50 (.I(GND_net), .O(MixerOutCos[50]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_49 (.I(GND_net), .O(MixerOutCos[49]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_48 (.I(GND_net), .O(MixerOutCos[48]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_47 (.I(GND_net), .O(MixerOutCos[47]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_46 (.I(GND_net), .O(MixerOutCos[46]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_45 (.I(GND_net), .O(MixerOutCos[45]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_44 (.I(GND_net), .O(MixerOutCos[44]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_43 (.I(GND_net), .O(MixerOutCos[43]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_42 (.I(GND_net), .O(MixerOutCos[42]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_41 (.I(GND_net), .O(MixerOutCos[41]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_40 (.I(GND_net), .O(MixerOutCos[40]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_39 (.I(GND_net), .O(MixerOutCos[39]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_38 (.I(GND_net), .O(MixerOutCos[38]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_37 (.I(GND_net), .O(MixerOutCos[37]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_36 (.I(GND_net), .O(MixerOutCos[36]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_35 (.I(GND_net), .O(MixerOutCos[35]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_34 (.I(GND_net), .O(MixerOutCos[34]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_33 (.I(GND_net), .O(MixerOutCos[33]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_32 (.I(GND_net), .O(MixerOutCos[32]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_31 (.I(GND_net), .O(MixerOutCos[31]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_30 (.I(GND_net), .O(MixerOutCos[30]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_29 (.I(GND_net), .O(MixerOutCos[29]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_28 (.I(GND_net), .O(MixerOutCos[28]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_27 (.I(GND_net), .O(MixerOutCos[27]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_26 (.I(GND_net), .O(MixerOutCos[26]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_25 (.I(GND_net), .O(MixerOutCos[25]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_24 (.I(GND_net), .O(MixerOutCos[24]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_23 (.I(GND_net), .O(MixerOutCos[23]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_22 (.I(GND_net), .O(MixerOutCos[22]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_21 (.I(GND_net), .O(MixerOutCos[21]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_20 (.I(GND_net), .O(MixerOutCos[20]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_19 (.I(GND_net), .O(MixerOutCos[19]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_18 (.I(GND_net), .O(MixerOutCos[18]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_17 (.I(GND_net), .O(MixerOutCos[17]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_16 (.I(GND_net), .O(MixerOutCos[16]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_15 (.I(GND_net), .O(MixerOutCos[15]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_14 (.I(GND_net), .O(MixerOutCos[14]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_13 (.I(GND_net), .O(MixerOutCos[13]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_12 (.I(GND_net), .O(MixerOutCos[12]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_11 (.I(GND_net), .O(MixerOutCos[11]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_10 (.I(GND_net), .O(MixerOutCos[10]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_9 (.I(GND_net), .O(MixerOutCos[9]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_8 (.I(GND_net), .O(MixerOutCos[8]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_7 (.I(GND_net), .O(MixerOutCos[7]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_6 (.I(GND_net), .O(MixerOutCos[6]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_5 (.I(GND_net), .O(MixerOutCos[5]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_4 (.I(GND_net), .O(MixerOutCos[4]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_3 (.I(GND_net), .O(MixerOutCos[3]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_2 (.I(GND_net), .O(MixerOutCos[2]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_1 (.I(GND_net), .O(MixerOutCos[1]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    OB MixerOutCos_pad_0 (.I(GND_net), .O(MixerOutCos[0]));   // c:/users/user/lattice/fpgasdr/mixer.v(16[15:26])
    IB clk_pad (.I(clk), .O(clk_c));   // c:/users/user/lattice/fpgasdr/mixer.v(11[7:10])
    IB RFIn_pad (.I(RFIn), .O(RFIn_c));   // c:/users/user/lattice/fpgasdr/mixer.v(14[7:11])
    GSR GSR_INST (.GSR(VCC_net));
    FD1S3AX RFInR_7 (.D(RFInR1), .CK(clk_c), .Q(MixerOutSin_c_0));   // c:/users/user/lattice/fpgasdr/mixer.v(20[8] 24[7])
    defparam RFInR_7.GSR = "ENABLED";
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    VLO i1 (.Z(GND_net));
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

