// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.11.2.446
// Netlist written on Sun Apr 05 22:59:51 2020
//
// Verilog Description of module top
//

module top (i_Rx_Serial, o_Tx_Serial, o_Rx_DV, o_Rx_Byte, MYLED, XOut, 
            RFIn, DiffOut, PWMOut, PWMOutP1, PWMOutP2, PWMOutP3, 
            PWMOutP4, PWMOutN1, PWMOutN2, PWMOutN3, PWMOutN4, sinGen, 
            sin_out, CIC_out_clkSin) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(45[8:11])
    input i_Rx_Serial;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(47[13:24])
    output o_Tx_Serial;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(48[11:22])
    output o_Rx_DV;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(49[13:20])
    output [7:0]o_Rx_Byte;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[16:25])
    output [7:0]MYLED;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(51[18:23])
    output XOut;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(55[9:13])
    input RFIn;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(56[9:13])
    output DiffOut;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(57[9:16])
    output PWMOut;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(58[9:15])
    output PWMOutP1;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(59[9:17])
    output PWMOutP2;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(60[9:17])
    output PWMOutP3;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(61[9:17])
    output PWMOutP4;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(62[9:17])
    output PWMOutN1;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(63[9:17])
    output PWMOutN2;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(64[9:17])
    output PWMOutN3;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(65[9:17])
    output PWMOutN4;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(66[9:17])
    output sinGen;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(67[9:15])
    output sin_out;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(68[9:16])
    output CIC_out_clkSin;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(69[9:23])
    
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(71[8:15])
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(82[6:21])
    
    wire GND_net, VCC_net, i_Rx_Serial_c, o_Rx_DV_c, o_Rx_Byte_c_7, 
        o_Rx_Byte_c_6, o_Rx_Byte_c_5, o_Rx_Byte_c_4, o_Rx_Byte_c_3, 
        o_Rx_Byte_c_2, n7349, o_Rx_Byte_c_0, MYLED_c_5, MYLED_c_4, 
        MYLED_c_3, MYLED_c_2, MYLED_c_1, MYLED_c_0, RFIn_c, DiffOut_c, 
        PWMOutP4_c, PWMOutN4_c, sinGen_c, n2303;
    wire [11:0]MixerOutSin;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(78[20:31])
    wire [11:0]MixerOutCos;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(79[20:31])
    wire [11:0]CIC1_outSin;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(81[20:31])
    wire [11:0]CIC1_outCos;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(84[20:31])
    wire [63:0]phase_accum;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(86[13:24])
    wire [12:0]LOSine;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(87[20:26])
    wire [12:0]LOCosine;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(88[20:28])
    wire [63:0]phase_inc_carrGen;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(90[19:36])
    wire [63:0]phase_inc_carrGen1;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(91[19:37])
    wire [11:0]DemodOut;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(94[20:28])
    wire [7:0]CICGain;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(96[11:18])
    
    wire n1134, n1133, n1132, n1131, n1130, n1129, n1128, n1127, 
        n1126, n1125, n1124, n1123, n1122, n1121, n1120, n1119, 
        n1118, n1117, n1116, n1115, n1114, n1113, n1112, n1111, 
        n1110, n1109, n1108, n1107, n1106, n1105, n1104, n1103, 
        n1102, n1101, n1100, n1099, n1098, n1097, n1096, n1095, 
        n1094, n1093, n1092, n1091, n1090, n1089, n1088, n1087, 
        n1086, n1085, n1084, n1083, n1082, n1081, n1080, n1079, 
        n1078, n1077, n1076, n1072, n1073, n1074, n1075, n7733, 
        n7735, n2364, n2359, n2353, n1012, n1011, n1013, n1014, 
        n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
        n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, 
        n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, 
        n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, 
        n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, 
        n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
        n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, 
        n11340, n11339, n11338, n11337, n11336, n11335, n11334, 
        n11333, n11332, n11331, n11330, n11329, n11328, n11327, 
        n11326, n11325, n11324, n11323, n11322, n11321, n11320, 
        n11319, n11318, n11317, n11316, n11315, n11314, n11313, 
        n11312, n11311, n11310, n11302, n11301, n11300, n11299, 
        n11298, n11297, n11296, n11295, n11294, n11293, n11292, 
        n11291, n11290, n11289, n11288, n11287, n11286, n11285, 
        n11284, n11283, n11282, n11281, n11280, n11279, n11278, 
        n11277, n11276, n11275, n11274, n11273, n11272, n11271, 
        n11129, n11128, n11127, n11126, n11125, n11124, n11123, 
        n11122, n11121, n11120, n11119, n11118, n11117, n11116, 
        n11115, n11114, n11113, n11112, n11111, n11110, n11109, 
        n11108, n11107, n11106, n11105, n11104, n11103, n11102, 
        n11101, n11100;
    wire [71:0]d10_adj_2550;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(47[26:29])
    wire [71:0]d_out_11__N_1819_adj_2575;
    
    wire n9571, n9593, n9591;
    wire [11:0]DataInReg_11__N_1856;
    
    wire n2305, n9589, n2302, n9547, n2300, n2299, n2298, n2297, 
        n2296, n2295, n2294, n2293, n2292, n2291, n2289, n13375, 
        n2288, n2287, n13376, n2286, n12803, n12931, n2285, n2284, 
        n2283, n2282, n3663, n3653, n3632, n3628, n3614, n6, 
        n2306, n2307, n12879, n13381, n2308, n2304, n13380, n9527, 
        n28, n29, n30, n2341, n2340, n2339, n2338, n2337, n2334, 
        n2333, n2332, n2331, n2330, n2328, n2327, n2326, n2324, 
        n8225, n2531, n2530, n2521, n2513, osc_clk_enable_1397, 
        n8016, n2492, n2486, n2485, n13390, n2608, n9535, osc_clk_enable_128, 
        n2860, n2859, n2858, n2857, n2856, n2855, n2854, n2853, 
        n2852, n2851, n2850, n2849, n2848, n2847, n2846, n2845, 
        n2844, n2843, n2842, n2841, n2840, n2839, n2838, n2837, 
        n2836, n2835, n2834, n2833, n2832, n2831, n2830, n2829, 
        n2828, n2827, n2826, n2825, n2824, n2823, n2822, n9000, 
        n61, n62, n63, n64, n65, n66, n67, n68, n70, n13411, 
        n2322, n2321, n2320, n2319, n2318, n2317, n2316, n2315, 
        n2314, n2313, n2312, n2311, n2310, n2309, n12919, n2821, 
        n2820, n2819, n2818, n2817, n2816, n2815, n2814, n2813, 
        n2812, n2811, n2810, n2809, n2808, n2807, n2806, n2805, 
        n2804, n2803, n2802, n2801, n2800, n2799, n2798, n2797, 
        n2795, osc_clk_enable_1457, n12970, osc_clk_enable_1447, n13372, 
        n13523, n13385, n13384, osc_clk_enable_1394, n13291, n7739, 
        n7741, n7743, n7749, n7751, n7755, n7759, n7763, n7765, 
        n7767, n7769, n7771, n7773, n7777, n7779, n7781, n7783, 
        n7785, n7787, n7789, n7791, n7793, n7795, n7799, n7801, 
        n7803, n7805, n7807, n7809, n7813, n7817, n7819, n7825, 
        n7827, n7829, n8341, n13383, n9563, n8014, n8012, n8010, 
        n8008, n8006, n7970, n8004, n8002, n8000;
    
    VHI i2 (.Z(VCC_net));
    PUR PUR_INST (.PUR(VCC_net)) /* synthesis syn_instantiated=1 */ ;
    defparam PUR_INST.RST_PULSE = 1;
    OSCH OSCH_inst (.STDBY(GND_net), .OSC(osc_clk)) /* synthesis syn_instantiated=1 */ ;
    defparam OSCH_inst.NOM_FREQ = "88.67";
    FD1S3AX phase_inc_carrGen1_i0 (.D(phase_inc_carrGen[0]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[0]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i0.GSR = "ENABLED";
    PWM PWM1 (.osc_clk(osc_clk), .\DataInReg_11__N_1856[0] (DataInReg_11__N_1856[0]), 
        .PWMOutP4_c(PWMOutP4_c), .GND_net(GND_net), .\DataInReg_11__N_1856[1] (DataInReg_11__N_1856[1]), 
        .\DataInReg_11__N_1856[2] (DataInReg_11__N_1856[2]), .\DataInReg_11__N_1856[3] (DataInReg_11__N_1856[3]), 
        .\DataInReg_11__N_1856[4] (DataInReg_11__N_1856[4]), .\DataInReg_11__N_1856[5] (DataInReg_11__N_1856[5]), 
        .\DataInReg_11__N_1856[6] (DataInReg_11__N_1856[6]), .\DataInReg_11__N_1856[7] (DataInReg_11__N_1856[7]), 
        .\DataInReg_11__N_1856[8] (DataInReg_11__N_1856[8]), .\DemodOut[9] (DemodOut[9])) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(186[5] 192[2])
    LUT4 mux_318_i55_4_lut (.A(n7819), .B(n1081), .C(n13376), .D(n13375), 
         .Z(n2288)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i55_4_lut.init = 16'hcfca;
    FD1S3AX phase_inc_carrGen1_i48 (.D(phase_inc_carrGen[48]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[48]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i48.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i47 (.D(phase_inc_carrGen[47]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[47]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i47.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i46 (.D(phase_inc_carrGen[46]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[46]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i46.GSR = "ENABLED";
    LUT4 i1806_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1014), .Z(n7829)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1806_3_lut_4_lut.init = 16'hfb0b;
    FD1P3AX CICGain__i1 (.D(o_Rx_Byte_c_0), .SP(osc_clk_enable_1394), .CK(osc_clk), 
            .Q(CICGain[0]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam CICGain__i1.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i45 (.D(phase_inc_carrGen[45]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[45]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i45.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i44 (.D(phase_inc_carrGen[44]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[44]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i44.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i43 (.D(phase_inc_carrGen[43]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[43]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i43.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i42 (.D(phase_inc_carrGen[42]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[42]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i42.GSR = "ENABLED";
    OB o_Rx_Byte_pad_7 (.I(o_Rx_Byte_c_7), .O(o_Rx_Byte[7]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[16:25])
    FD1S3AX phase_inc_carrGen1_i41 (.D(phase_inc_carrGen[41]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[41]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i41.GSR = "ENABLED";
    LUT4 i1802_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1016), .Z(n7825)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1802_3_lut_4_lut.init = 16'hfb0b;
    FD1S3AX phase_inc_carrGen1_i40 (.D(phase_inc_carrGen[40]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[40]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i40.GSR = "ENABLED";
    LUT4 mux_318_i56_4_lut (.A(n2353), .B(n1080), .C(n13376), .D(n7970), 
         .Z(n2287)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i56_4_lut.init = 16'hcfca;
    FD1S3AX phase_inc_carrGen1_i39 (.D(phase_inc_carrGen[39]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[39]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i39.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i38 (.D(phase_inc_carrGen[38]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[38]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i38.GSR = "ENABLED";
    LUT4 i2967_2_lut (.A(n1019), .B(o_Rx_Byte_c_3), .Z(n2353)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i2967_2_lut.init = 16'h8888;
    FD1S3AX phase_inc_carrGen1_i37 (.D(phase_inc_carrGen[37]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[37]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i37.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i36 (.D(phase_inc_carrGen[36]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[36]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i36.GSR = "ENABLED";
    LUT4 i1975_4_lut (.A(n1083), .B(n1022), .C(o_Rx_Byte_c_3), .D(n13383), 
         .Z(n8010)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1975_4_lut.init = 16'hcac0;
    FD1S3AX phase_inc_carrGen1_i35 (.D(phase_inc_carrGen[35]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[35]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i35.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i34 (.D(phase_inc_carrGen[34]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[34]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i34.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i33 (.D(phase_inc_carrGen[33]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[33]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i33.GSR = "ENABLED";
    LUT4 i1804_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1015), .Z(n7827)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1804_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i1754_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1044), .Z(n7777)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i1754_3_lut_4_lut.init = 16'hf808;
    LUT4 i1796_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1020), .Z(n7819)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1796_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i1784_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1027), .Z(n7807)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1784_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_318_i44_4_lut (.A(n7801), .B(n1092), .C(n13376), .D(n13375), 
         .Z(n2299)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i44_4_lut.init = 16'hc0ca;
    LUT4 mux_318_i54_4_lut (.A(n7817), .B(n1082), .C(n13376), .D(n13375), 
         .Z(n2289)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i54_4_lut.init = 16'hc0ca;
    LUT4 mux_318_i51_4_lut (.A(n2492), .B(n1085), .C(n13376), .D(n13375), 
         .Z(n2292)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i51_4_lut.init = 16'hcfca;
    FD1S3AX phase_inc_carrGen1_i32 (.D(phase_inc_carrGen[32]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[32]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i32.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i31 (.D(phase_inc_carrGen[31]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[31]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i31.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i30 (.D(phase_inc_carrGen[30]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[30]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i30.GSR = "ENABLED";
    VLO i1 (.Z(GND_net));
    FD1S3AX phase_inc_carrGen1_i29 (.D(phase_inc_carrGen[29]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[29]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i29.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i28 (.D(phase_inc_carrGen[28]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[28]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i28.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i27 (.D(phase_inc_carrGen[27]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[27]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i27.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i26 (.D(phase_inc_carrGen[26]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[26]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i26.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i25 (.D(phase_inc_carrGen[25]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[25]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i25.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i24 (.D(phase_inc_carrGen[24]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[24]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i24.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i23 (.D(phase_inc_carrGen[23]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[23]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i23.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i22 (.D(phase_inc_carrGen[22]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[22]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i22.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i21 (.D(phase_inc_carrGen[21]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[21]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i21.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i20 (.D(phase_inc_carrGen[20]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[20]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i20.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i19 (.D(phase_inc_carrGen[19]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[19]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i19.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i18 (.D(phase_inc_carrGen[18]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[18]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i18.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i17 (.D(phase_inc_carrGen[17]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[17]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i17.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i16 (.D(phase_inc_carrGen[16]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[16]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i16.GSR = "ENABLED";
    LUT4 i3027_2_lut (.A(n1024), .B(o_Rx_Byte_c_3), .Z(n2492)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i3027_2_lut.init = 16'h8888;
    LUT4 mux_318_i52_4_lut (.A(n7813), .B(n1084), .C(n13376), .D(n13375), 
         .Z(n2291)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i52_4_lut.init = 16'hc0ca;
    LUT4 mux_318_i41_4_lut (.A(n13375), .B(n1095), .C(n13376), .D(n30), 
         .Z(n2302)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i41_4_lut.init = 16'hcfca;
    LUT4 i1778_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1031), .Z(n7801)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1778_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i1973_4_lut (.A(n1094), .B(n1033), .C(o_Rx_Byte_c_3), .D(n13383), 
         .Z(n8008)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1973_4_lut.init = 16'hcac0;
    FD1S3AX phase_inc_carrGen1_i15 (.D(phase_inc_carrGen[15]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[15]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i15.GSR = "ENABLED";
    LUT4 i1758_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1042), .Z(n7781)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1758_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i1760_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1041), .Z(n7783)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1760_3_lut_4_lut.init = 16'hfb0b;
    FD1S3AX phase_inc_carrGen1_i14 (.D(phase_inc_carrGen[14]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[14]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i14.GSR = "ENABLED";
    TSALL TSALL_INST (.TSALL(GND_net));
    FD1S3AX phase_inc_carrGen1_i13 (.D(phase_inc_carrGen[13]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[13]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i13.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i12 (.D(phase_inc_carrGen[12]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[12]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i12.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i11 (.D(phase_inc_carrGen[11]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[11]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i11.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i10 (.D(phase_inc_carrGen[10]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[10]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i10.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i9 (.D(phase_inc_carrGen[9]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[9]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i9.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i8 (.D(phase_inc_carrGen[8]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[8]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i8.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i7 (.D(phase_inc_carrGen[7]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[7]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i7.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i6 (.D(phase_inc_carrGen[6]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[6]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i6.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i5 (.D(phase_inc_carrGen[5]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[5]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i5.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i4 (.D(phase_inc_carrGen[4]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[4]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i4.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i3 (.D(phase_inc_carrGen[3]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[3]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i3.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i2 (.D(phase_inc_carrGen[2]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[2]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i2.GSR = "ENABLED";
    OB o_Rx_Byte_pad_6 (.I(o_Rx_Byte_c_6), .O(o_Rx_Byte[6]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[16:25])
    FD1S3AX phase_inc_carrGen1_i1 (.D(phase_inc_carrGen[1]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[1]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i1.GSR = "ENABLED";
    LUT4 i1768_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1037), .Z(n7791)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;
    defparam i1768_3_lut_4_lut.init = 16'hf707;
    LUT4 i1776_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1032), .Z(n7799)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i1776_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_318_i49_4_lut (.A(n7809), .B(n1087), .C(n13376), .D(n13375), 
         .Z(n2294)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i49_4_lut.init = 16'hc0ca;
    LUT4 mux_318_i50_4_lut (.A(n2359), .B(n1086), .C(n13376), .D(n7970), 
         .Z(n2293)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i50_4_lut.init = 16'hcfca;
    LUT4 i1_2_lut_rep_73_3_lut_3_lut_3_lut (.A(o_Rx_Byte_c_0), .B(n7349), 
         .C(o_Rx_Byte_c_4), .Z(n13384)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i1_2_lut_rep_73_3_lut_3_lut_3_lut.init = 16'h0404;
    LUT4 i1_2_lut_rep_70_3_lut_4_lut_4_lut_4_lut (.A(o_Rx_Byte_c_0), .B(n7349), 
         .C(n8225), .D(o_Rx_Byte_c_4), .Z(n13381)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_rep_70_3_lut_4_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i2966_2_lut (.A(n1025), .B(o_Rx_Byte_c_3), .Z(n2359)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i2966_2_lut.init = 16'h8888;
    LUT4 mux_743_i3_3_lut (.A(o_Rx_Byte_c_2), .B(o_Rx_Byte_c_4), .C(n2795), 
         .Z(n3632)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_743_i3_3_lut.init = 16'hcaca;
    LUT4 i2306_2_lut_3_lut_4_lut_4_lut (.A(o_Rx_Byte_c_0), .B(n8225), .C(o_Rx_Byte_c_3), 
         .D(n13385), .Z(n8341)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;
    defparam i2306_2_lut_3_lut_4_lut_4_lut.init = 16'hf4f0;
    LUT4 i1_4_lut_4_lut_4_lut (.A(o_Rx_Byte_c_0), .B(n8225), .C(o_Rx_Byte_c_2), 
         .D(o_Rx_Byte_c_4), .Z(n12919)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A ((D)+!B))) */ ;
    defparam i1_4_lut_4_lut_4_lut.init = 16'h00c4;
    LUT4 i1_3_lut_rep_79 (.A(o_Rx_Byte_c_7), .B(o_Rx_DV_c), .C(o_Rx_Byte_c_5), 
         .Z(n13390)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_3_lut_rep_79.init = 16'h4040;
    LUT4 i1746_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1048), .Z(n7769)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i1746_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_2_lut_4_lut (.A(o_Rx_Byte_c_7), .B(o_Rx_DV_c), .C(o_Rx_Byte_c_5), 
         .D(o_Rx_Byte_c_6), .Z(n8225)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h4000;
    LUT4 i1728_3_lut_4_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n1058), .C(o_Rx_Byte_c_3), 
         .D(n13381), .Z(n7751)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1728_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 mux_318_i47_4_lut (.A(n7805), .B(n1089), .C(n13376), .D(n13375), 
         .Z(n2296)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i47_4_lut.init = 16'hc0ca;
    LUT4 mux_318_i48_4_lut (.A(n7807), .B(n1088), .C(n13376), .D(n13375), 
         .Z(n2295)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i48_4_lut.init = 16'hcfca;
    LUT4 i1764_3_lut_4_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n1039), .C(o_Rx_Byte_c_3), 
         .D(n13381), .Z(n7787)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1764_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i1766_3_lut_4_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n1038), .C(o_Rx_Byte_c_3), 
         .D(n13381), .Z(n7789)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1766_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i1748_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1047), .Z(n7771)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;
    defparam i1748_3_lut_4_lut.init = 16'hf707;
    LUT4 mux_318_i45_4_lut (.A(n2364), .B(n1091), .C(n13376), .D(n7970), 
         .Z(n2298)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i45_4_lut.init = 16'hc0ca;
    LUT4 i1720_3_lut_4_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n1064), .C(o_Rx_Byte_c_3), 
         .D(n13381), .Z(n7743)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1720_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i1772_3_lut_4_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n1035), .C(o_Rx_Byte_c_3), 
         .D(n13381), .Z(n7795)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1772_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i1750_3_lut_4_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n1046), .C(o_Rx_Byte_c_3), 
         .D(n13381), .Z(n7773)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1750_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 mux_318_i46_4_lut (.A(n7803), .B(n1090), .C(n13376), .D(n13375), 
         .Z(n2297)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i46_4_lut.init = 16'hcfca;
    LUT4 i2884_2_lut (.A(o_Rx_Byte_c_4), .B(n2795), .Z(n3653)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i2884_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_4_lut (.A(o_Rx_Byte_c_2), .B(o_Rx_Byte_c_0), .C(o_Rx_Byte_c_6), 
         .D(n13390), .Z(n12931)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1_4_lut_4_lut.init = 16'h4000;
    LUT4 i1744_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1049), .Z(n7767)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i1744_3_lut_4_lut.init = 16'hf808;
    LUT4 i1756_3_lut_4_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n1043), .C(o_Rx_Byte_c_3), 
         .D(n13381), .Z(n7779)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1756_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i1710_3_lut_4_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n1070), .C(o_Rx_Byte_c_3), 
         .D(n13381), .Z(n7733)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1710_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 mux_743_i2_3_lut_3_lut (.A(o_Rx_Byte_c_2), .B(n2795), .C(o_Rx_Byte_c_4), 
         .Z(n3663)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_743_i2_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i1770_3_lut_4_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n1036), .C(o_Rx_Byte_c_3), 
         .D(n13381), .Z(n7793)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1770_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i1790_3_lut_4_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n1023), .C(o_Rx_Byte_c_3), 
         .D(n13381), .Z(n7813)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1790_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i1740_3_lut_4_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n1051), .C(o_Rx_Byte_c_3), 
         .D(n13381), .Z(n7763)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1740_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i1736_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1054), .Z(n7759)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;
    defparam i1736_3_lut_4_lut.init = 16'hf707;
    LUT4 i1742_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1050), .Z(n7765)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1742_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i1780_3_lut_4_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n1029), .C(o_Rx_Byte_c_3), 
         .D(n13381), .Z(n7803)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1780_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 mux_318_i39_4_lut (.A(n7793), .B(n1097), .C(n13376), .D(n13375), 
         .Z(n2304)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i39_4_lut.init = 16'hc0ca;
    LUT4 i1726_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1060), .Z(n7749)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i1726_3_lut_4_lut.init = 16'hf808;
    OB o_Rx_DV_pad (.I(o_Rx_DV_c), .O(o_Rx_DV));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(49[13:20])
    OB o_Tx_Serial_pad (.I(GND_net), .O(o_Tx_Serial));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(48[11:22])
    \uart_rx(CLKS_PER_BIT=87)  uart_rx1 (.o_Rx_Byte_c_2(o_Rx_Byte_c_2), .n8225(n8225), 
            .n2795(n2795), .o_Rx_Byte_c_4(o_Rx_Byte_c_4), .n13291(n13291), 
            .n12970(n12970), .n13523(n13523), .osc_clk(osc_clk), .i_Rx_Serial_c(i_Rx_Serial_c), 
            .o_Rx_Byte_c_0(o_Rx_Byte_c_0), .osc_clk_enable_1447(osc_clk_enable_1447), 
            .n3614(n3614), .o_Rx_Byte_c_3(o_Rx_Byte_c_3), .n6(n6), .n12803(n12803), 
            .n13380(n13380), .n3628(n3628), .osc_clk_enable_1457(osc_clk_enable_1457), 
            .n7349(n7349), .n13385(n13385), .n2608(n2608), .n1132(n1132), 
            .n13383(n13383), .n2339(n2339), .n1030(n1030), .n2364(n2364), 
            .n1018(n1018), .n2486(n2486), .n12919(n12919), .n12931(n12931), 
            .n13372(n13372), .n1034(n1034), .n13381(n13381), .n30(n30), 
            .n7970(n7970), .n13376(n13376), .n13375(n13375), .n1052(n1052), 
            .n28(n28), .n1045(n1045), .n2513(n2513), .n1059(n1059), 
            .n29(n29), .GND_net(GND_net), .o_Rx_Byte_c_5(o_Rx_Byte_c_5), 
            .o_Rx_Byte_c_6(o_Rx_Byte_c_6), .o_Rx_Byte_c_7(o_Rx_Byte_c_7), 
            .n9000(n9000), .osc_clk_enable_128(osc_clk_enable_128), .n1128(n1128), 
            .n1067(n1067), .n13384(n13384), .n1062(n1062), .n2530(n2530), 
            .o_Rx_DV_c(o_Rx_DV_c), .n13411(n13411)) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(217[32] 222[2])
    LUT4 i1732_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1056), .Z(n7755)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1732_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i1716_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1066), .Z(n7739)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i1716_3_lut_4_lut.init = 16'hf808;
    OB o_Rx_Byte_pad_5 (.I(o_Rx_Byte_c_5), .O(o_Rx_Byte[5]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[16:25])
    OB o_Rx_Byte_pad_4 (.I(o_Rx_Byte_c_4), .O(o_Rx_Byte[4]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[16:25])
    OB o_Rx_Byte_pad_3 (.I(o_Rx_Byte_c_3), .O(o_Rx_Byte[3]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[16:25])
    OB o_Rx_Byte_pad_2 (.I(o_Rx_Byte_c_2), .O(o_Rx_Byte[2]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[16:25])
    OB o_Rx_Byte_pad_1 (.I(n7349), .O(o_Rx_Byte[1]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[16:25])
    OB o_Rx_Byte_pad_0 (.I(o_Rx_Byte_c_0), .O(o_Rx_Byte[0]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[16:25])
    OB MYLED_pad_7 (.I(GND_net), .O(MYLED[7]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(51[18:23])
    OB MYLED_pad_6 (.I(n7349), .O(MYLED[6]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(51[18:23])
    OB MYLED_pad_5 (.I(MYLED_c_5), .O(MYLED[5]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(51[18:23])
    OB MYLED_pad_4 (.I(MYLED_c_4), .O(MYLED[4]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(51[18:23])
    OB MYLED_pad_3 (.I(MYLED_c_3), .O(MYLED[3]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(51[18:23])
    OB MYLED_pad_2 (.I(MYLED_c_2), .O(MYLED[2]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(51[18:23])
    OB MYLED_pad_1 (.I(MYLED_c_1), .O(MYLED[1]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(51[18:23])
    OB MYLED_pad_0 (.I(MYLED_c_0), .O(MYLED[0]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(51[18:23])
    OB XOut_pad (.I(GND_net), .O(XOut));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(55[9:13])
    OB DiffOut_pad (.I(DiffOut_c), .O(DiffOut));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(57[9:16])
    OB PWMOut_pad (.I(PWMOutP4_c), .O(PWMOut));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(58[9:15])
    OB PWMOutP1_pad (.I(PWMOutP4_c), .O(PWMOutP1));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(59[9:17])
    OB PWMOutP2_pad (.I(PWMOutP4_c), .O(PWMOutP2));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(60[9:17])
    OB PWMOutP3_pad (.I(PWMOutP4_c), .O(PWMOutP3));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(61[9:17])
    OB PWMOutP4_pad (.I(PWMOutP4_c), .O(PWMOutP4));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(62[9:17])
    OB PWMOutN1_pad (.I(PWMOutN4_c), .O(PWMOutN1));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(63[9:17])
    OB PWMOutN2_pad (.I(PWMOutN4_c), .O(PWMOutN2));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(64[9:17])
    OB PWMOutN3_pad (.I(PWMOutN4_c), .O(PWMOutN3));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(65[9:17])
    OB PWMOutN4_pad (.I(PWMOutN4_c), .O(PWMOutN4));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(66[9:17])
    OB sinGen_pad (.I(sinGen_c), .O(sinGen));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(67[9:15])
    OB sin_out_pad (.I(GND_net), .O(sin_out));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(68[9:16])
    OB CIC_out_clkSin_pad (.I(GND_net), .O(CIC_out_clkSin));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(69[9:23])
    IB i_Rx_Serial_pad (.I(i_Rx_Serial), .O(i_Rx_Serial_c));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(47[13:24])
    IB RFIn_pad (.I(RFIn), .O(RFIn_c));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(56[9:13])
    LUT4 mux_318_i40_4_lut (.A(n7795), .B(n1096), .C(n13376), .D(n13375), 
         .Z(n2303)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i40_4_lut.init = 16'hcfca;
    FD1P3AX phase_inc_carrGen_i0_i0 (.D(n2860), .SP(osc_clk_enable_128), 
            .CK(osc_clk), .Q(phase_inc_carrGen[0]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i0.GSR = "ENABLED";
    LUT4 mux_318_i37_4_lut (.A(n7789), .B(n1099), .C(n13376), .D(n13375), 
         .Z(n2306)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i37_4_lut.init = 16'hcfca;
    LUT4 i3496_3_lut (.A(phase_inc_carrGen[37]), .B(n2305), .C(n9000), 
         .Z(n9527)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i3496_3_lut.init = 16'hacac;
    FD1S3AX phase_inc_carrGen1_i49 (.D(phase_inc_carrGen[49]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[49]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i49.GSR = "ENABLED";
    LUT4 mux_318_i43_4_lut (.A(n7799), .B(n1093), .C(n13376), .D(n13375), 
         .Z(n2300)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i43_4_lut.init = 16'hc0ca;
    FD1S3AX phase_inc_carrGen1_i50 (.D(phase_inc_carrGen[50]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[50]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i50.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i51 (.D(phase_inc_carrGen[51]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[51]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i51.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i52 (.D(phase_inc_carrGen[52]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[52]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i52.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i53 (.D(phase_inc_carrGen[53]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[53]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i53.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i54 (.D(phase_inc_carrGen[54]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[54]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i54.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i55 (.D(phase_inc_carrGen[55]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[55]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i55.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i56 (.D(phase_inc_carrGen[56]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[56]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i56.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i57 (.D(phase_inc_carrGen[57]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[57]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i57.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i58 (.D(phase_inc_carrGen[58]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[58]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i58.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i59 (.D(phase_inc_carrGen[59]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[59]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i59.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i60 (.D(phase_inc_carrGen[60]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[60]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i60.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i61 (.D(phase_inc_carrGen[61]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[61]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i61.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i62 (.D(phase_inc_carrGen[62]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[62]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i62.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i63 (.D(phase_inc_carrGen[63]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[63]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen1_i63.GSR = "ENABLED";
    FD1P3AX CICGain__i2 (.D(n7349), .SP(osc_clk_enable_1394), .CK(osc_clk), 
            .Q(CICGain[1]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam CICGain__i2.GSR = "ENABLED";
    LUT4 i1718_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1065), .Z(n7741)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;
    defparam i1718_3_lut_4_lut.init = 16'hf707;
    FD1P3AX phase_inc_carrGen_i0_i1 (.D(n2859), .SP(osc_clk_enable_1397), 
            .CK(osc_clk), .Q(phase_inc_carrGen[1]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i1.GSR = "ENABLED";
    LUT4 i1712_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1069), .Z(n7735)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i1712_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_318_i38_4_lut (.A(n7791), .B(n1098), .C(n13376), .D(n13375), 
         .Z(n2305)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i38_4_lut.init = 16'hc0ca;
    CCU2D sub_42_add_2_63 (.A0(phase_inc_carrGen[62]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[63]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11340), .S0(n1073), .S1(n1072));
    defparam sub_42_add_2_63.INIT0 = 16'h5555;
    defparam sub_42_add_2_63.INIT1 = 16'h5555;
    defparam sub_42_add_2_63.INJECT1_0 = "NO";
    defparam sub_42_add_2_63.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_61 (.A0(phase_inc_carrGen[60]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[61]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11339), .COUT(n11340), .S0(n1075), .S1(n1074));
    defparam sub_42_add_2_61.INIT0 = 16'h5555;
    defparam sub_42_add_2_61.INIT1 = 16'h5555;
    defparam sub_42_add_2_61.INJECT1_0 = "NO";
    defparam sub_42_add_2_61.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_59 (.A0(phase_inc_carrGen[58]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[59]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11338), .COUT(n11339), .S0(n1077), .S1(n1076));
    defparam sub_42_add_2_59.INIT0 = 16'h5555;
    defparam sub_42_add_2_59.INIT1 = 16'h5555;
    defparam sub_42_add_2_59.INJECT1_0 = "NO";
    defparam sub_42_add_2_59.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_57 (.A0(phase_inc_carrGen[56]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[57]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11337), .COUT(n11338), .S0(n1079), .S1(n1078));
    defparam sub_42_add_2_57.INIT0 = 16'h5555;
    defparam sub_42_add_2_57.INIT1 = 16'h5555;
    defparam sub_42_add_2_57.INJECT1_0 = "NO";
    defparam sub_42_add_2_57.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_55 (.A0(phase_inc_carrGen[54]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[55]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11336), .COUT(n11337), .S0(n1081), .S1(n1080));
    defparam sub_42_add_2_55.INIT0 = 16'h5555;
    defparam sub_42_add_2_55.INIT1 = 16'h5555;
    defparam sub_42_add_2_55.INJECT1_0 = "NO";
    defparam sub_42_add_2_55.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_53 (.A0(phase_inc_carrGen[52]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[53]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11335), .COUT(n11336), .S0(n1083), .S1(n1082));
    defparam sub_42_add_2_53.INIT0 = 16'h5555;
    defparam sub_42_add_2_53.INIT1 = 16'h5555;
    defparam sub_42_add_2_53.INJECT1_0 = "NO";
    defparam sub_42_add_2_53.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_51 (.A0(phase_inc_carrGen[50]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[51]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11334), .COUT(n11335), .S0(n1085), .S1(n1084));
    defparam sub_42_add_2_51.INIT0 = 16'h5aaa;
    defparam sub_42_add_2_51.INIT1 = 16'h5aaa;
    defparam sub_42_add_2_51.INJECT1_0 = "NO";
    defparam sub_42_add_2_51.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_49 (.A0(phase_inc_carrGen[48]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[49]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11333), .COUT(n11334), .S0(n1087), .S1(n1086));
    defparam sub_42_add_2_49.INIT0 = 16'h5555;
    defparam sub_42_add_2_49.INIT1 = 16'h5555;
    defparam sub_42_add_2_49.INJECT1_0 = "NO";
    defparam sub_42_add_2_49.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_47 (.A0(phase_inc_carrGen[46]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[47]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11332), .COUT(n11333), .S0(n1089), .S1(n1088));
    defparam sub_42_add_2_47.INIT0 = 16'h5555;
    defparam sub_42_add_2_47.INIT1 = 16'h5aaa;
    defparam sub_42_add_2_47.INJECT1_0 = "NO";
    defparam sub_42_add_2_47.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_45 (.A0(phase_inc_carrGen[44]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[45]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11331), .COUT(n11332), .S0(n1091), .S1(n1090));
    defparam sub_42_add_2_45.INIT0 = 16'h5555;
    defparam sub_42_add_2_45.INIT1 = 16'h5aaa;
    defparam sub_42_add_2_45.INJECT1_0 = "NO";
    defparam sub_42_add_2_45.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_43 (.A0(phase_inc_carrGen[42]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[43]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11330), .COUT(n11331), .S0(n1093), .S1(n1092));
    defparam sub_42_add_2_43.INIT0 = 16'h5555;
    defparam sub_42_add_2_43.INIT1 = 16'h5555;
    defparam sub_42_add_2_43.INJECT1_0 = "NO";
    defparam sub_42_add_2_43.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_41 (.A0(phase_inc_carrGen[40]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[41]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11329), .COUT(n11330), .S0(n1095), .S1(n1094));
    defparam sub_42_add_2_41.INIT0 = 16'h5555;
    defparam sub_42_add_2_41.INIT1 = 16'h5aaa;
    defparam sub_42_add_2_41.INJECT1_0 = "NO";
    defparam sub_42_add_2_41.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_39 (.A0(phase_inc_carrGen[38]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[39]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11328), .COUT(n11329), .S0(n1097), .S1(n1096));
    defparam sub_42_add_2_39.INIT0 = 16'h5555;
    defparam sub_42_add_2_39.INIT1 = 16'h5555;
    defparam sub_42_add_2_39.INJECT1_0 = "NO";
    defparam sub_42_add_2_39.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_37 (.A0(phase_inc_carrGen[36]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[37]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11327), .COUT(n11328), .S0(n1099), .S1(n1098));
    defparam sub_42_add_2_37.INIT0 = 16'h5555;
    defparam sub_42_add_2_37.INIT1 = 16'h5aaa;
    defparam sub_42_add_2_37.INJECT1_0 = "NO";
    defparam sub_42_add_2_37.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_35 (.A0(phase_inc_carrGen[34]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[35]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11326), .COUT(n11327), .S0(n1101), .S1(n1100));
    defparam sub_42_add_2_35.INIT0 = 16'h5555;
    defparam sub_42_add_2_35.INIT1 = 16'h5aaa;
    defparam sub_42_add_2_35.INJECT1_0 = "NO";
    defparam sub_42_add_2_35.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_33 (.A0(phase_inc_carrGen[32]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[33]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11325), .COUT(n11326), .S0(n1103), .S1(n1102));
    defparam sub_42_add_2_33.INIT0 = 16'h5aaa;
    defparam sub_42_add_2_33.INIT1 = 16'h5555;
    defparam sub_42_add_2_33.INJECT1_0 = "NO";
    defparam sub_42_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_31 (.A0(phase_inc_carrGen[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11324), .COUT(n11325), .S0(n1105), .S1(n1104));
    defparam sub_42_add_2_31.INIT0 = 16'h5555;
    defparam sub_42_add_2_31.INIT1 = 16'h5aaa;
    defparam sub_42_add_2_31.INJECT1_0 = "NO";
    defparam sub_42_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_29 (.A0(phase_inc_carrGen[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11323), .COUT(n11324), .S0(n1107), .S1(n1106));
    defparam sub_42_add_2_29.INIT0 = 16'h5555;
    defparam sub_42_add_2_29.INIT1 = 16'h5555;
    defparam sub_42_add_2_29.INJECT1_0 = "NO";
    defparam sub_42_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_27 (.A0(phase_inc_carrGen[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11322), .COUT(n11323), .S0(n1109), .S1(n1108));
    defparam sub_42_add_2_27.INIT0 = 16'h5555;
    defparam sub_42_add_2_27.INIT1 = 16'h5555;
    defparam sub_42_add_2_27.INJECT1_0 = "NO";
    defparam sub_42_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_25 (.A0(phase_inc_carrGen[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11321), .COUT(n11322), .S0(n1111), .S1(n1110));
    defparam sub_42_add_2_25.INIT0 = 16'h5555;
    defparam sub_42_add_2_25.INIT1 = 16'h5555;
    defparam sub_42_add_2_25.INJECT1_0 = "NO";
    defparam sub_42_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_23 (.A0(phase_inc_carrGen[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11320), .COUT(n11321), .S0(n1113), .S1(n1112));
    defparam sub_42_add_2_23.INIT0 = 16'h5555;
    defparam sub_42_add_2_23.INIT1 = 16'h5aaa;
    defparam sub_42_add_2_23.INJECT1_0 = "NO";
    defparam sub_42_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_21 (.A0(phase_inc_carrGen[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11319), .COUT(n11320), .S0(n1115), .S1(n1114));
    defparam sub_42_add_2_21.INIT0 = 16'h5aaa;
    defparam sub_42_add_2_21.INIT1 = 16'h5aaa;
    defparam sub_42_add_2_21.INJECT1_0 = "NO";
    defparam sub_42_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_19 (.A0(phase_inc_carrGen[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11318), .COUT(n11319), .S0(n1117), .S1(n1116));
    defparam sub_42_add_2_19.INIT0 = 16'h5555;
    defparam sub_42_add_2_19.INIT1 = 16'h5aaa;
    defparam sub_42_add_2_19.INJECT1_0 = "NO";
    defparam sub_42_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_17 (.A0(phase_inc_carrGen[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11317), .COUT(n11318), .S0(n1119), .S1(n1118));
    defparam sub_42_add_2_17.INIT0 = 16'h5555;
    defparam sub_42_add_2_17.INIT1 = 16'h5aaa;
    defparam sub_42_add_2_17.INJECT1_0 = "NO";
    defparam sub_42_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_15 (.A0(phase_inc_carrGen[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11316), .COUT(n11317), .S0(n1121), .S1(n1120));
    defparam sub_42_add_2_15.INIT0 = 16'h5aaa;
    defparam sub_42_add_2_15.INIT1 = 16'h5555;
    defparam sub_42_add_2_15.INJECT1_0 = "NO";
    defparam sub_42_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_13 (.A0(phase_inc_carrGen[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11315), .COUT(n11316), .S0(n1123), .S1(n1122));
    defparam sub_42_add_2_13.INIT0 = 16'h5aaa;
    defparam sub_42_add_2_13.INIT1 = 16'h5555;
    defparam sub_42_add_2_13.INJECT1_0 = "NO";
    defparam sub_42_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_11 (.A0(phase_inc_carrGen[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11314), .COUT(n11315), .S0(n1125), .S1(n1124));
    defparam sub_42_add_2_11.INIT0 = 16'h5aaa;
    defparam sub_42_add_2_11.INIT1 = 16'h5555;
    defparam sub_42_add_2_11.INJECT1_0 = "NO";
    defparam sub_42_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_9 (.A0(phase_inc_carrGen[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11313), .COUT(n11314), .S0(n1127), .S1(n1126));
    defparam sub_42_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_42_add_2_9.INIT1 = 16'h5aaa;
    defparam sub_42_add_2_9.INJECT1_0 = "NO";
    defparam sub_42_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_7 (.A0(phase_inc_carrGen[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11312), .COUT(n11313), .S0(n1129), .S1(n1128));
    defparam sub_42_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_42_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_42_add_2_7.INJECT1_0 = "NO";
    defparam sub_42_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_5 (.A0(phase_inc_carrGen[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11311), .COUT(n11312), .S0(n1131), .S1(n1130));
    defparam sub_42_add_2_5.INIT0 = 16'h5555;
    defparam sub_42_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_42_add_2_5.INJECT1_0 = "NO";
    defparam sub_42_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_3 (.A0(phase_inc_carrGen[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11310), .COUT(n11311), .S0(n1133), .S1(n1132));
    defparam sub_42_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_42_add_2_3.INIT1 = 16'h5555;
    defparam sub_42_add_2_3.INJECT1_0 = "NO";
    defparam sub_42_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_42_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(phase_inc_carrGen[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n11310), .S1(n1134));
    defparam sub_42_add_2_1.INIT0 = 16'hF000;
    defparam sub_42_add_2_1.INIT1 = 16'h5555;
    defparam sub_42_add_2_1.INJECT1_0 = "NO";
    defparam sub_42_add_2_1.INJECT1_1 = "NO";
    CCU2D add_745_65 (.A0(n3614), .B0(n9000), .C0(n8014), .D0(phase_inc_carrGen[62]), 
          .A1(n3614), .B1(n9000), .C1(n8016), .D1(phase_inc_carrGen[63]), 
          .CIN(n11302), .S0(n2798), .S1(n2797));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_65.INIT0 = 16'h74b8;
    defparam add_745_65.INIT1 = 16'h74b8;
    defparam add_745_65.INJECT1_0 = "NO";
    defparam add_745_65.INJECT1_1 = "NO";
    CCU2D add_745_63 (.A0(n3614), .B0(n9000), .C0(n2282), .D0(phase_inc_carrGen[60]), 
          .A1(n3614), .B1(n9000), .C1(n8012), .D1(phase_inc_carrGen[61]), 
          .CIN(n11301), .COUT(n11302), .S0(n2800), .S1(n2799));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_63.INIT0 = 16'h74b8;
    defparam add_745_63.INIT1 = 16'h74b8;
    defparam add_745_63.INJECT1_0 = "NO";
    defparam add_745_63.INJECT1_1 = "NO";
    CCU2D add_745_61 (.A0(n3614), .B0(n9000), .C0(n2284), .D0(phase_inc_carrGen[58]), 
          .A1(n3614), .B1(n9000), .C1(n2283), .D1(phase_inc_carrGen[59]), 
          .CIN(n11300), .COUT(n11301), .S0(n2802), .S1(n2801));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_61.INIT0 = 16'h74b8;
    defparam add_745_61.INIT1 = 16'h74b8;
    defparam add_745_61.INJECT1_0 = "NO";
    defparam add_745_61.INJECT1_1 = "NO";
    CCU2D add_745_59 (.A0(n3614), .B0(n9000), .C0(n2286), .D0(phase_inc_carrGen[56]), 
          .A1(n3614), .B1(n9000), .C1(n2285), .D1(phase_inc_carrGen[57]), 
          .CIN(n11299), .COUT(n11300), .S0(n2804), .S1(n2803));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_59.INIT0 = 16'h74b8;
    defparam add_745_59.INIT1 = 16'h74b8;
    defparam add_745_59.INJECT1_0 = "NO";
    defparam add_745_59.INJECT1_1 = "NO";
    CCU2D add_745_57 (.A0(n3614), .B0(n9000), .C0(n2288), .D0(phase_inc_carrGen[54]), 
          .A1(n3614), .B1(n9000), .C1(n2287), .D1(phase_inc_carrGen[55]), 
          .CIN(n11298), .COUT(n11299), .S0(n2806), .S1(n2805));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_57.INIT0 = 16'h74b8;
    defparam add_745_57.INIT1 = 16'h74b8;
    defparam add_745_57.INJECT1_0 = "NO";
    defparam add_745_57.INJECT1_1 = "NO";
    CCU2D add_745_55 (.A0(n3614), .B0(n9000), .C0(n8010), .D0(phase_inc_carrGen[52]), 
          .A1(n3614), .B1(n9000), .C1(n2289), .D1(phase_inc_carrGen[53]), 
          .CIN(n11297), .COUT(n11298), .S0(n2808), .S1(n2807));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_55.INIT0 = 16'h74b8;
    defparam add_745_55.INIT1 = 16'h74b8;
    defparam add_745_55.INJECT1_0 = "NO";
    defparam add_745_55.INJECT1_1 = "NO";
    CCU2D add_745_53 (.A0(n3628), .B0(n9000), .C0(n2292), .D0(phase_inc_carrGen[50]), 
          .A1(n3614), .B1(n9000), .C1(n2291), .D1(phase_inc_carrGen[51]), 
          .CIN(n11296), .COUT(n11297), .S0(n2810), .S1(n2809));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_53.INIT0 = 16'h74b8;
    defparam add_745_53.INIT1 = 16'h74b8;
    defparam add_745_53.INJECT1_0 = "NO";
    defparam add_745_53.INJECT1_1 = "NO";
    CCU2D add_745_51 (.A0(n3628), .B0(n9000), .C0(n2294), .D0(phase_inc_carrGen[48]), 
          .A1(n3628), .B1(n9000), .C1(n2293), .D1(phase_inc_carrGen[49]), 
          .CIN(n11295), .COUT(n11296), .S0(n2812), .S1(n2811));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_51.INIT0 = 16'h74b8;
    defparam add_745_51.INIT1 = 16'h74b8;
    defparam add_745_51.INJECT1_0 = "NO";
    defparam add_745_51.INJECT1_1 = "NO";
    CCU2D add_745_49 (.A0(n3632), .B0(n9000), .C0(n2296), .D0(phase_inc_carrGen[46]), 
          .A1(n3632), .B1(n9000), .C1(n2295), .D1(phase_inc_carrGen[47]), 
          .CIN(n11294), .COUT(n11295), .S0(n2814), .S1(n2813));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_49.INIT0 = 16'hb874;
    defparam add_745_49.INIT1 = 16'hb874;
    defparam add_745_49.INJECT1_0 = "NO";
    defparam add_745_49.INJECT1_1 = "NO";
    CCU2D add_745_47 (.A0(n3632), .B0(n9000), .C0(n2298), .D0(phase_inc_carrGen[44]), 
          .A1(n3614), .B1(n9000), .C1(n2297), .D1(phase_inc_carrGen[45]), 
          .CIN(n11293), .COUT(n11294), .S0(n2816), .S1(n2815));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_47.INIT0 = 16'h74b8;
    defparam add_745_47.INIT1 = 16'h74b8;
    defparam add_745_47.INJECT1_0 = "NO";
    defparam add_745_47.INJECT1_1 = "NO";
    CCU2D add_745_45 (.A0(n3653), .B0(n9000), .C0(n2300), .D0(phase_inc_carrGen[42]), 
          .A1(n3653), .B1(n9000), .C1(n2299), .D1(phase_inc_carrGen[43]), 
          .CIN(n11292), .COUT(n11293), .S0(n2818), .S1(n2817));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_45.INIT0 = 16'h74b8;
    defparam add_745_45.INIT1 = 16'hb874;
    defparam add_745_45.INJECT1_0 = "NO";
    defparam add_745_45.INJECT1_1 = "NO";
    CCU2D add_745_43 (.A0(n3628), .B0(n9000), .C0(n2302), .D0(phase_inc_carrGen[40]), 
          .A1(n3653), .B1(n9000), .C1(n8008), .D1(phase_inc_carrGen[41]), 
          .CIN(n11291), .COUT(n11292), .S0(n2820), .S1(n2819));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_43.INIT0 = 16'h74b8;
    defparam add_745_43.INIT1 = 16'hb874;
    defparam add_745_43.INJECT1_0 = "NO";
    defparam add_745_43.INJECT1_1 = "NO";
    CCU2D add_745_41 (.A0(n3614), .B0(n9000), .C0(n2304), .D0(phase_inc_carrGen[38]), 
          .A1(n3614), .B1(n9000), .C1(n2303), .D1(phase_inc_carrGen[39]), 
          .CIN(n11290), .COUT(n11291), .S0(n2822), .S1(n2821));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_41.INIT0 = 16'h74b8;
    defparam add_745_41.INIT1 = 16'h74b8;
    defparam add_745_41.INJECT1_0 = "NO";
    defparam add_745_41.INJECT1_1 = "NO";
    CCU2D add_745_39 (.A0(n3632), .B0(n9000), .C0(n2306), .D0(phase_inc_carrGen[36]), 
          .A1(n9527), .B1(n2795), .C1(n9000), .D1(o_Rx_Byte_c_4), .CIN(n11289), 
          .COUT(n11290), .S0(n2824), .S1(n2823));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_39.INIT0 = 16'h74b8;
    defparam add_745_39.INIT1 = 16'h5a9a;
    defparam add_745_39.INJECT1_0 = "NO";
    defparam add_745_39.INJECT1_1 = "NO";
    CCU2D add_745_37 (.A0(n3632), .B0(n9000), .C0(n2308), .D0(phase_inc_carrGen[34]), 
          .A1(n3614), .B1(n9000), .C1(n2307), .D1(phase_inc_carrGen[35]), 
          .CIN(n11288), .COUT(n11289), .S0(n2826), .S1(n2825));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_37.INIT0 = 16'h74b8;
    defparam add_745_37.INIT1 = 16'h74b8;
    defparam add_745_37.INJECT1_0 = "NO";
    defparam add_745_37.INJECT1_1 = "NO";
    CCU2D add_745_35 (.A0(n3628), .B0(n9000), .C0(n2310), .D0(phase_inc_carrGen[32]), 
          .A1(n9535), .B1(n2795), .C1(n9000), .D1(o_Rx_Byte_c_4), .CIN(n11287), 
          .COUT(n11288), .S0(n2828), .S1(n2827));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_35.INIT0 = 16'h74b8;
    defparam add_745_35.INIT1 = 16'h5a9a;
    defparam add_745_35.INJECT1_0 = "NO";
    defparam add_745_35.INJECT1_1 = "NO";
    CCU2D add_745_33 (.A0(n3628), .B0(n9000), .C0(n2312), .D0(phase_inc_carrGen[30]), 
          .A1(n3663), .B1(n9000), .C1(n2311), .D1(phase_inc_carrGen[31]), 
          .CIN(n11286), .COUT(n11287), .S0(n2830), .S1(n2829));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_33.INIT0 = 16'h74b8;
    defparam add_745_33.INIT1 = 16'h74b8;
    defparam add_745_33.INJECT1_0 = "NO";
    defparam add_745_33.INJECT1_1 = "NO";
    CCU2D add_745_31 (.A0(n3653), .B0(n9000), .C0(n2314), .D0(phase_inc_carrGen[28]), 
          .A1(n3653), .B1(n9000), .C1(n2313), .D1(phase_inc_carrGen[29]), 
          .CIN(n11285), .COUT(n11286), .S0(n2832), .S1(n2831));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_31.INIT0 = 16'hb874;
    defparam add_745_31.INIT1 = 16'h74b8;
    defparam add_745_31.INJECT1_0 = "NO";
    defparam add_745_31.INJECT1_1 = "NO";
    CCU2D add_745_29 (.A0(n3614), .B0(n9000), .C0(n2316), .D0(phase_inc_carrGen[26]), 
          .A1(n9547), .B1(n2795), .C1(n9000), .D1(o_Rx_Byte_c_4), .CIN(n11284), 
          .COUT(n11285), .S0(n2834), .S1(n2833));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_29.INIT0 = 16'h74b8;
    defparam add_745_29.INIT1 = 16'h5a9a;
    defparam add_745_29.INJECT1_0 = "NO";
    defparam add_745_29.INJECT1_1 = "NO";
    CCU2D add_745_27 (.A0(n3614), .B0(n9000), .C0(n2318), .D0(phase_inc_carrGen[24]), 
          .A1(n3614), .B1(n9000), .C1(n2317), .D1(phase_inc_carrGen[25]), 
          .CIN(n11283), .COUT(n11284), .S0(n2836), .S1(n2835));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_27.INIT0 = 16'h74b8;
    defparam add_745_27.INIT1 = 16'h74b8;
    defparam add_745_27.INJECT1_0 = "NO";
    defparam add_745_27.INJECT1_1 = "NO";
    CCU2D add_745_25 (.A0(n3632), .B0(n9000), .C0(n2320), .D0(phase_inc_carrGen[22]), 
          .A1(n3653), .B1(n9000), .C1(n2319), .D1(phase_inc_carrGen[23]), 
          .CIN(n11282), .COUT(n11283), .S0(n2838), .S1(n2837));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_25.INIT0 = 16'h74b8;
    defparam add_745_25.INIT1 = 16'h74b8;
    defparam add_745_25.INJECT1_0 = "NO";
    defparam add_745_25.INJECT1_1 = "NO";
    CCU2D add_745_23 (.A0(n3614), .B0(n9000), .C0(n2322), .D0(phase_inc_carrGen[20]), 
          .A1(n3628), .B1(n9000), .C1(n2321), .D1(phase_inc_carrGen[21]), 
          .CIN(n11281), .COUT(n11282), .S0(n2840), .S1(n2839));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_23.INIT0 = 16'h74b8;
    defparam add_745_23.INIT1 = 16'h74b8;
    defparam add_745_23.INJECT1_0 = "NO";
    defparam add_745_23.INJECT1_1 = "NO";
    CCU2D add_745_21 (.A0(n3653), .B0(n9000), .C0(n2324), .D0(phase_inc_carrGen[18]), 
          .A1(n9563), .B1(n2795), .C1(n9000), .D1(o_Rx_Byte_c_4), .CIN(n11280), 
          .COUT(n11281), .S0(n2842), .S1(n2841));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_21.INIT0 = 16'h74b8;
    defparam add_745_21.INIT1 = 16'h5a9a;
    defparam add_745_21.INJECT1_0 = "NO";
    defparam add_745_21.INJECT1_1 = "NO";
    CCU2D add_745_19 (.A0(n3663), .B0(n9000), .C0(n2326), .D0(phase_inc_carrGen[16]), 
          .A1(n3632), .B1(n9000), .C1(n8004), .D1(phase_inc_carrGen[17]), 
          .CIN(n11279), .COUT(n11280), .S0(n2844), .S1(n2843));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_19.INIT0 = 16'h74b8;
    defparam add_745_19.INIT1 = 16'hb874;
    defparam add_745_19.INJECT1_0 = "NO";
    defparam add_745_19.INJECT1_1 = "NO";
    CCU2D add_745_17 (.A0(n3632), .B0(n9000), .C0(n2328), .D0(phase_inc_carrGen[14]), 
          .A1(n9571), .B1(n2795), .C1(n9000), .D1(o_Rx_Byte_c_4), .CIN(n11278), 
          .COUT(n11279), .S0(n2846), .S1(n2845));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_17.INIT0 = 16'h74b8;
    defparam add_745_17.INIT1 = 16'h5a9a;
    defparam add_745_17.INJECT1_0 = "NO";
    defparam add_745_17.INJECT1_1 = "NO";
    CCU2D add_745_15 (.A0(n3632), .B0(n9000), .C0(n2330), .D0(phase_inc_carrGen[12]), 
          .A1(n3663), .B1(n9000), .C1(n8002), .D1(phase_inc_carrGen[13]), 
          .CIN(n11277), .COUT(n11278), .S0(n2848), .S1(n2847));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_15.INIT0 = 16'h74b8;
    defparam add_745_15.INIT1 = 16'h74b8;
    defparam add_745_15.INJECT1_0 = "NO";
    defparam add_745_15.INJECT1_1 = "NO";
    CCU2D add_745_13 (.A0(n3663), .B0(n9000), .C0(n2332), .D0(phase_inc_carrGen[10]), 
          .A1(n3614), .B1(n9000), .C1(n2331), .D1(phase_inc_carrGen[11]), 
          .CIN(n11276), .COUT(n11277), .S0(n2850), .S1(n2849));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_13.INIT0 = 16'h74b8;
    defparam add_745_13.INIT1 = 16'h74b8;
    defparam add_745_13.INJECT1_0 = "NO";
    defparam add_745_13.INJECT1_1 = "NO";
    CCU2D add_745_11 (.A0(n3653), .B0(n9000), .C0(n2334), .D0(phase_inc_carrGen[8]), 
          .A1(n3653), .B1(n9000), .C1(n2333), .D1(phase_inc_carrGen[9]), 
          .CIN(n11275), .COUT(n11276), .S0(n2852), .S1(n2851));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_11.INIT0 = 16'hb874;
    defparam add_745_11.INIT1 = 16'h74b8;
    defparam add_745_11.INJECT1_0 = "NO";
    defparam add_745_11.INJECT1_1 = "NO";
    CCU2D add_745_9 (.A0(n9589), .B0(n2795), .C0(n9000), .D0(o_Rx_Byte_c_4), 
          .A1(n3653), .B1(n9000), .C1(n13411), .D1(phase_inc_carrGen[7]), 
          .CIN(n11274), .COUT(n11275), .S0(n2854), .S1(n2853));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_9.INIT0 = 16'h5a9a;
    defparam add_745_9.INIT1 = 16'h74b8;
    defparam add_745_9.INJECT1_0 = "NO";
    defparam add_745_9.INJECT1_1 = "NO";
    CCU2D add_745_7 (.A0(n9593), .B0(n2795), .C0(n9000), .D0(o_Rx_Byte_c_4), 
          .A1(n9591), .B1(n2795), .C1(n9000), .D1(o_Rx_Byte_c_4), .CIN(n11273), 
          .COUT(n11274), .S0(n2856), .S1(n2855));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_7.INIT0 = 16'h5a9a;
    defparam add_745_7.INIT1 = 16'h5a9a;
    defparam add_745_7.INJECT1_0 = "NO";
    defparam add_745_7.INJECT1_1 = "NO";
    CCU2D add_745_5 (.A0(n3632), .B0(n9000), .C0(n2340), .D0(phase_inc_carrGen[2]), 
          .A1(n3632), .B1(n9000), .C1(n2339), .D1(phase_inc_carrGen[3]), 
          .CIN(n11272), .COUT(n11273), .S0(n2858), .S1(n2857));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_5.INIT0 = 16'hb874;
    defparam add_745_5.INIT1 = 16'hb874;
    defparam add_745_5.INJECT1_0 = "NO";
    defparam add_745_5.INJECT1_1 = "NO";
    CCU2D add_745_3 (.A0(n3653), .B0(n9000), .C0(n2608), .D0(phase_inc_carrGen[0]), 
          .A1(n3663), .B1(n9000), .C1(n2341), .D1(phase_inc_carrGen[1]), 
          .CIN(n11271), .COUT(n11272), .S0(n2860), .S1(n2859));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_3.INIT0 = 16'h74b8;
    defparam add_745_3.INIT1 = 16'h74b8;
    defparam add_745_3.INJECT1_0 = "NO";
    defparam add_745_3.INJECT1_1 = "NO";
    CCU2D add_745_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n3614), .B1(n9000), .C1(GND_net), .D1(GND_net), .COUT(n11271));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam add_745_1.INIT0 = 16'hF000;
    defparam add_745_1.INIT1 = 16'h7777;
    defparam add_745_1.INJECT1_0 = "NO";
    defparam add_745_1.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_61 (.A0(phase_inc_carrGen[63]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11129), .S0(n1011));
    defparam sub_41_add_2_61.INIT0 = 16'h5555;
    defparam sub_41_add_2_61.INIT1 = 16'h0000;
    defparam sub_41_add_2_61.INJECT1_0 = "NO";
    defparam sub_41_add_2_61.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_59 (.A0(phase_inc_carrGen[61]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[62]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11128), .COUT(n11129), .S0(n1013), .S1(n1012));
    defparam sub_41_add_2_59.INIT0 = 16'h5555;
    defparam sub_41_add_2_59.INIT1 = 16'h5555;
    defparam sub_41_add_2_59.INJECT1_0 = "NO";
    defparam sub_41_add_2_59.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_57 (.A0(phase_inc_carrGen[59]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[60]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11127), .COUT(n11128), .S0(n1015), .S1(n1014));
    defparam sub_41_add_2_57.INIT0 = 16'h5555;
    defparam sub_41_add_2_57.INIT1 = 16'h5555;
    defparam sub_41_add_2_57.INJECT1_0 = "NO";
    defparam sub_41_add_2_57.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_55 (.A0(phase_inc_carrGen[57]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[58]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11126), .COUT(n11127), .S0(n1017), .S1(n1016));
    defparam sub_41_add_2_55.INIT0 = 16'h5555;
    defparam sub_41_add_2_55.INIT1 = 16'h5555;
    defparam sub_41_add_2_55.INJECT1_0 = "NO";
    defparam sub_41_add_2_55.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_53 (.A0(phase_inc_carrGen[55]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[56]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11125), .COUT(n11126), .S0(n1019), .S1(n1018));
    defparam sub_41_add_2_53.INIT0 = 16'h5555;
    defparam sub_41_add_2_53.INIT1 = 16'h5555;
    defparam sub_41_add_2_53.INJECT1_0 = "NO";
    defparam sub_41_add_2_53.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_51 (.A0(phase_inc_carrGen[53]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[54]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11124), .COUT(n11125), .S0(n1021), .S1(n1020));
    defparam sub_41_add_2_51.INIT0 = 16'h5555;
    defparam sub_41_add_2_51.INIT1 = 16'h5555;
    defparam sub_41_add_2_51.INJECT1_0 = "NO";
    defparam sub_41_add_2_51.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_49 (.A0(phase_inc_carrGen[51]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[52]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11123), .COUT(n11124), .S0(n1023), .S1(n1022));
    defparam sub_41_add_2_49.INIT0 = 16'h5555;
    defparam sub_41_add_2_49.INIT1 = 16'h5555;
    defparam sub_41_add_2_49.INJECT1_0 = "NO";
    defparam sub_41_add_2_49.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_47 (.A0(phase_inc_carrGen[49]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[50]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11122), .COUT(n11123), .S0(n1025), .S1(n1024));
    defparam sub_41_add_2_47.INIT0 = 16'h5aaa;
    defparam sub_41_add_2_47.INIT1 = 16'h5aaa;
    defparam sub_41_add_2_47.INJECT1_0 = "NO";
    defparam sub_41_add_2_47.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_45 (.A0(phase_inc_carrGen[47]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[48]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11121), .COUT(n11122), .S0(n1027), .S1(n1026));
    defparam sub_41_add_2_45.INIT0 = 16'h5555;
    defparam sub_41_add_2_45.INIT1 = 16'h5aaa;
    defparam sub_41_add_2_45.INJECT1_0 = "NO";
    defparam sub_41_add_2_45.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_43 (.A0(phase_inc_carrGen[45]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[46]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11120), .COUT(n11121), .S0(n1029), .S1(n1028));
    defparam sub_41_add_2_43.INIT0 = 16'h5555;
    defparam sub_41_add_2_43.INIT1 = 16'h5555;
    defparam sub_41_add_2_43.INJECT1_0 = "NO";
    defparam sub_41_add_2_43.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_41 (.A0(phase_inc_carrGen[43]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[44]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11119), .COUT(n11120), .S0(n1031), .S1(n1030));
    defparam sub_41_add_2_41.INIT0 = 16'h5aaa;
    defparam sub_41_add_2_41.INIT1 = 16'h5aaa;
    defparam sub_41_add_2_41.INJECT1_0 = "NO";
    defparam sub_41_add_2_41.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_39 (.A0(phase_inc_carrGen[41]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[42]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11118), .COUT(n11119), .S0(n1033), .S1(n1032));
    defparam sub_41_add_2_39.INIT0 = 16'h5aaa;
    defparam sub_41_add_2_39.INIT1 = 16'h5555;
    defparam sub_41_add_2_39.INJECT1_0 = "NO";
    defparam sub_41_add_2_39.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_37 (.A0(phase_inc_carrGen[39]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[40]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11117), .COUT(n11118), .S0(n1035), .S1(n1034));
    defparam sub_41_add_2_37.INIT0 = 16'h5555;
    defparam sub_41_add_2_37.INIT1 = 16'h5aaa;
    defparam sub_41_add_2_37.INJECT1_0 = "NO";
    defparam sub_41_add_2_37.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_35 (.A0(phase_inc_carrGen[37]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[38]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11116), .COUT(n11117), .S0(n1037), .S1(n1036));
    defparam sub_41_add_2_35.INIT0 = 16'h5aaa;
    defparam sub_41_add_2_35.INIT1 = 16'h5555;
    defparam sub_41_add_2_35.INJECT1_0 = "NO";
    defparam sub_41_add_2_35.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_33 (.A0(phase_inc_carrGen[35]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[36]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11115), .COUT(n11116), .S0(n1039), .S1(n1038));
    defparam sub_41_add_2_33.INIT0 = 16'h5555;
    defparam sub_41_add_2_33.INIT1 = 16'h5aaa;
    defparam sub_41_add_2_33.INJECT1_0 = "NO";
    defparam sub_41_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_31 (.A0(phase_inc_carrGen[33]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[34]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11114), .COUT(n11115), .S0(n1041), .S1(n1040));
    defparam sub_41_add_2_31.INIT0 = 16'h5aaa;
    defparam sub_41_add_2_31.INIT1 = 16'h5aaa;
    defparam sub_41_add_2_31.INJECT1_0 = "NO";
    defparam sub_41_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_29 (.A0(phase_inc_carrGen[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[32]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11113), .COUT(n11114), .S0(n1043), .S1(n1042));
    defparam sub_41_add_2_29.INIT0 = 16'h5555;
    defparam sub_41_add_2_29.INIT1 = 16'h5aaa;
    defparam sub_41_add_2_29.INJECT1_0 = "NO";
    defparam sub_41_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_27 (.A0(phase_inc_carrGen[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11112), .COUT(n11113), .S0(n1045), .S1(n1044));
    defparam sub_41_add_2_27.INIT0 = 16'h5555;
    defparam sub_41_add_2_27.INIT1 = 16'h5aaa;
    defparam sub_41_add_2_27.INJECT1_0 = "NO";
    defparam sub_41_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_25 (.A0(phase_inc_carrGen[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11111), .COUT(n11112), .S0(n1047), .S1(n1046));
    defparam sub_41_add_2_25.INIT0 = 16'h5aaa;
    defparam sub_41_add_2_25.INIT1 = 16'h5aaa;
    defparam sub_41_add_2_25.INJECT1_0 = "NO";
    defparam sub_41_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_23 (.A0(phase_inc_carrGen[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11110), .COUT(n11111), .S0(n1049), .S1(n1048));
    defparam sub_41_add_2_23.INIT0 = 16'h5555;
    defparam sub_41_add_2_23.INIT1 = 16'h5555;
    defparam sub_41_add_2_23.INJECT1_0 = "NO";
    defparam sub_41_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_21 (.A0(phase_inc_carrGen[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11109), .COUT(n11110), .S0(n1051), .S1(n1050));
    defparam sub_41_add_2_21.INIT0 = 16'h5555;
    defparam sub_41_add_2_21.INIT1 = 16'h5555;
    defparam sub_41_add_2_21.INJECT1_0 = "NO";
    defparam sub_41_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_19 (.A0(phase_inc_carrGen[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11108), .COUT(n11109), .S0(n1053), .S1(n1052));
    defparam sub_41_add_2_19.INIT0 = 16'h5aaa;
    defparam sub_41_add_2_19.INIT1 = 16'h5aaa;
    defparam sub_41_add_2_19.INJECT1_0 = "NO";
    defparam sub_41_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_17 (.A0(phase_inc_carrGen[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11107), .COUT(n11108), .S0(n1055), .S1(n1054));
    defparam sub_41_add_2_17.INIT0 = 16'h5aaa;
    defparam sub_41_add_2_17.INIT1 = 16'h5555;
    defparam sub_41_add_2_17.INJECT1_0 = "NO";
    defparam sub_41_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_15 (.A0(phase_inc_carrGen[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11106), .COUT(n11107), .S0(n1057), .S1(n1056));
    defparam sub_41_add_2_15.INIT0 = 16'h5555;
    defparam sub_41_add_2_15.INIT1 = 16'h5555;
    defparam sub_41_add_2_15.INJECT1_0 = "NO";
    defparam sub_41_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_13 (.A0(phase_inc_carrGen[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11105), .COUT(n11106), .S0(n1059), .S1(n1058));
    defparam sub_41_add_2_13.INIT0 = 16'h5aaa;
    defparam sub_41_add_2_13.INIT1 = 16'h5555;
    defparam sub_41_add_2_13.INJECT1_0 = "NO";
    defparam sub_41_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_11 (.A0(phase_inc_carrGen[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11104), .COUT(n11105), .S0(n1061), .S1(n1060));
    defparam sub_41_add_2_11.INIT0 = 16'h5555;
    defparam sub_41_add_2_11.INIT1 = 16'h5aaa;
    defparam sub_41_add_2_11.INJECT1_0 = "NO";
    defparam sub_41_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_9 (.A0(phase_inc_carrGen[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11103), .COUT(n11104), .S0(n1063), .S1(n1062));
    defparam sub_41_add_2_9.INIT0 = 16'h5555;
    defparam sub_41_add_2_9.INIT1 = 16'h5aaa;
    defparam sub_41_add_2_9.INJECT1_0 = "NO";
    defparam sub_41_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_7 (.A0(phase_inc_carrGen[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11102), .COUT(n11103), .S0(n1065), .S1(n1064));
    defparam sub_41_add_2_7.INIT0 = 16'h5555;
    defparam sub_41_add_2_7.INIT1 = 16'h5555;
    defparam sub_41_add_2_7.INJECT1_0 = "NO";
    defparam sub_41_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_5 (.A0(phase_inc_carrGen[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11101), .COUT(n11102), .S0(n1067), .S1(n1066));
    defparam sub_41_add_2_5.INIT0 = 16'h5555;
    defparam sub_41_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_41_add_2_5.INJECT1_0 = "NO";
    defparam sub_41_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_3 (.A0(phase_inc_carrGen[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11100), .COUT(n11101), .S0(n1069), .S1(n1068));
    defparam sub_41_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_41_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_41_add_2_3.INJECT1_0 = "NO";
    defparam sub_41_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_41_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(phase_inc_carrGen[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n11100), .S1(n1070));
    defparam sub_41_add_2_1.INIT0 = 16'hF000;
    defparam sub_41_add_2_1.INIT1 = 16'h5555;
    defparam sub_41_add_2_1.INJECT1_0 = "NO";
    defparam sub_41_add_2_1.INJECT1_1 = "NO";
    LUT4 mux_318_i35_4_lut (.A(n7785), .B(n1101), .C(n13376), .D(n13375), 
         .Z(n2308)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i35_4_lut.init = 16'hcfca;
    LUT4 mux_318_i36_4_lut (.A(n7787), .B(n1100), .C(n13376), .D(n13375), 
         .Z(n2307)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i36_4_lut.init = 16'hcfca;
    LUT4 mux_318_i33_4_lut (.A(n7781), .B(n1103), .C(n13376), .D(n13375), 
         .Z(n2310)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i33_4_lut.init = 16'hc0ca;
    LUT4 PWMOut_I_0_1_lut (.A(PWMOutP4_c), .Z(PWMOutN4_c)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(132[19:26])
    defparam PWMOut_I_0_1_lut.init = 16'h5555;
    LUT4 i3504_3_lut (.A(phase_inc_carrGen[33]), .B(n2309), .C(n9000), 
         .Z(n9535)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i3504_3_lut.init = 16'hacac;
    LUT4 mux_318_i34_4_lut (.A(n7783), .B(n1102), .C(n13376), .D(n13375), 
         .Z(n2309)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i34_4_lut.init = 16'hcfca;
    LUT4 mux_318_i31_4_lut (.A(n7777), .B(n1105), .C(n13376), .D(n13375), 
         .Z(n2312)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i31_4_lut.init = 16'hc0ca;
    LUT4 i3558_3_lut (.A(phase_inc_carrGen[6]), .B(n8000), .C(n9000), 
         .Z(n9589)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i3558_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_rep_72 (.A(o_Rx_Byte_c_4), .B(n12803), .Z(n13383)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_72.init = 16'h8888;
    LUT4 i1965_4_lut (.A(n1129), .B(n1068), .C(o_Rx_Byte_c_3), .D(n13383), 
         .Z(n8000)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1965_4_lut.init = 16'hcacf;
    LUT4 i5699_4_lut (.A(n13384), .B(n13372), .C(n8225), .D(o_Rx_Byte_c_2), 
         .Z(n9000)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B))) */ ;
    defparam i5699_4_lut.init = 16'h1333;
    LUT4 o_Rx_Byte_c_0_bdd_4_lut_5762 (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(n7349), .D(o_Rx_Byte_c_3), .Z(n13291)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;
    defparam o_Rx_Byte_c_0_bdd_4_lut_5762.init = 16'hc9d0;
    LUT4 i3562_3_lut (.A(phase_inc_carrGen[4]), .B(n2338), .C(n9000), 
         .Z(n9593)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i3562_3_lut.init = 16'hacac;
    LUT4 i1_4_lut (.A(o_Rx_Byte_c_2), .B(n8225), .C(o_Rx_Byte_c_0), .D(n7349), 
         .Z(n12803)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut.init = 16'h0040;
    SinCos SinCos1 (.osc_clk(osc_clk), .VCC_net(VCC_net), .GND_net(GND_net), 
           .\phase_accum[57] (phase_accum[57]), .\phase_accum[58] (phase_accum[58]), 
           .\phase_accum[59] (phase_accum[59]), .\phase_accum[60] (phase_accum[60]), 
           .\phase_accum[61] (phase_accum[61]), .\phase_accum[62] (phase_accum[62]), 
           .\phase_accum[63] (phase_accum[63]), .\LOSine[1] (LOSine[1]), 
           .\LOSine[2] (LOSine[2]), .\LOSine[3] (LOSine[3]), .\LOSine[4] (LOSine[4]), 
           .\LOSine[5] (LOSine[5]), .\LOSine[6] (LOSine[6]), .\LOSine[7] (LOSine[7]), 
           .\LOSine[8] (LOSine[8]), .\LOSine[9] (LOSine[9]), .\LOSine[10] (LOSine[10]), 
           .\LOSine[11] (LOSine[11]), .\LOSine[12] (LOSine[12]), .\LOCosine[1] (LOCosine[1]), 
           .\LOCosine[2] (LOCosine[2]), .\LOCosine[3] (LOCosine[3]), .\LOCosine[4] (LOCosine[4]), 
           .\LOCosine[5] (LOCosine[5]), .\LOCosine[6] (LOCosine[6]), .\LOCosine[7] (LOCosine[7]), 
           .\LOCosine[8] (LOCosine[8]), .\LOCosine[9] (LOCosine[9]), .\LOCosine[10] (LOCosine[10]), 
           .\LOCosine[11] (LOCosine[11]), .\LOCosine[12] (LOCosine[12]), 
           .\phase_accum[56] (phase_accum[56])) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    LUT4 mux_318_i5_4_lut (.A(n7733), .B(n1131), .C(n13376), .D(n13375), 
         .Z(n2338)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i5_4_lut.init = 16'hc0ca;
    LUT4 i3560_3_lut (.A(phase_inc_carrGen[5]), .B(n2337), .C(n9000), 
         .Z(n9591)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i3560_3_lut.init = 16'hacac;
    LUT4 mux_318_i6_4_lut (.A(n7735), .B(n1130), .C(n13376), .D(n13375), 
         .Z(n2337)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i6_4_lut.init = 16'hcfca;
    LUT4 mux_318_i32_4_lut (.A(n7779), .B(n1104), .C(n13376), .D(n13375), 
         .Z(n2311)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i32_4_lut.init = 16'hcfca;
    LUT4 mux_318_i3_4_lut (.A(o_Rx_Byte_c_3), .B(n1133), .C(n13376), .D(n13380), 
         .Z(n2340)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i3_4_lut.init = 16'hc0c5;
    LUT4 i1794_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1021), .Z(n7817)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;
    defparam i1794_3_lut_4_lut.init = 16'hf707;
    LUT4 i2_4_lut (.A(o_Rx_Byte_c_2), .B(n12879), .C(n7349), .D(o_Rx_Byte_c_3), 
         .Z(n12970)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i2_4_lut.init = 16'hfffb;
    LUT4 i1786_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1026), .Z(n7809)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i1786_3_lut_4_lut.init = 16'hf808;
    LUT4 i5413_2_lut (.A(o_Rx_Byte_c_4), .B(o_Rx_Byte_c_0), .Z(n12879)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i5413_2_lut.init = 16'heeee;
    LUT4 mux_318_i29_4_lut (.A(n7773), .B(n1107), .C(n13376), .D(n13375), 
         .Z(n2314)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i29_4_lut.init = 16'hc0ca;
    LUT4 mux_318_i30_4_lut (.A(n2513), .B(n1106), .C(n13376), .D(n13375), 
         .Z(n2313)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i30_4_lut.init = 16'hc0ca;
    LUT4 mux_318_i27_4_lut (.A(n7769), .B(n1109), .C(n13376), .D(n13375), 
         .Z(n2316)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i27_4_lut.init = 16'hc0ca;
    LUT4 mux_318_i2_4_lut (.A(n8341), .B(n1134), .C(n13376), .D(n13375), 
         .Z(n2341)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i2_4_lut.init = 16'hcfc5;
    LUT4 i3516_3_lut (.A(phase_inc_carrGen[27]), .B(n2315), .C(n9000), 
         .Z(n9547)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i3516_3_lut.init = 16'hacac;
    LUT4 mux_318_i28_4_lut (.A(n7771), .B(n1108), .C(n13376), .D(n13375), 
         .Z(n2315)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i28_4_lut.init = 16'hcfca;
    LUT4 mux_318_i25_4_lut (.A(n7765), .B(n1111), .C(n13376), .D(n13375), 
         .Z(n2318)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i25_4_lut.init = 16'hc0ca;
    LUT4 mux_318_i26_4_lut (.A(n7767), .B(n1110), .C(n13376), .D(n13375), 
         .Z(n2317)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i26_4_lut.init = 16'hc0ca;
    LUT4 mux_318_i23_4_lut (.A(n13375), .B(n1113), .C(n13376), .D(n28), 
         .Z(n2320)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i23_4_lut.init = 16'hcfca;
    LUT4 mux_318_i24_4_lut (.A(n7763), .B(n1112), .C(n13376), .D(n13375), 
         .Z(n2319)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i24_4_lut.init = 16'hcfca;
    LUT4 mux_318_i21_4_lut (.A(n7759), .B(n1115), .C(n13376), .D(n13375), 
         .Z(n2322)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i21_4_lut.init = 16'hcfca;
    LUT4 i1782_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1028), .Z(n7805)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;
    defparam i1782_3_lut_4_lut.init = 16'hf707;
    LUT4 mux_318_i22_4_lut (.A(n2521), .B(n1114), .C(n13376), .D(n13375), 
         .Z(n2321)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i22_4_lut.init = 16'hcfca;
    LUT4 i3022_2_lut (.A(n1053), .B(o_Rx_Byte_c_3), .Z(n2521)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i3022_2_lut.init = 16'h8888;
    LUT4 mux_318_i19_4_lut (.A(n7755), .B(n1117), .C(n13376), .D(n13375), 
         .Z(n2324)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i19_4_lut.init = 16'hc0ca;
    Mixer Mixer1 (.\LOCosine[12] (LOCosine[12]), .MixerOutSin({MixerOutSin}), 
          .osc_clk(osc_clk), .DiffOut_c(DiffOut_c), .MixerOutCos({MixerOutCos}), 
          .RFIn_c(RFIn_c), .GND_net(GND_net), .\LOCosine[10] (LOCosine[10]), 
          .\LOCosine[11] (LOCosine[11]), .\LOCosine[8] (LOCosine[8]), .\LOCosine[9] (LOCosine[9]), 
          .\LOCosine[6] (LOCosine[6]), .\LOCosine[7] (LOCosine[7]), .\LOCosine[4] (LOCosine[4]), 
          .\LOCosine[5] (LOCosine[5]), .\LOCosine[2] (LOCosine[2]), .\LOCosine[3] (LOCosine[3]), 
          .\LOCosine[1] (LOCosine[1]), .\LOSine[12] (LOSine[12]), .\LOSine[10] (LOSine[10]), 
          .\LOSine[11] (LOSine[11]), .\LOSine[8] (LOSine[8]), .\LOSine[9] (LOSine[9]), 
          .\LOSine[6] (LOSine[6]), .\LOSine[7] (LOSine[7]), .\LOSine[4] (LOSine[4]), 
          .\LOSine[5] (LOSine[5]), .\LOSine[2] (LOSine[2]), .\LOSine[3] (LOSine[3]), 
          .\LOSine[1] (LOSine[1])) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(157[7] 165[2])
    FD1P3AX phase_inc_carrGen_i0_i2 (.D(n2858), .SP(osc_clk_enable_1397), 
            .CK(osc_clk), .Q(phase_inc_carrGen[2]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i2.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i3 (.D(n2857), .SP(osc_clk_enable_1397), 
            .CK(osc_clk), .Q(phase_inc_carrGen[3]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i3.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i4 (.D(n2856), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[4]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i4.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i5 (.D(n2855), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[5]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i5.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i6 (.D(n2854), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[6]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i6.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i7 (.D(n2853), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[7]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i7.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i8 (.D(n2852), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[8]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i8.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i9 (.D(n2851), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[9]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i9.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i10 (.D(n2850), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[10]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i10.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i11 (.D(n2849), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[11]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i11.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i12 (.D(n2848), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[12]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i12.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i13 (.D(n2847), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[13]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i13.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i14 (.D(n2846), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[14]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i14.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i15 (.D(n2845), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[15]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i15.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i16 (.D(n2844), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[16]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i16.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i17 (.D(n2843), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[17]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i17.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i18 (.D(n2842), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[18]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i18.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i19 (.D(n2841), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[19]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i19.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i20 (.D(n2840), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[20]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i20.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i21 (.D(n2839), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[21]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i21.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i22 (.D(n2838), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[22]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i22.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i23 (.D(n2837), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[23]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i23.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i24 (.D(n2836), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[24]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i24.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i25 (.D(n2835), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[25]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i25.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i26 (.D(n2834), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[26]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i26.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i27 (.D(n2833), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[27]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i27.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i28 (.D(n2832), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[28]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i28.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i29 (.D(n2831), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[29]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i29.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i30 (.D(n2830), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[30]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i30.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i31 (.D(n2829), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[31]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i31.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i32 (.D(n2828), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[32]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i32.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i33 (.D(n2827), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[33]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i33.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i34 (.D(n2826), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[34]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i34.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i35 (.D(n2825), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[35]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i35.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i36 (.D(n2824), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[36]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i36.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i37 (.D(n2823), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[37]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i37.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i38 (.D(n2822), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[38]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i38.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i39 (.D(n2821), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[39]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i39.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i40 (.D(n2820), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[40]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i40.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i41 (.D(n2819), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[41]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i41.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i42 (.D(n2818), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[42]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i42.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i43 (.D(n2817), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[43]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i43.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i44 (.D(n2816), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[44]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i44.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i45 (.D(n2815), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[45]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i45.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i46 (.D(n2814), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[46]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i46.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i47 (.D(n2813), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[47]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i47.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i48 (.D(n2812), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[48]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i48.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i49 (.D(n2811), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[49]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i49.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i50 (.D(n2810), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[50]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i50.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i51 (.D(n2809), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[51]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i51.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i52 (.D(n2808), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[52]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i52.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i53 (.D(n2807), .SP(osc_clk_enable_1447), 
            .CK(osc_clk), .Q(phase_inc_carrGen[53]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i53.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i54 (.D(n2806), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[54]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i54.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i55 (.D(n2805), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[55]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i55.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i56 (.D(n2804), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[56]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i56.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i57 (.D(n2803), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[57]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i57.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i58 (.D(n2802), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[58]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i58.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i59 (.D(n2801), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[59]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i59.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i60 (.D(n2800), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[60]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i60.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i61 (.D(n2799), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[61]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i61.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i62 (.D(n2798), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[62]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i62.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i63 (.D(n2797), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[63]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(235[8] 282[4])
    defparam phase_inc_carrGen_i0_i63.GSR = "ENABLED";
    LUT4 i5751_4_lut (.A(o_Rx_Byte_c_2), .B(n13390), .C(o_Rx_Byte_c_6), 
         .D(n6), .Z(osc_clk_enable_1394)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i5751_4_lut.init = 16'h0004;
    LUT4 i3532_3_lut (.A(phase_inc_carrGen[19]), .B(n8006), .C(n9000), 
         .Z(n9563)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i3532_3_lut.init = 16'hacac;
    LUT4 i1971_4_lut (.A(n1116), .B(n1055), .C(o_Rx_Byte_c_3), .D(n13383), 
         .Z(n8006)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1971_4_lut.init = 16'hcac0;
    LUT4 mux_318_i17_4_lut (.A(n7751), .B(n1119), .C(n13376), .D(n13375), 
         .Z(n2326)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i17_4_lut.init = 16'hcfca;
    LUT4 i1969_4_lut (.A(n1118), .B(n1057), .C(o_Rx_Byte_c_3), .D(n13383), 
         .Z(n8004)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1969_4_lut.init = 16'hcac0;
    GSR GSR_INST (.GSR(VCC_net));
    LUT4 mux_318_i15_4_lut (.A(n7749), .B(n1121), .C(n13376), .D(n13375), 
         .Z(n2328)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i15_4_lut.init = 16'hcfca;
    LUT4 i5737_3_lut (.A(o_Rx_Byte_c_3), .B(n13523), .C(n9000), .Z(osc_clk_enable_1397)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;
    defparam i5737_3_lut.init = 16'hc4c4;
    LUT4 i3540_3_lut (.A(phase_inc_carrGen[15]), .B(n2327), .C(n9000), 
         .Z(n9571)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i3540_3_lut.init = 16'hacac;
    LUT4 i1979_4_lut (.A(n1073), .B(n1012), .C(o_Rx_Byte_c_3), .D(n13383), 
         .Z(n8014)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1979_4_lut.init = 16'hcac0;
    LUT4 mux_318_i16_4_lut (.A(n13375), .B(n1120), .C(n13376), .D(n29), 
         .Z(n2327)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i16_4_lut.init = 16'hcfca;
    LUT4 i1981_4_lut (.A(n1072), .B(n1011), .C(o_Rx_Byte_c_3), .D(n13383), 
         .Z(n8016)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1981_4_lut.init = 16'hcac0;
    LUT4 mux_318_i61_4_lut (.A(n7829), .B(n1075), .C(n13376), .D(n13375), 
         .Z(n2282)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i61_4_lut.init = 16'hc0ca;
    LUT4 mux_318_i13_4_lut (.A(n2530), .B(n1123), .C(n13376), .D(n13375), 
         .Z(n2330)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i13_4_lut.init = 16'hc0ca;
    LUT4 i1977_4_lut (.A(n1074), .B(n1013), .C(o_Rx_Byte_c_3), .D(n13383), 
         .Z(n8012)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1977_4_lut.init = 16'hcac0;
    LUT4 i1967_4_lut (.A(n1122), .B(n1061), .C(o_Rx_Byte_c_3), .D(n13383), 
         .Z(n8002)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i1967_4_lut.init = 16'hcac0;
    LUT4 mux_318_i11_4_lut (.A(n7743), .B(n1125), .C(n13376), .D(n13375), 
         .Z(n2332)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i11_4_lut.init = 16'hcfca;
    LUT4 mux_318_i12_4_lut (.A(n2531), .B(n1124), .C(n13376), .D(n13375), 
         .Z(n2331)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i12_4_lut.init = 16'hcfca;
    LUT4 i3017_2_lut (.A(n1063), .B(o_Rx_Byte_c_3), .Z(n2531)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i3017_2_lut.init = 16'h8888;
    LUT4 mux_318_i9_4_lut (.A(n7739), .B(n1127), .C(n13376), .D(n13375), 
         .Z(n2334)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i9_4_lut.init = 16'hcfca;
    LUT4 mux_318_i10_4_lut (.A(n7741), .B(n1126), .C(n13376), .D(n13375), 
         .Z(n2333)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i10_4_lut.init = 16'hcfca;
    LUT4 mux_318_i59_4_lut (.A(n7825), .B(n1077), .C(n13376), .D(n13375), 
         .Z(n2284)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i59_4_lut.init = 16'hc0ca;
    LUT4 mux_318_i60_4_lut (.A(n7827), .B(n1076), .C(n13376), .D(n13375), 
         .Z(n2283)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i60_4_lut.init = 16'hc0ca;
    LUT4 i1762_3_lut_4_lut (.A(o_Rx_Byte_c_2), .B(n13381), .C(o_Rx_Byte_c_3), 
         .D(n1040), .Z(n7785)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i1762_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_318_i57_4_lut (.A(n2486), .B(n1079), .C(n13376), .D(n13375), 
         .Z(n2286)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i57_4_lut.init = 16'hc0ca;
    nco_sig ncoGen (.osc_clk(osc_clk), .\phase_accum[56] (phase_accum[56]), 
            .\phase_accum[57] (phase_accum[57]), .\phase_accum[58] (phase_accum[58]), 
            .\phase_accum[59] (phase_accum[59]), .\phase_accum[60] (phase_accum[60]), 
            .\phase_accum[61] (phase_accum[61]), .\phase_accum[62] (phase_accum[62]), 
            .\phase_accum[63] (phase_accum[63]), .phase_inc_carrGen1({phase_inc_carrGen1}), 
            .GND_net(GND_net), .sinGen_c(sinGen_c)) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(148[10] 154[2])
    LUT4 mux_318_i58_4_lut (.A(n2485), .B(n1078), .C(n13376), .D(n13375), 
         .Z(n2285)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam mux_318_i58_4_lut.init = 16'hcfca;
    \CIC(width=72,decimation_ratio=4096)  CIC1Sin (.osc_clk(osc_clk), .MixerOutSin({MixerOutSin}), 
            .GND_net(GND_net), .CIC1_out_clkSin(CIC1_out_clkSin), .\CICGain[1] (CICGain[1]), 
            .\CICGain[0] (CICGain[0]), .\CIC1_outSin[0] (CIC1_outSin[0]), 
            .n63(n63), .\d_out_11__N_1819[2] (d_out_11__N_1819_adj_2575[2]), 
            .n64(n64), .\d_out_11__N_1819[3] (d_out_11__N_1819_adj_2575[3]), 
            .n65(n65), .\d_out_11__N_1819[4] (d_out_11__N_1819_adj_2575[4]), 
            .n66(n66), .\d_out_11__N_1819[5] (d_out_11__N_1819_adj_2575[5]), 
            .n67(n67), .\d_out_11__N_1819[6] (d_out_11__N_1819_adj_2575[6]), 
            .n68(n68), .\d_out_11__N_1819[7] (d_out_11__N_1819_adj_2575[7]), 
            .\d10[68] (d10_adj_2550[68]), .\d_out_11__N_1819[8] (d_out_11__N_1819_adj_2575[8]), 
            .n70(n70), .\d_out_11__N_1819[9] (d_out_11__N_1819_adj_2575[9]), 
            .\d10[71] (d10_adj_2550[71]), .\d_out_11__N_1819[11] (d_out_11__N_1819_adj_2575[11]), 
            .\d10[65] (d10_adj_2550[65]), .\d10[66] (d10_adj_2550[66]), 
            .\d10[63] (d10_adj_2550[63]), .\d10[64] (d10_adj_2550[64]), 
            .\d10[61] (d10_adj_2550[61]), .\d10[62] (d10_adj_2550[62]), 
            .n61(n61), .\d10[59] (d10_adj_2550[59]), .n62(n62), .\d10[60] (d10_adj_2550[60]), 
            .\CIC1_outSin[1] (CIC1_outSin[1]), .\CIC1_outSin[2] (CIC1_outSin[2]), 
            .\CIC1_outSin[3] (CIC1_outSin[3]), .\CIC1_outSin[4] (CIC1_outSin[4]), 
            .\CIC1_outSin[5] (CIC1_outSin[5]), .MYLED_c_0(MYLED_c_0), .MYLED_c_1(MYLED_c_1), 
            .MYLED_c_2(MYLED_c_2), .MYLED_c_3(MYLED_c_3), .MYLED_c_4(MYLED_c_4), 
            .MYLED_c_5(MYLED_c_5), .\d10[67] (d10_adj_2550[67]), .\d10[69] (d10_adj_2550[69]), 
            .\d10[70] (d10_adj_2550[70]), .\d_out_11__N_1819[10] (d_out_11__N_1819_adj_2575[10])) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(168[45] 174[2])
    LUT4 i3033_2_lut (.A(n1017), .B(o_Rx_Byte_c_3), .Z(n2485)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(239[2] 281[6])
    defparam i3033_2_lut.init = 16'h8888;
    \CIC(width=72,decimation_ratio=4096)_U1  CIC1Cos (.GND_net(GND_net), .MixerOutCos({MixerOutCos}), 
            .osc_clk(osc_clk), .CIC1_outCos({CIC1_outCos}), .\d10[59] (d10_adj_2550[59]), 
            .\d10[60] (d10_adj_2550[60]), .\d10[61] (d10_adj_2550[61]), 
            .\d10[62] (d10_adj_2550[62]), .\d10[63] (d10_adj_2550[63]), 
            .\d10[64] (d10_adj_2550[64]), .\d10[65] (d10_adj_2550[65]), 
            .\d10[66] (d10_adj_2550[66]), .\d10[67] (d10_adj_2550[67]), 
            .\d10[68] (d10_adj_2550[68]), .\d10[69] (d10_adj_2550[69]), 
            .\d10[70] (d10_adj_2550[70]), .\d10[71] (d10_adj_2550[71]), 
            .\d_out_11__N_1819[2] (d_out_11__N_1819_adj_2575[2]), .\d_out_11__N_1819[3] (d_out_11__N_1819_adj_2575[3]), 
            .\d_out_11__N_1819[4] (d_out_11__N_1819_adj_2575[4]), .\d_out_11__N_1819[5] (d_out_11__N_1819_adj_2575[5]), 
            .\d_out_11__N_1819[6] (d_out_11__N_1819_adj_2575[6]), .\d_out_11__N_1819[7] (d_out_11__N_1819_adj_2575[7]), 
            .\d_out_11__N_1819[8] (d_out_11__N_1819_adj_2575[8]), .\d_out_11__N_1819[9] (d_out_11__N_1819_adj_2575[9]), 
            .\d_out_11__N_1819[10] (d_out_11__N_1819_adj_2575[10]), .\d_out_11__N_1819[11] (d_out_11__N_1819_adj_2575[11]), 
            .\CICGain[0] (CICGain[0]), .n61(n61), .n70(n70), .\CICGain[1] (CICGain[1]), 
            .n62(n62), .n63(n63), .n64(n64), .n65(n65), .n66(n66), 
            .n67(n67), .n68(n68)) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(177[45] 183[2])
    AMDemodulator AMDemodulator1 (.CIC1_out_clkSin(CIC1_out_clkSin), .\CIC1_outSin[0] (CIC1_outSin[0]), 
            .CIC1_outCos({CIC1_outCos}), .\DataInReg_11__N_1856[0] (DataInReg_11__N_1856[0]), 
            .GND_net(GND_net), .\CIC1_outSin[1] (CIC1_outSin[1]), .\CIC1_outSin[2] (CIC1_outSin[2]), 
            .\CIC1_outSin[3] (CIC1_outSin[3]), .\CIC1_outSin[4] (CIC1_outSin[4]), 
            .\CIC1_outSin[5] (CIC1_outSin[5]), .MYLED_c_0(MYLED_c_0), .MYLED_c_1(MYLED_c_1), 
            .MYLED_c_2(MYLED_c_2), .MYLED_c_3(MYLED_c_3), .MYLED_c_4(MYLED_c_4), 
            .MYLED_c_5(MYLED_c_5), .\DataInReg_11__N_1856[1] (DataInReg_11__N_1856[1]), 
            .\DataInReg_11__N_1856[2] (DataInReg_11__N_1856[2]), .\DataInReg_11__N_1856[3] (DataInReg_11__N_1856[3]), 
            .\DataInReg_11__N_1856[4] (DataInReg_11__N_1856[4]), .\DataInReg_11__N_1856[5] (DataInReg_11__N_1856[5]), 
            .\DataInReg_11__N_1856[6] (DataInReg_11__N_1856[6]), .\DataInReg_11__N_1856[7] (DataInReg_11__N_1856[7]), 
            .\DataInReg_11__N_1856[8] (DataInReg_11__N_1856[8]), .\DemodOut[9] (DemodOut[9]), 
            .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(209[15] 214[10])
    
endmodule
//
// Verilog Description of module PWM
//

module PWM (osc_clk, \DataInReg_11__N_1856[0] , PWMOutP4_c, GND_net, 
            \DataInReg_11__N_1856[1] , \DataInReg_11__N_1856[2] , \DataInReg_11__N_1856[3] , 
            \DataInReg_11__N_1856[4] , \DataInReg_11__N_1856[5] , \DataInReg_11__N_1856[6] , 
            \DataInReg_11__N_1856[7] , \DataInReg_11__N_1856[8] , \DemodOut[9] ) /* synthesis syn_module_defined=1 */ ;
    input osc_clk;
    input \DataInReg_11__N_1856[0] ;
    output PWMOutP4_c;
    input GND_net;
    input \DataInReg_11__N_1856[1] ;
    input \DataInReg_11__N_1856[2] ;
    input \DataInReg_11__N_1856[3] ;
    input \DataInReg_11__N_1856[4] ;
    input \DataInReg_11__N_1856[5] ;
    input \DataInReg_11__N_1856[6] ;
    input \DataInReg_11__N_1856[7] ;
    input \DataInReg_11__N_1856[8] ;
    input \DemodOut[9] ;
    
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(71[8:15])
    wire [11:0]DataInReg;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(10[12:21])
    
    wire osc_clk_enable_1393, PWMOut_N_1869;
    wire [9:0]counter;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(7[11:18])
    wire [9:0]n45;
    
    wire n11802, n11801, n11800, n11799, n11798;
    wire [11:0]n3926;
    
    wire n11267, n11266, n11265, n11264, n11263, n17, n15, n11, 
        n12;
    
    FD1P3AX DataInReg__i1 (.D(\DataInReg_11__N_1856[0] ), .SP(osc_clk_enable_1393), 
            .CK(osc_clk), .Q(DataInReg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i1.GSR = "ENABLED";
    FD1S3AX PWMOut_15 (.D(PWMOut_N_1869), .CK(osc_clk), .Q(PWMOutP4_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam PWMOut_15.GSR = "ENABLED";
    FD1S3AX counter_999__i0 (.D(n45[0]), .CK(osc_clk), .Q(counter[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_999__i0.GSR = "ENABLED";
    CCU2D counter_999_add_4_11 (.A0(counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11802), .S0(n45[9]));   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_999_add_4_11.INIT0 = 16'hfaaa;
    defparam counter_999_add_4_11.INIT1 = 16'h0000;
    defparam counter_999_add_4_11.INJECT1_0 = "NO";
    defparam counter_999_add_4_11.INJECT1_1 = "NO";
    CCU2D counter_999_add_4_9 (.A0(counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11801), .COUT(n11802), .S0(n45[7]), .S1(n45[8]));   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_999_add_4_9.INIT0 = 16'hfaaa;
    defparam counter_999_add_4_9.INIT1 = 16'hfaaa;
    defparam counter_999_add_4_9.INJECT1_0 = "NO";
    defparam counter_999_add_4_9.INJECT1_1 = "NO";
    CCU2D counter_999_add_4_7 (.A0(counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11800), .COUT(n11801), .S0(n45[5]), .S1(n45[6]));   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_999_add_4_7.INIT0 = 16'hfaaa;
    defparam counter_999_add_4_7.INIT1 = 16'hfaaa;
    defparam counter_999_add_4_7.INJECT1_0 = "NO";
    defparam counter_999_add_4_7.INJECT1_1 = "NO";
    CCU2D counter_999_add_4_5 (.A0(counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11799), .COUT(n11800), .S0(n45[3]), .S1(n45[4]));   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_999_add_4_5.INIT0 = 16'hfaaa;
    defparam counter_999_add_4_5.INIT1 = 16'hfaaa;
    defparam counter_999_add_4_5.INJECT1_0 = "NO";
    defparam counter_999_add_4_5.INJECT1_1 = "NO";
    CCU2D counter_999_add_4_3 (.A0(counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11798), .COUT(n11799), .S0(n45[1]), .S1(n45[2]));   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_999_add_4_3.INIT0 = 16'hfaaa;
    defparam counter_999_add_4_3.INIT1 = 16'hfaaa;
    defparam counter_999_add_4_3.INJECT1_0 = "NO";
    defparam counter_999_add_4_3.INJECT1_1 = "NO";
    CCU2D counter_999_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n11798), .S1(n45[0]));   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_999_add_4_1.INIT0 = 16'hF000;
    defparam counter_999_add_4_1.INIT1 = 16'h0555;
    defparam counter_999_add_4_1.INJECT1_0 = "NO";
    defparam counter_999_add_4_1.INJECT1_1 = "NO";
    FD1P3AX DataInReg__i2 (.D(\DataInReg_11__N_1856[1] ), .SP(osc_clk_enable_1393), 
            .CK(osc_clk), .Q(DataInReg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i2.GSR = "ENABLED";
    FD1P3AX DataInReg__i3 (.D(\DataInReg_11__N_1856[2] ), .SP(osc_clk_enable_1393), 
            .CK(osc_clk), .Q(DataInReg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i3.GSR = "ENABLED";
    FD1P3AX DataInReg__i4 (.D(\DataInReg_11__N_1856[3] ), .SP(osc_clk_enable_1393), 
            .CK(osc_clk), .Q(DataInReg[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i4.GSR = "ENABLED";
    FD1P3AX DataInReg__i5 (.D(\DataInReg_11__N_1856[4] ), .SP(osc_clk_enable_1393), 
            .CK(osc_clk), .Q(DataInReg[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i5.GSR = "ENABLED";
    FD1P3AX DataInReg__i6 (.D(\DataInReg_11__N_1856[5] ), .SP(osc_clk_enable_1393), 
            .CK(osc_clk), .Q(DataInReg[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i6.GSR = "ENABLED";
    FD1P3AX DataInReg__i7 (.D(\DataInReg_11__N_1856[6] ), .SP(osc_clk_enable_1393), 
            .CK(osc_clk), .Q(DataInReg[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i7.GSR = "ENABLED";
    FD1P3AX DataInReg__i8 (.D(\DataInReg_11__N_1856[7] ), .SP(osc_clk_enable_1393), 
            .CK(osc_clk), .Q(DataInReg[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i8.GSR = "ENABLED";
    FD1P3AX DataInReg__i9 (.D(\DataInReg_11__N_1856[8] ), .SP(osc_clk_enable_1393), 
            .CK(osc_clk), .Q(DataInReg[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i9.GSR = "ENABLED";
    FD1P3AX DataInReg__i10 (.D(n3926[9]), .SP(osc_clk_enable_1393), .CK(osc_clk), 
            .Q(DataInReg[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=192 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i10.GSR = "ENABLED";
    FD1S3AX counter_999__i1 (.D(n45[1]), .CK(osc_clk), .Q(counter[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_999__i1.GSR = "ENABLED";
    FD1S3AX counter_999__i2 (.D(n45[2]), .CK(osc_clk), .Q(counter[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_999__i2.GSR = "ENABLED";
    FD1S3AX counter_999__i3 (.D(n45[3]), .CK(osc_clk), .Q(counter[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_999__i3.GSR = "ENABLED";
    FD1S3AX counter_999__i4 (.D(n45[4]), .CK(osc_clk), .Q(counter[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_999__i4.GSR = "ENABLED";
    FD1S3AX counter_999__i5 (.D(n45[5]), .CK(osc_clk), .Q(counter[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_999__i5.GSR = "ENABLED";
    FD1S3AX counter_999__i6 (.D(n45[6]), .CK(osc_clk), .Q(counter[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_999__i6.GSR = "ENABLED";
    FD1S3AX counter_999__i7 (.D(n45[7]), .CK(osc_clk), .Q(counter[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_999__i7.GSR = "ENABLED";
    FD1S3AX counter_999__i8 (.D(n45[8]), .CK(osc_clk), .Q(counter[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_999__i8.GSR = "ENABLED";
    FD1S3AX counter_999__i9 (.D(n45[9]), .CK(osc_clk), .Q(counter[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_999__i9.GSR = "ENABLED";
    CCU2D sub_761_add_2_11 (.A0(DataInReg[9]), .B0(counter[9]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11267), .S1(PWMOut_N_1869));
    defparam sub_761_add_2_11.INIT0 = 16'h5999;
    defparam sub_761_add_2_11.INIT1 = 16'h0000;
    defparam sub_761_add_2_11.INJECT1_0 = "NO";
    defparam sub_761_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_761_add_2_9 (.A0(DataInReg[7]), .B0(counter[7]), .C0(GND_net), 
          .D0(GND_net), .A1(DataInReg[8]), .B1(counter[8]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11266), .COUT(n11267));
    defparam sub_761_add_2_9.INIT0 = 16'h5999;
    defparam sub_761_add_2_9.INIT1 = 16'h5999;
    defparam sub_761_add_2_9.INJECT1_0 = "NO";
    defparam sub_761_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_761_add_2_7 (.A0(DataInReg[5]), .B0(counter[5]), .C0(GND_net), 
          .D0(GND_net), .A1(DataInReg[6]), .B1(counter[6]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11265), .COUT(n11266));
    defparam sub_761_add_2_7.INIT0 = 16'h5999;
    defparam sub_761_add_2_7.INIT1 = 16'h5999;
    defparam sub_761_add_2_7.INJECT1_0 = "NO";
    defparam sub_761_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_761_add_2_5 (.A0(DataInReg[3]), .B0(counter[3]), .C0(GND_net), 
          .D0(GND_net), .A1(DataInReg[4]), .B1(counter[4]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11264), .COUT(n11265));
    defparam sub_761_add_2_5.INIT0 = 16'h5999;
    defparam sub_761_add_2_5.INIT1 = 16'h5999;
    defparam sub_761_add_2_5.INJECT1_0 = "NO";
    defparam sub_761_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_761_add_2_3 (.A0(DataInReg[1]), .B0(counter[1]), .C0(GND_net), 
          .D0(GND_net), .A1(DataInReg[2]), .B1(counter[2]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11263), .COUT(n11264));
    defparam sub_761_add_2_3.INIT0 = 16'h5999;
    defparam sub_761_add_2_3.INIT1 = 16'h5999;
    defparam sub_761_add_2_3.INJECT1_0 = "NO";
    defparam sub_761_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_761_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(DataInReg[0]), .B1(counter[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n11263));
    defparam sub_761_add_2_1.INIT0 = 16'h0000;
    defparam sub_761_add_2_1.INIT1 = 16'h5999;
    defparam sub_761_add_2_1.INJECT1_0 = "NO";
    defparam sub_761_add_2_1.INJECT1_1 = "NO";
    LUT4 i5754_4_lut (.A(n17), .B(n15), .C(n11), .D(n12), .Z(osc_clk_enable_1393)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(26[7:19])
    defparam i5754_4_lut.init = 16'h0001;
    LUT4 i7_4_lut (.A(counter[3]), .B(counter[2]), .C(counter[1]), .D(counter[9]), 
         .Z(n17)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(26[7:19])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut (.A(counter[6]), .B(counter[4]), .Z(n15)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(26[7:19])
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i1147_1_lut (.A(\DemodOut[9] ), .Z(n3926[9])) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(26[3] 27[35])
    defparam i1147_1_lut.init = 16'h5555;
    LUT4 i1_2_lut (.A(counter[0]), .B(counter[5]), .Z(n11)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(26[7:19])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i2_2_lut (.A(counter[7]), .B(counter[8]), .Z(n12)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(26[7:19])
    defparam i2_2_lut.init = 16'heeee;
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module \uart_rx(CLKS_PER_BIT=87) 
//

module \uart_rx(CLKS_PER_BIT=87)  (o_Rx_Byte_c_2, n8225, n2795, o_Rx_Byte_c_4, 
            n13291, n12970, n13523, osc_clk, i_Rx_Serial_c, o_Rx_Byte_c_0, 
            osc_clk_enable_1447, n3614, o_Rx_Byte_c_3, n6, n12803, 
            n13380, n3628, osc_clk_enable_1457, n7349, n13385, n2608, 
            n1132, n13383, n2339, n1030, n2364, n1018, n2486, 
            n12919, n12931, n13372, n1034, n13381, n30, n7970, 
            n13376, n13375, n1052, n28, n1045, n2513, n1059, n29, 
            GND_net, o_Rx_Byte_c_5, o_Rx_Byte_c_6, o_Rx_Byte_c_7, n9000, 
            osc_clk_enable_128, n1128, n1067, n13384, n1062, n2530, 
            o_Rx_DV_c, n13411) /* synthesis syn_module_defined=1 */ ;
    output o_Rx_Byte_c_2;
    input n8225;
    output n2795;
    output o_Rx_Byte_c_4;
    input n13291;
    input n12970;
    output n13523;
    input osc_clk;
    input i_Rx_Serial_c;
    output o_Rx_Byte_c_0;
    output osc_clk_enable_1447;
    output n3614;
    output o_Rx_Byte_c_3;
    output n6;
    input n12803;
    output n13380;
    output n3628;
    output osc_clk_enable_1457;
    output n7349;
    output n13385;
    output n2608;
    input n1132;
    input n13383;
    output n2339;
    input n1030;
    output n2364;
    input n1018;
    output n2486;
    input n12919;
    input n12931;
    output n13372;
    input n1034;
    input n13381;
    output n30;
    output n7970;
    output n13376;
    output n13375;
    input n1052;
    output n28;
    input n1045;
    output n2513;
    input n1059;
    output n29;
    input GND_net;
    output o_Rx_Byte_c_5;
    output o_Rx_Byte_c_6;
    output o_Rx_Byte_c_7;
    input n9000;
    output osc_clk_enable_128;
    input n1128;
    input n1067;
    input n13384;
    input n1062;
    output n2530;
    output o_Rx_DV_c;
    output n13411;
    
    wire [7:0]UartClk /* synthesis SET_AS_NETWORK=\uart_rx1/UartClk[2], is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(37[14:21])
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(71[8:15])
    wire [2:0]r_Bit_Index;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(40[17:28])
    
    wire n13374, UartClk_2_enable_18, n13287, n13286, UartClk_2_enable_3;
    wire [2:0]r_SM_Main;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(43[17:26])
    
    wire n3, r_Rx_DV_last, r_Rx_DV, r_Rx_Data_R, r_Rx_Data;
    wire [7:0]r_Rx_Byte;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(41[17:26])
    
    wire UartClk_2_enable_1, r_Rx_DV_N_2484, UartClk_2_enable_25, n12821, 
        n12511, n13387, n1, n12841;
    wire [2:0]n4;
    wire [2:0]n17;
    
    wire n9118, UartClk_2_enable_5, n11803, UartClk_2_enable_4, n12819;
    wire [2:0]r_SM_Main_2__N_2418;
    
    wire n9085, n12796;
    wire [15:0]r_Clock_Count;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(39[18:31])
    
    wire n13414, UartClk_2_enable_23, n8374;
    wire [15:0]n69;
    
    wire n13061, n13063, n13055, n13059, n13073, n12406, n12405, 
        n12404, n12403, n12402, n12401, n12400, n12399, n13338, 
        n13379, n13378, n13386, UartClk_2_enable_26, n13410, n13409, 
        n13413, n13412, UartClk_2_enable_28, UartClk_2_enable_27, UartClk_2_enable_11, 
        n8372, r_Rx_DV_last_N_2483, n13377, n13079, n24, n13014, 
        n12822;
    
    LUT4 i5683_2_lut_3_lut_4_lut (.A(r_Bit_Index[1]), .B(n13374), .C(r_Bit_Index[0]), 
         .D(r_Bit_Index[2]), .Z(UartClk_2_enable_18)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(112[17:39])
    defparam i5683_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 n13287_bdd_4_lut (.A(n13287), .B(n13286), .C(o_Rx_Byte_c_2), 
         .D(n8225), .Z(n2795)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n13287_bdd_4_lut.init = 16'hca00;
    LUT4 i5716_2_lut_3_lut_4_lut (.A(r_Bit_Index[1]), .B(n13374), .C(r_Bit_Index[0]), 
         .D(r_Bit_Index[2]), .Z(UartClk_2_enable_3)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(112[17:39])
    defparam i5716_2_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 i5743_4_lut_4_lut_rep_113 (.A(o_Rx_Byte_c_4), .B(n13291), .C(n8225), 
         .D(n12970), .Z(n13523)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B (C)+!B !((D)+!C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam i5743_4_lut_4_lut_rep_113.init = 16'h40f0;
    FD1S3IX r_SM_Main_i0 (.D(n3), .CK(UartClk[2]), .CD(r_SM_Main[2]), 
            .Q(r_SM_Main[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_SM_Main_i0.GSR = "ENABLED";
    FD1S3AX r_Rx_DV_last_60 (.D(r_Rx_DV), .CK(osc_clk), .Q(r_Rx_DV_last)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(47[11] 52[8])
    defparam r_Rx_DV_last_60.GSR = "ENABLED";
    FD1S3AY r_Rx_Data_R_61 (.D(i_Rx_Serial_c), .CK(UartClk[2]), .Q(r_Rx_Data_R)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(57[12] 61[8])
    defparam r_Rx_Data_R_61.GSR = "ENABLED";
    FD1S3AY r_Rx_Data_62 (.D(r_Rx_Data_R), .CK(UartClk[2]), .Q(r_Rx_Data)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(57[12] 61[8])
    defparam r_Rx_Data_62.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i4 (.D(r_Rx_Data), .SP(UartClk_2_enable_1), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Rx_Byte_i4.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i1 (.D(r_Rx_Byte[0]), .SP(r_Rx_DV_N_2484), .CK(UartClk[2]), 
            .Q(o_Rx_Byte_c_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam o_Rx_Byte_i1.GSR = "ENABLED";
    FD1P3AX r_Bit_Index_i0 (.D(n12821), .SP(UartClk_2_enable_25), .CK(UartClk[2]), 
            .Q(r_Bit_Index[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Bit_Index_i0.GSR = "ENABLED";
    LUT4 r_SM_Main_2__I_0_69_Mux_0_i1_3_lut_4_lut_4_lut (.A(r_Rx_Data), .B(r_SM_Main[0]), 
         .C(n12511), .D(n13387), .Z(n1)) /* synthesis lut_function=(A (B (C+!(D)))+!A ((C+!(D))+!B)) */ ;
    defparam r_SM_Main_2__I_0_69_Mux_0_i1_3_lut_4_lut_4_lut.init = 16'hd1dd;
    LUT4 i5743_4_lut_4_lut_rep_114 (.A(o_Rx_Byte_c_4), .B(n13291), .C(n8225), 
         .D(n12970), .Z(osc_clk_enable_1447)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B (C)+!B !((D)+!C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam i5743_4_lut_4_lut_rep_114.init = 16'h40f0;
    LUT4 i2874_2_lut_2_lut (.A(o_Rx_Byte_c_4), .B(n2795), .Z(n3614)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam i2874_2_lut_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_2_lut (.A(o_Rx_Byte_c_4), .B(o_Rx_Byte_c_3), .Z(n6)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam i1_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_rep_69_2_lut (.A(o_Rx_Byte_c_4), .B(n12803), .Z(n13380)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam i1_2_lut_rep_69_2_lut.init = 16'h4444;
    LUT4 mux_743_i22_3_lut_3_lut (.A(o_Rx_Byte_c_4), .B(n2795), .C(o_Rx_Byte_c_2), 
         .Z(n3628)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam mux_743_i22_3_lut_3_lut.init = 16'h7474;
    LUT4 i5743_4_lut_4_lut (.A(o_Rx_Byte_c_4), .B(n13291), .C(n8225), 
         .D(n12970), .Z(osc_clk_enable_1457)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B (C)+!B !((D)+!C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam i5743_4_lut_4_lut.init = 16'h40f0;
    LUT4 i1_2_lut (.A(r_Bit_Index[0]), .B(r_Bit_Index[2]), .Z(n12841)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(112[17:39])
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 n2632_bdd_4_lut_5756_4_lut (.A(o_Rx_Byte_c_4), .B(o_Rx_Byte_c_3), 
         .C(n7349), .D(o_Rx_Byte_c_0), .Z(n13286)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam n2632_bdd_4_lut_5756_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_rep_74_2_lut (.A(o_Rx_Byte_c_4), .B(n7349), .Z(n13385)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam i1_2_lut_rep_74_2_lut.init = 16'h4444;
    LUT4 mux_318_i4_3_lut_4_lut_4_lut (.A(o_Rx_Byte_c_3), .B(n2608), .C(n1132), 
         .D(n13383), .Z(n2339)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[16:25])
    defparam mux_318_i4_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 n2632_bdd_4_lut_5779_4_lut (.A(o_Rx_Byte_c_3), .B(n7349), .C(o_Rx_Byte_c_4), 
         .D(o_Rx_Byte_c_0), .Z(n13287)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[16:25])
    defparam n2632_bdd_4_lut_5779_4_lut.init = 16'h0010;
    FD1S3AX UartClk_1000_1022__i0 (.D(n17[0]), .CK(osc_clk), .Q(n4[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(49[15:29])
    defparam UartClk_1000_1022__i0.GSR = "ENABLED";
    LUT4 i2965_2_lut_2_lut (.A(o_Rx_Byte_c_3), .B(n1030), .Z(n2364)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[16:25])
    defparam i2965_2_lut_2_lut.init = 16'hdddd;
    LUT4 i3032_2_lut_2_lut (.A(o_Rx_Byte_c_3), .B(n1018), .Z(n2486)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[16:25])
    defparam i3032_2_lut_2_lut.init = 16'hdddd;
    PFUMX r_SM_Main_2__I_0_69_Mux_0_i3 (.BLUT(n1), .ALUT(n9118), .C0(r_SM_Main[1]), 
          .Z(n3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;
    LUT4 n12931_bdd_4_lut_4_lut (.A(o_Rx_Byte_c_3), .B(n7349), .C(n12919), 
         .D(n12931), .Z(n13372)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[16:25])
    defparam n12931_bdd_4_lut_4_lut.init = 16'h5140;
    LUT4 i1_3_lut_4_lut_3_lut (.A(o_Rx_Byte_c_3), .B(n1034), .C(n13381), 
         .Z(n30)) /* synthesis lut_function=(A (B)+!A !(C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[16:25])
    defparam i1_3_lut_4_lut_3_lut.init = 16'h8d8d;
    LUT4 i1940_3_lut_4_lut_4_lut_4_lut (.A(o_Rx_Byte_c_3), .B(n12803), .C(n13381), 
         .D(o_Rx_Byte_c_4), .Z(n7970)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[16:25])
    defparam i1940_3_lut_4_lut_4_lut_4_lut.init = 16'h5054;
    LUT4 i1_2_lut_rep_65_3_lut_3_lut (.A(o_Rx_Byte_c_3), .B(n12803), .C(o_Rx_Byte_c_4), 
         .Z(n13376)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[16:25])
    defparam i1_2_lut_rep_65_3_lut_3_lut.init = 16'h4040;
    LUT4 i352_2_lut_rep_64_3_lut_3_lut_3_lut (.A(o_Rx_Byte_c_3), .B(n12803), 
         .C(o_Rx_Byte_c_4), .Z(n13375)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[16:25])
    defparam i352_2_lut_rep_64_3_lut_3_lut_3_lut.init = 16'h0404;
    LUT4 i1_3_lut_4_lut_3_lut_adj_44 (.A(o_Rx_Byte_c_3), .B(n1052), .C(n13381), 
         .Z(n28)) /* synthesis lut_function=(A (B)+!A !(C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[16:25])
    defparam i1_3_lut_4_lut_3_lut_adj_44.init = 16'h8d8d;
    LUT4 i3023_2_lut_2_lut (.A(o_Rx_Byte_c_3), .B(n1045), .Z(n2513)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[16:25])
    defparam i3023_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_3_lut_4_lut_3_lut_adj_45 (.A(o_Rx_Byte_c_3), .B(n1059), .C(n13381), 
         .Z(n29)) /* synthesis lut_function=(A (B)+!A !(C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[16:25])
    defparam i1_3_lut_4_lut_3_lut_adj_45.init = 16'h8d8d;
    LUT4 i1_4_lut_4_lut (.A(o_Rx_Byte_c_3), .B(o_Rx_Byte_c_2), .C(n13380), 
         .D(n13381), .Z(n2608)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[16:25])
    defparam i1_4_lut_4_lut.init = 16'h0400;
    FD1P3AX r_Rx_Byte_i3 (.D(r_Rx_Data), .SP(UartClk_2_enable_3), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Rx_Byte_i3.GSR = "ENABLED";
    LUT4 i5711_2_lut_3_lut_4_lut (.A(r_Bit_Index[1]), .B(n13374), .C(r_Bit_Index[0]), 
         .D(r_Bit_Index[2]), .Z(UartClk_2_enable_5)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(112[17:39])
    defparam i5711_2_lut_3_lut_4_lut.init = 16'h0010;
    CCU2D UartClk_1000_1022_add_4_3 (.A0(n4[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(UartClk[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11803), .S0(n17[1]), .S1(n17[2]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(49[15:29])
    defparam UartClk_1000_1022_add_4_3.INIT0 = 16'hfaaa;
    defparam UartClk_1000_1022_add_4_3.INIT1 = 16'hfaaa;
    defparam UartClk_1000_1022_add_4_3.INJECT1_0 = "NO";
    defparam UartClk_1000_1022_add_4_3.INJECT1_1 = "NO";
    CCU2D UartClk_1000_1022_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n4[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n11803), .S1(n17[0]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(49[15:29])
    defparam UartClk_1000_1022_add_4_1.INIT0 = 16'hF000;
    defparam UartClk_1000_1022_add_4_1.INIT1 = 16'h0555;
    defparam UartClk_1000_1022_add_4_1.INJECT1_0 = "NO";
    defparam UartClk_1000_1022_add_4_1.INJECT1_1 = "NO";
    FD1P3AX r_Rx_Byte_i2 (.D(r_Rx_Data), .SP(UartClk_2_enable_4), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Rx_Byte_i2.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i1 (.D(r_Rx_Data), .SP(UartClk_2_enable_5), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Rx_Byte_i1.GSR = "ENABLED";
    FD1S3IX r_SM_Main_i2 (.D(r_SM_Main_2__N_2418[2]), .CK(UartClk[2]), .CD(n12819), 
            .Q(r_SM_Main[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_SM_Main_i2.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(n9085), .B(n12796), .C(r_Clock_Count[6]), .D(r_Clock_Count[5]), 
         .Z(r_SM_Main_2__N_2418[2])) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(83[17:52])
    defparam i1_4_lut.init = 16'hfcec;
    FD1S3IX r_SM_Main_i1 (.D(n13414), .CK(UartClk[2]), .CD(r_SM_Main[2]), 
            .Q(r_SM_Main[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_SM_Main_i1.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i2 (.D(r_Rx_Byte[1]), .SP(r_Rx_DV_N_2484), .CK(UartClk[2]), 
            .Q(n7349)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam o_Rx_Byte_i2.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1002__i0 (.D(n69[0]), .SP(UartClk_2_enable_23), 
            .CD(n8374), .CK(UartClk[2]), .Q(r_Clock_Count[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002__i0.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i3 (.D(r_Rx_Byte[2]), .SP(r_Rx_DV_N_2484), .CK(UartClk[2]), 
            .Q(o_Rx_Byte_c_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam o_Rx_Byte_i3.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i4 (.D(r_Rx_Byte[3]), .SP(r_Rx_DV_N_2484), .CK(UartClk[2]), 
            .Q(o_Rx_Byte_c_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam o_Rx_Byte_i4.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i5 (.D(r_Rx_Byte[4]), .SP(r_Rx_DV_N_2484), .CK(UartClk[2]), 
            .Q(o_Rx_Byte_c_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam o_Rx_Byte_i5.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i6 (.D(r_Rx_Byte[5]), .SP(r_Rx_DV_N_2484), .CK(UartClk[2]), 
            .Q(o_Rx_Byte_c_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam o_Rx_Byte_i6.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i7 (.D(r_Rx_Byte[6]), .SP(r_Rx_DV_N_2484), .CK(UartClk[2]), 
            .Q(o_Rx_Byte_c_6)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam o_Rx_Byte_i7.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i8 (.D(r_Rx_Byte[7]), .SP(r_Rx_DV_N_2484), .CK(UartClk[2]), 
            .Q(o_Rx_Byte_c_7)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam o_Rx_Byte_i8.GSR = "ENABLED";
    LUT4 i3055_4_lut (.A(r_Clock_Count[1]), .B(r_Clock_Count[4]), .C(r_Clock_Count[3]), 
         .D(r_Clock_Count[2]), .Z(n9085)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i3055_4_lut.init = 16'hc8c0;
    FD1S3AX UartClk_1000_1022__i1 (.D(n17[1]), .CK(osc_clk), .Q(n4[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(49[15:29])
    defparam UartClk_1000_1022__i1.GSR = "ENABLED";
    FD1S3AX UartClk_1000_1022__i2 (.D(n17[2]), .CK(osc_clk), .Q(UartClk[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(49[15:29])
    defparam UartClk_1000_1022__i2.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1002__i15 (.D(n69[15]), .SP(UartClk_2_enable_23), 
            .CD(n8374), .CK(UartClk[2]), .Q(r_Clock_Count[15])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002__i15.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_46 (.A(n13061), .B(n13063), .C(n13055), .D(n13059), 
         .Z(n12796)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(83[17:52])
    defparam i1_4_lut_adj_46.init = 16'hfffe;
    LUT4 i1_2_lut_adj_47 (.A(r_Clock_Count[7]), .B(r_Clock_Count[10]), .Z(n13061)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(83[17:52])
    defparam i1_2_lut_adj_47.init = 16'heeee;
    LUT4 i1_4_lut_adj_48 (.A(r_Clock_Count[1]), .B(n12796), .C(n13073), 
         .D(r_Clock_Count[6]), .Z(n12511)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(83[17:52])
    defparam i1_4_lut_adj_48.init = 16'hfffd;
    FD1P3IX r_Clock_Count_1002__i14 (.D(n69[14]), .SP(UartClk_2_enable_23), 
            .CD(n8374), .CK(UartClk[2]), .Q(r_Clock_Count[14])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002__i14.GSR = "ENABLED";
    CCU2D r_Clock_Count_1002_add_4_17 (.A0(r_Clock_Count[15]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12406), .S0(n69[15]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002_add_4_17.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_1002_add_4_17.INIT1 = 16'h0000;
    defparam r_Clock_Count_1002_add_4_17.INJECT1_0 = "NO";
    defparam r_Clock_Count_1002_add_4_17.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_1002_add_4_15 (.A0(r_Clock_Count[13]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[14]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12405), .COUT(n12406), .S0(n69[13]), 
          .S1(n69[14]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002_add_4_15.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_1002_add_4_15.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_1002_add_4_15.INJECT1_0 = "NO";
    defparam r_Clock_Count_1002_add_4_15.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_1002_add_4_13 (.A0(r_Clock_Count[11]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[12]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12404), .COUT(n12405), .S0(n69[11]), 
          .S1(n69[12]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002_add_4_13.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_1002_add_4_13.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_1002_add_4_13.INJECT1_0 = "NO";
    defparam r_Clock_Count_1002_add_4_13.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_1002_add_4_11 (.A0(r_Clock_Count[9]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[10]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12403), .COUT(n12404), .S0(n69[9]), 
          .S1(n69[10]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002_add_4_11.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_1002_add_4_11.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_1002_add_4_11.INJECT1_0 = "NO";
    defparam r_Clock_Count_1002_add_4_11.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_1002_add_4_9 (.A0(r_Clock_Count[7]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[8]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12402), .COUT(n12403), .S0(n69[7]), 
          .S1(n69[8]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002_add_4_9.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_1002_add_4_9.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_1002_add_4_9.INJECT1_0 = "NO";
    defparam r_Clock_Count_1002_add_4_9.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_1002_add_4_7 (.A0(r_Clock_Count[5]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[6]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12401), .COUT(n12402), .S0(n69[5]), 
          .S1(n69[6]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002_add_4_7.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_1002_add_4_7.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_1002_add_4_7.INJECT1_0 = "NO";
    defparam r_Clock_Count_1002_add_4_7.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_1002_add_4_5 (.A0(r_Clock_Count[3]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[4]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12400), .COUT(n12401), .S0(n69[3]), 
          .S1(n69[4]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002_add_4_5.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_1002_add_4_5.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_1002_add_4_5.INJECT1_0 = "NO";
    defparam r_Clock_Count_1002_add_4_5.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_1002_add_4_3 (.A0(r_Clock_Count[1]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[2]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12399), .COUT(n12400), .S0(n69[1]), 
          .S1(n69[2]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002_add_4_3.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_1002_add_4_3.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_1002_add_4_3.INJECT1_0 = "NO";
    defparam r_Clock_Count_1002_add_4_3.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_1002_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(r_Clock_Count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n12399), .S1(n69[0]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002_add_4_1.INIT0 = 16'hF000;
    defparam r_Clock_Count_1002_add_4_1.INIT1 = 16'h0555;
    defparam r_Clock_Count_1002_add_4_1.INJECT1_0 = "NO";
    defparam r_Clock_Count_1002_add_4_1.INJECT1_1 = "NO";
    LUT4 i1_3_lut (.A(r_Clock_Count[13]), .B(r_Clock_Count[8]), .C(r_Clock_Count[15]), 
         .Z(n13063)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(83[17:52])
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_adj_49 (.A(r_Clock_Count[14]), .B(r_Clock_Count[11]), 
         .Z(n13055)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(83[17:52])
    defparam i1_2_lut_adj_49.init = 16'heeee;
    LUT4 i1_2_lut_adj_50 (.A(r_Clock_Count[9]), .B(r_Clock_Count[12]), .Z(n13059)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(83[17:52])
    defparam i1_2_lut_adj_50.init = 16'heeee;
    LUT4 i1_2_lut_adj_51 (.A(r_Clock_Count[2]), .B(r_Clock_Count[4]), .Z(n13073)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(83[17:52])
    defparam i1_2_lut_adj_51.init = 16'heeee;
    LUT4 i5714_2_lut_3_lut_4_lut (.A(r_Bit_Index[1]), .B(n13374), .C(r_Bit_Index[0]), 
         .D(r_Bit_Index[2]), .Z(UartClk_2_enable_4)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(112[17:39])
    defparam i5714_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i5734_4_lut (.A(n13523), .B(o_Rx_Byte_c_3), .C(n9000), .D(n13383), 
         .Z(osc_clk_enable_128)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))) */ ;
    defparam i5734_4_lut.init = 16'ha0a2;
    LUT4 r_Bit_Index_2__bdd_3_lut (.A(r_Bit_Index[2]), .B(r_Bit_Index[1]), 
         .C(r_Bit_Index[0]), .Z(n13338)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;
    defparam r_Bit_Index_2__bdd_3_lut.init = 16'h6a6a;
    LUT4 i1_3_lut_rep_68 (.A(r_SM_Main[0]), .B(r_SM_Main_2__N_2418[2]), 
         .C(r_SM_Main[1]), .Z(n13379)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_3_lut_rep_68.init = 16'h4040;
    LUT4 i1_2_lut_4_lut (.A(r_SM_Main[0]), .B(r_SM_Main_2__N_2418[2]), .C(r_SM_Main[1]), 
         .D(r_Bit_Index[0]), .Z(n12821)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0040;
    LUT4 i1_4_lut_adj_52 (.A(r_SM_Main[0]), .B(r_SM_Main_2__N_2418[2]), 
         .C(r_SM_Main[2]), .D(r_SM_Main[1]), .Z(UartClk_2_enable_25)) /* synthesis lut_function=(!(A+(B (C)+!B (C+(D))))) */ ;
    defparam i1_4_lut_adj_52.init = 16'h0405;
    LUT4 i5726_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n13378), .C(n13386), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_26)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(112[17:39])
    defparam i5726_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i5787_then_4_lut (.A(n1128), .B(n1067), .C(o_Rx_Byte_c_3), .D(o_Rx_Byte_c_4), 
         .Z(n13410)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;
    defparam i5787_then_4_lut.init = 16'hcacf;
    LUT4 i5787_else_4_lut (.A(n1067), .B(o_Rx_Byte_c_3), .C(n13381), .Z(n13409)) /* synthesis lut_function=(A (B+!(C))+!A !(B+(C))) */ ;
    defparam i5787_else_4_lut.init = 16'h8b8b;
    LUT4 r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_then_3_lut (.A(r_SM_Main[0]), 
         .B(r_SM_Main_2__N_2418[2]), .C(r_SM_Main[1]), .Z(n13413)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(67[7] 159[14])
    defparam r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_then_3_lut.init = 16'h7070;
    LUT4 r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_else_3_lut (.A(r_SM_Main[0]), 
         .B(r_SM_Main_2__N_2418[2]), .C(r_SM_Main[1]), .D(r_Rx_Data), 
         .Z(n13412)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A !(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(67[7] 159[14])
    defparam r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_else_3_lut.init = 16'h707a;
    LUT4 i3086_3_lut_4_lut (.A(r_Bit_Index[1]), .B(n13386), .C(r_SM_Main[0]), 
         .D(r_SM_Main_2__N_2418[2]), .Z(n9118)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((D)+!C))) */ ;
    defparam i3086_3_lut_4_lut.init = 16'h08f0;
    LUT4 i5721_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n13378), .C(n13386), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_28)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(112[17:39])
    defparam i5721_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i5724_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n13378), .C(n12841), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_27)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(112[17:39])
    defparam i5724_2_lut_3_lut_4_lut.init = 16'h0100;
    FD1P3IX r_Clock_Count_1002__i13 (.D(n69[13]), .SP(UartClk_2_enable_23), 
            .CD(n8374), .CK(UartClk[2]), .Q(r_Clock_Count[13])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002__i13.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1002__i12 (.D(n69[12]), .SP(UartClk_2_enable_23), 
            .CD(n8374), .CK(UartClk[2]), .Q(r_Clock_Count[12])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002__i12.GSR = "ENABLED";
    FD1P3AX r_Rx_DV_64 (.D(r_Rx_DV_N_2484), .SP(UartClk_2_enable_11), .CK(UartClk[2]), 
            .Q(r_Rx_DV)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Rx_DV_64.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1002__i11 (.D(n69[11]), .SP(UartClk_2_enable_23), 
            .CD(n8374), .CK(UartClk[2]), .Q(r_Clock_Count[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002__i11.GSR = "ENABLED";
    LUT4 i5709_2_lut_3_lut (.A(r_SM_Main[1]), .B(r_SM_Main[2]), .C(r_SM_Main[0]), 
         .Z(n12819)) /* synthesis lut_function=((B+!(C))+!A) */ ;
    defparam i5709_2_lut_3_lut.init = 16'hdfdf;
    FD1P3IX r_Clock_Count_1002__i10 (.D(n69[10]), .SP(UartClk_2_enable_23), 
            .CD(n8374), .CK(UartClk[2]), .Q(r_Clock_Count[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002__i10.GSR = "ENABLED";
    LUT4 i3089_3_lut_4_lut (.A(n8225), .B(n13384), .C(o_Rx_Byte_c_3), 
         .D(n1062), .Z(n2530)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(47[11] 52[8])
    defparam i3089_3_lut_4_lut.init = 16'hf808;
    FD1S3IX o_Rx_DV_59 (.D(r_Rx_DV_last_N_2483), .CK(osc_clk), .CD(n8372), 
            .Q(o_Rx_DV_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(47[11] 52[8])
    defparam o_Rx_DV_59.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1002__i9 (.D(n69[9]), .SP(UartClk_2_enable_23), 
            .CD(n8374), .CK(UartClk[2]), .Q(r_Clock_Count[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002__i9.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1002__i8 (.D(n69[8]), .SP(UartClk_2_enable_23), 
            .CD(n8374), .CK(UartClk[2]), .Q(r_Clock_Count[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002__i8.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1002__i7 (.D(n69[7]), .SP(UartClk_2_enable_23), 
            .CD(n8374), .CK(UartClk[2]), .Q(r_Clock_Count[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002__i7.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1002__i6 (.D(n69[6]), .SP(UartClk_2_enable_23), 
            .CD(n8374), .CK(UartClk[2]), .Q(r_Clock_Count[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002__i6.GSR = "ENABLED";
    LUT4 i5719_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n13378), .C(n12841), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_1)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(112[17:39])
    defparam i5719_2_lut_3_lut_4_lut.init = 16'h0001;
    FD1P3AX r_Rx_Byte_i0 (.D(r_Rx_Data), .SP(UartClk_2_enable_18), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Rx_Byte_i0.GSR = "ENABLED";
    LUT4 i21_4_lut_4_lut (.A(r_SM_Main[1]), .B(r_SM_Main[2]), .C(r_SM_Main[0]), 
         .D(r_SM_Main_2__N_2418[2]), .Z(UartClk_2_enable_11)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (C))) */ ;
    defparam i21_4_lut_4_lut.init = 16'h2505;
    LUT4 i1_2_lut_rep_75 (.A(r_Bit_Index[2]), .B(r_Bit_Index[0]), .Z(n13386)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_75.init = 16'h8888;
    LUT4 i1_3_lut_rep_76 (.A(r_Clock_Count[3]), .B(r_Clock_Count[5]), .C(r_Clock_Count[0]), 
         .Z(n13387)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_rep_76.init = 16'h8080;
    LUT4 i1_2_lut_rep_66_4_lut (.A(r_Clock_Count[3]), .B(r_Clock_Count[5]), 
         .C(r_Clock_Count[0]), .D(n12511), .Z(n13377)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_2_lut_rep_66_4_lut.init = 16'hff7f;
    LUT4 i1_2_lut_rep_67_3_lut (.A(r_SM_Main[2]), .B(r_SM_Main[1]), .C(r_SM_Main_2__N_2418[2]), 
         .Z(n13378)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i1_2_lut_rep_67_3_lut.init = 16'hbfbf;
    LUT4 i5746_4_lut (.A(r_SM_Main[2]), .B(r_SM_Main[1]), .C(n13377), 
         .D(n13079), .Z(UartClk_2_enable_23)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(67[7] 159[14])
    defparam i5746_4_lut.init = 16'h5455;
    LUT4 i1_2_lut_adj_53 (.A(r_Rx_Data), .B(r_SM_Main[0]), .Z(n13079)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_53.init = 16'h8888;
    LUT4 i1_2_lut_rep_63_3_lut_4_lut (.A(r_SM_Main[2]), .B(r_SM_Main[1]), 
         .C(r_SM_Main[0]), .D(r_SM_Main_2__N_2418[2]), .Z(n13374)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;
    defparam i1_2_lut_rep_63_3_lut_4_lut.init = 16'hfbff;
    LUT4 i1_4_lut_adj_54 (.A(r_SM_Main[2]), .B(n24), .C(r_SM_Main_2__N_2418[2]), 
         .D(r_SM_Main[1]), .Z(n8374)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;
    defparam i1_4_lut_adj_54.init = 16'h5044;
    FD1P3IX r_Clock_Count_1002__i5 (.D(n69[5]), .SP(UartClk_2_enable_23), 
            .CD(n8374), .CK(UartClk[2]), .Q(r_Clock_Count[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002__i5.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1002__i4 (.D(n69[4]), .SP(UartClk_2_enable_23), 
            .CD(n8374), .CK(UartClk[2]), .Q(r_Clock_Count[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002__i4.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1002__i3 (.D(n69[3]), .SP(UartClk_2_enable_23), 
            .CD(n8374), .CK(UartClk[2]), .Q(r_Clock_Count[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002__i3.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1002__i2 (.D(n69[2]), .SP(UartClk_2_enable_23), 
            .CD(n8374), .CK(UartClk[2]), .Q(r_Clock_Count[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002__i2.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1002__i1 (.D(n69[1]), .SP(UartClk_2_enable_23), 
            .CD(n8374), .CK(UartClk[2]), .Q(r_Clock_Count[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_1002__i1.GSR = "ENABLED";
    FD1P3AX r_Bit_Index_i2 (.D(n13014), .SP(UartClk_2_enable_25), .CK(UartClk[2]), 
            .Q(r_Bit_Index[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Bit_Index_i2.GSR = "ENABLED";
    FD1P3AX r_Bit_Index_i1 (.D(n12822), .SP(UartClk_2_enable_25), .CK(UartClk[2]), 
            .Q(r_Bit_Index[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Bit_Index_i1.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i7 (.D(r_Rx_Data), .SP(UartClk_2_enable_26), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Rx_Byte_i7.GSR = "ENABLED";
    LUT4 i2337_1_lut (.A(r_Rx_DV), .Z(n8372)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam i2337_1_lut.init = 16'h5555;
    LUT4 r_Rx_DV_last_I_0_1_lut (.A(r_Rx_DV_last), .Z(r_Rx_DV_last_N_2483)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(50[30:43])
    defparam r_Rx_DV_last_I_0_1_lut.init = 16'h5555;
    LUT4 i4_4_lut (.A(n13338), .B(r_SM_Main[0]), .C(r_SM_Main[1]), .D(r_SM_Main_2__N_2418[2]), 
         .Z(n13014)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i4_4_lut.init = 16'h2000;
    LUT4 i1_3_lut_adj_55 (.A(r_Bit_Index[0]), .B(n13379), .C(r_Bit_Index[1]), 
         .Z(n12822)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam i1_3_lut_adj_55.init = 16'h4848;
    FD1P3AX r_Rx_Byte_i6 (.D(r_Rx_Data), .SP(UartClk_2_enable_27), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Rx_Byte_i6.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i5 (.D(r_Rx_Data), .SP(UartClk_2_enable_28), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=217, LSE_RLINE=222 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Rx_Byte_i5.GSR = "ENABLED";
    PFUMX i5806 (.BLUT(n13412), .ALUT(n13413), .C0(n13377), .Z(n13414));
    LUT4 i5739_2_lut_3_lut_4_lut (.A(r_SM_Main[2]), .B(r_SM_Main[1]), .C(r_SM_Main[0]), 
         .D(r_SM_Main_2__N_2418[2]), .Z(r_Rx_DV_N_2484)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i5739_2_lut_3_lut_4_lut.init = 16'h4000;
    PFUMX i5804 (.BLUT(n13409), .ALUT(n13410), .C0(n12803), .Z(n13411));
    LUT4 i1_4_lut_4_lut_adj_56 (.A(r_Rx_Data), .B(n13387), .C(n12511), 
         .D(r_SM_Main[0]), .Z(n24)) /* synthesis lut_function=(!(A (D)+!A (B (C (D))+!B (D)))) */ ;
    defparam i1_4_lut_4_lut_adj_56.init = 16'h04ff;
    
endmodule
//
// Verilog Description of module SinCos
//

module SinCos (osc_clk, VCC_net, GND_net, \phase_accum[57] , \phase_accum[58] , 
            \phase_accum[59] , \phase_accum[60] , \phase_accum[61] , \phase_accum[62] , 
            \phase_accum[63] , \LOSine[1] , \LOSine[2] , \LOSine[3] , 
            \LOSine[4] , \LOSine[5] , \LOSine[6] , \LOSine[7] , \LOSine[8] , 
            \LOSine[9] , \LOSine[10] , \LOSine[11] , \LOSine[12] , \LOCosine[1] , 
            \LOCosine[2] , \LOCosine[3] , \LOCosine[4] , \LOCosine[5] , 
            \LOCosine[6] , \LOCosine[7] , \LOCosine[8] , \LOCosine[9] , 
            \LOCosine[10] , \LOCosine[11] , \LOCosine[12] , \phase_accum[56] ) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input osc_clk;
    input VCC_net;
    input GND_net;
    input \phase_accum[57] ;
    input \phase_accum[58] ;
    input \phase_accum[59] ;
    input \phase_accum[60] ;
    input \phase_accum[61] ;
    input \phase_accum[62] ;
    input \phase_accum[63] ;
    output \LOSine[1] ;
    output \LOSine[2] ;
    output \LOSine[3] ;
    output \LOSine[4] ;
    output \LOSine[5] ;
    output \LOSine[6] ;
    output \LOSine[7] ;
    output \LOSine[8] ;
    output \LOSine[9] ;
    output \LOSine[10] ;
    output \LOSine[11] ;
    output \LOSine[12] ;
    output \LOCosine[1] ;
    output \LOCosine[2] ;
    output \LOCosine[3] ;
    output \LOCosine[4] ;
    output \LOCosine[5] ;
    output \LOCosine[6] ;
    output \LOCosine[7] ;
    output \LOCosine[8] ;
    output \LOCosine[9] ;
    output \LOCosine[10] ;
    output \LOCosine[11] ;
    output \LOCosine[12] ;
    input \phase_accum[56] ;
    
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(71[8:15])
    
    wire rom_addr0_r_1, rom_addr0_r_1_inv, rom_addr0_r_2, rom_addr0_r_3, 
        rom_addr0_r_4, rom_addr0_r_5, mx_ctrl_r, mx_ctrl_r_1, rom_addr0_r, 
        rom_addr0_r_n, rom_addr0_r_6, rom_dout_11, rom_dout_11_ffin, 
        rom_dout_10, rom_dout_10_ffin, rom_dout_9, rom_dout_9_ffin, 
        rom_dout_8, rom_dout_8_ffin, rom_dout_7, rom_dout_7_ffin, rom_dout_6, 
        rom_dout_6_ffin, rom_dout_5, rom_dout_5_ffin, rom_dout_4, rom_dout_4_ffin, 
        rom_dout_3, rom_dout_3_ffin, rom_dout_2, rom_dout_2_ffin, rom_dout_1, 
        rom_dout_1_ffin, rom_dout, rom_dout_ffin, rom_dout_25, rom_dout_25_ffin, 
        rom_dout_24, rom_dout_24_ffin, rom_dout_23, rom_dout_23_ffin, 
        rom_dout_22, rom_dout_22_ffin, rom_dout_21, rom_dout_21_ffin, 
        rom_dout_20, rom_dout_20_ffin, rom_dout_19, rom_dout_19_ffin, 
        rom_dout_18, rom_dout_18_ffin, rom_dout_17, rom_dout_17_ffin, 
        rom_dout_16, rom_dout_16_ffin, rom_dout_15, rom_dout_15_ffin, 
        rom_dout_14, rom_dout_14_ffin, rom_dout_13, rom_dout_13_ffin, 
        cosromoutsel_i, cosromoutsel, sinromoutsel, sinout_pre_1, sinout_pre_2, 
        sinout_pre_3, sinout_pre_4, sinout_pre_5, sinout_pre_6, sinout_pre_7, 
        sinout_pre_8, sinout_pre_9, sinout_pre_10, sinout_pre_11, sinout_pre_12, 
        cosout_pre_1, cosout_pre_2, cosout_pre_3, cosout_pre_4, cosout_pre_5, 
        cosout_pre_6, cosout_pre_7, cosout_pre_8, cosout_pre_9, cosout_pre_10, 
        cosout_pre_11, cosout_pre_12, rom_addr0_r_inv, co0, rom_addr0_r_n_1, 
        rom_addr0_r_n_2, rom_addr0_r_2_inv, co1, rom_addr0_r_n_3, rom_addr0_r_n_4, 
        rom_addr0_r_3_inv, rom_addr0_r_4_inv, co2, rom_addr0_r_n_5, 
        rom_addr0_r_5_inv, rom_dout_12_ffin, rom_addr0_r_7, rom_addr0_r_8, 
        rom_addr0_r_9, rom_addr0_r_10, rom_addr0_r_11, rom_dout_s_n_1, 
        rom_dout_s_n_2, co0_1, rom_dout_1_inv, rom_dout_2_inv, co1_1, 
        rom_dout_s_n_3, rom_dout_s_n_4, rom_dout_3_inv, rom_dout_4_inv, 
        co2_1, rom_dout_s_n_5, rom_dout_s_n_6, rom_dout_5_inv, rom_dout_6_inv, 
        co3, rom_dout_s_n_7, rom_dout_s_n_8, rom_dout_7_inv, rom_dout_8_inv, 
        co4, rom_dout_s_n_9, rom_dout_s_n_10, rom_dout_9_inv, rom_dout_10_inv, 
        co5, rom_dout_s_n_11, rom_dout_s_n_12, rom_dout_11_inv, rom_dout_12_inv, 
        rom_dout_13_inv, co0_2, rom_dout_c_n_1, rom_dout_c_n_2, rom_dout_14_inv, 
        rom_dout_15_inv, co1_2, rom_dout_c_n_3, rom_dout_c_n_4, rom_dout_16_inv, 
        rom_dout_17_inv, co2_2, rom_dout_c_n_5, rom_dout_c_n_6, rom_dout_18_inv, 
        rom_dout_19_inv, co3_1, rom_dout_c_n_7, rom_dout_c_n_8, rom_dout_20_inv, 
        rom_dout_21_inv, co4_1, rom_dout_c_n_9, rom_dout_c_n_10, rom_dout_22_inv, 
        rom_dout_23_inv, co5_1, rom_dout_c_n_11, rom_dout_c_n_12, rom_dout_24_inv, 
        rom_dout_25_inv, rom_dout_12, rom_dout_inv, func_or_inet, lx_ne0, 
        lx_ne0_inv, out_sel_i, rom_dout_s_1, rom_dout_s_2, rom_dout_s_3, 
        rom_dout_s_4, rom_dout_s_5, rom_dout_s_6, rom_dout_s_7, rom_dout_s_8, 
        rom_dout_s_9, rom_dout_s_10, rom_dout_s_11, rom_dout_s_12, rom_dout_c_1, 
        rom_dout_c_2, rom_dout_c_3, rom_dout_c_4, rom_dout_c_5, rom_dout_c_6, 
        rom_dout_c_7, rom_dout_c_8, rom_dout_c_9, rom_dout_c_10, rom_dout_c_11, 
        rom_dout_c_12, out_sel;
    
    INV INV_29 (.A(rom_addr0_r_1), .Z(rom_addr0_r_1_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    FD1P3DX FF_61 (.D(\phase_accum[57] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(rom_addr0_r_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(312[13:88])
    defparam FF_61.GSR = "ENABLED";
    FD1P3DX FF_60 (.D(\phase_accum[58] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(rom_addr0_r_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(315[13:88])
    defparam FF_60.GSR = "ENABLED";
    FD1P3DX FF_59 (.D(\phase_accum[59] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(rom_addr0_r_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(318[13:88])
    defparam FF_59.GSR = "ENABLED";
    FD1P3DX FF_58 (.D(\phase_accum[60] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(rom_addr0_r_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(321[13:88])
    defparam FF_58.GSR = "ENABLED";
    FD1P3DX FF_57 (.D(\phase_accum[61] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(rom_addr0_r_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(324[13:88])
    defparam FF_57.GSR = "ENABLED";
    FD1P3DX FF_56 (.D(\phase_accum[62] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(mx_ctrl_r)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(327[13:84])
    defparam FF_56.GSR = "ENABLED";
    FD1P3DX FF_55 (.D(\phase_accum[63] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(mx_ctrl_r_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(330[13:86])
    defparam FF_55.GSR = "ENABLED";
    MUX21 muxb_57 (.D0(rom_addr0_r), .D1(rom_addr0_r_n), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    FD1P3DX FF_53 (.D(rom_dout_11_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(355[13] 356[25])
    defparam FF_53.GSR = "ENABLED";
    FD1P3DX FF_52 (.D(rom_dout_10_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(359[13] 360[25])
    defparam FF_52.GSR = "ENABLED";
    FD1P3DX FF_51 (.D(rom_dout_9_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(363[13] 364[24])
    defparam FF_51.GSR = "ENABLED";
    FD1P3DX FF_50 (.D(rom_dout_8_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(367[13] 368[24])
    defparam FF_50.GSR = "ENABLED";
    FD1P3DX FF_49 (.D(rom_dout_7_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(371[13] 372[24])
    defparam FF_49.GSR = "ENABLED";
    FD1P3DX FF_48 (.D(rom_dout_6_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(375[13] 376[24])
    defparam FF_48.GSR = "ENABLED";
    FD1P3DX FF_47 (.D(rom_dout_5_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(379[13] 380[24])
    defparam FF_47.GSR = "ENABLED";
    FD1P3DX FF_46 (.D(rom_dout_4_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(383[13] 384[24])
    defparam FF_46.GSR = "ENABLED";
    FD1P3DX FF_45 (.D(rom_dout_3_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(387[13] 388[24])
    defparam FF_45.GSR = "ENABLED";
    FD1P3DX FF_44 (.D(rom_dout_2_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(391[13] 392[24])
    defparam FF_44.GSR = "ENABLED";
    FD1P3DX FF_43 (.D(rom_dout_1_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(395[13] 396[24])
    defparam FF_43.GSR = "ENABLED";
    FD1P3DX FF_42 (.D(rom_dout_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(399[13] 400[22])
    defparam FF_42.GSR = "ENABLED";
    FD1P3DX FF_41 (.D(rom_dout_25_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_25)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(403[13] 404[25])
    defparam FF_41.GSR = "ENABLED";
    FD1P3DX FF_40 (.D(rom_dout_24_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_24)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(407[13] 408[25])
    defparam FF_40.GSR = "ENABLED";
    FD1P3DX FF_39 (.D(rom_dout_23_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_23)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(411[13] 412[25])
    defparam FF_39.GSR = "ENABLED";
    FD1P3DX FF_38 (.D(rom_dout_22_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_22)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(415[13] 416[25])
    defparam FF_38.GSR = "ENABLED";
    FD1P3DX FF_37 (.D(rom_dout_21_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(419[13] 420[25])
    defparam FF_37.GSR = "ENABLED";
    FD1P3DX FF_36 (.D(rom_dout_20_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(423[13] 424[25])
    defparam FF_36.GSR = "ENABLED";
    FD1P3DX FF_35 (.D(rom_dout_19_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(427[13] 428[25])
    defparam FF_35.GSR = "ENABLED";
    FD1P3DX FF_34 (.D(rom_dout_18_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(431[13] 432[25])
    defparam FF_34.GSR = "ENABLED";
    FD1P3DX FF_33 (.D(rom_dout_17_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(435[13] 436[25])
    defparam FF_33.GSR = "ENABLED";
    FD1P3DX FF_32 (.D(rom_dout_16_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(439[13] 440[25])
    defparam FF_32.GSR = "ENABLED";
    FD1P3DX FF_31 (.D(rom_dout_15_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(443[13] 444[25])
    defparam FF_31.GSR = "ENABLED";
    FD1P3DX FF_30 (.D(rom_dout_14_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(447[13] 448[25])
    defparam FF_30.GSR = "ENABLED";
    FD1P3DX FF_29 (.D(rom_dout_13_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(451[13] 452[25])
    defparam FF_29.GSR = "ENABLED";
    FD1P3DX FF_28 (.D(cosromoutsel_i), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(cosromoutsel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(455[13] 456[26])
    defparam FF_28.GSR = "ENABLED";
    FD1P3DX FF_27 (.D(mx_ctrl_r_1), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(sinromoutsel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(459[13] 460[26])
    defparam FF_27.GSR = "ENABLED";
    FD1P3DX FF_24 (.D(sinout_pre_1), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[1] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(599[13] 600[21])
    defparam FF_24.GSR = "ENABLED";
    FD1P3DX FF_23 (.D(sinout_pre_2), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[2] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(603[13] 604[21])
    defparam FF_23.GSR = "ENABLED";
    FD1P3DX FF_22 (.D(sinout_pre_3), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[3] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(607[13] 608[21])
    defparam FF_22.GSR = "ENABLED";
    FD1P3DX FF_21 (.D(sinout_pre_4), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[4] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(611[13] 612[21])
    defparam FF_21.GSR = "ENABLED";
    FD1P3DX FF_20 (.D(sinout_pre_5), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[5] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(615[13] 616[21])
    defparam FF_20.GSR = "ENABLED";
    FD1P3DX FF_19 (.D(sinout_pre_6), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[6] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(619[13] 620[21])
    defparam FF_19.GSR = "ENABLED";
    FD1P3DX FF_18 (.D(sinout_pre_7), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[7] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(623[13] 624[21])
    defparam FF_18.GSR = "ENABLED";
    FD1P3DX FF_17 (.D(sinout_pre_8), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[8] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(627[13] 628[21])
    defparam FF_17.GSR = "ENABLED";
    FD1P3DX FF_16 (.D(sinout_pre_9), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[9] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(631[13] 632[21])
    defparam FF_16.GSR = "ENABLED";
    FD1P3DX FF_15 (.D(sinout_pre_10), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[10] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(635[13] 636[22])
    defparam FF_15.GSR = "ENABLED";
    FD1P3DX FF_14 (.D(sinout_pre_11), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[11] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(639[13] 640[22])
    defparam FF_14.GSR = "ENABLED";
    FD1P3DX FF_13 (.D(sinout_pre_12), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[12] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(643[13] 644[22])
    defparam FF_13.GSR = "ENABLED";
    FD1P3DX FF_11 (.D(cosout_pre_1), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[1] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(650[13] 651[23])
    defparam FF_11.GSR = "ENABLED";
    FD1P3DX FF_10 (.D(cosout_pre_2), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[2] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(654[13] 655[23])
    defparam FF_10.GSR = "ENABLED";
    FD1P3DX FF_9 (.D(cosout_pre_3), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[3] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(658[13] 659[23])
    defparam FF_9.GSR = "ENABLED";
    FD1P3DX FF_8 (.D(cosout_pre_4), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[4] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(662[13] 663[23])
    defparam FF_8.GSR = "ENABLED";
    FD1P3DX FF_7 (.D(cosout_pre_5), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[5] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(666[13] 667[23])
    defparam FF_7.GSR = "ENABLED";
    FD1P3DX FF_6 (.D(cosout_pre_6), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[6] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(670[13] 671[23])
    defparam FF_6.GSR = "ENABLED";
    FD1P3DX FF_5 (.D(cosout_pre_7), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[7] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(674[13] 675[23])
    defparam FF_5.GSR = "ENABLED";
    FD1P3DX FF_4 (.D(cosout_pre_8), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[8] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(678[13] 679[23])
    defparam FF_4.GSR = "ENABLED";
    FD1P3DX FF_3 (.D(cosout_pre_9), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[9] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(682[13] 683[23])
    defparam FF_3.GSR = "ENABLED";
    FD1P3DX FF_2 (.D(cosout_pre_10), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[10] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(686[13] 687[24])
    defparam FF_2.GSR = "ENABLED";
    FD1P3DX FF_1 (.D(cosout_pre_11), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[11] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(690[13] 691[24])
    defparam FF_1.GSR = "ENABLED";
    FD1P3DX FF_0 (.D(cosout_pre_12), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[12] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(694[13] 695[24])
    defparam FF_0.GSR = "ENABLED";
    FADD2B neg_rom_addr0_r_n_0 (.A0(GND_net), .A1(rom_addr0_r_inv), .B0(GND_net), 
           .B1(VCC_net), .CI(GND_net), .COUT(co0), .S1(rom_addr0_r_n)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    FADD2B neg_rom_addr0_r_n_1 (.A0(rom_addr0_r_1_inv), .A1(rom_addr0_r_2_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co0), .COUT(co1), .S0(rom_addr0_r_n_1), 
           .S1(rom_addr0_r_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    FADD2B neg_rom_addr0_r_n_2 (.A0(rom_addr0_r_3_inv), .A1(rom_addr0_r_4_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co1), .COUT(co2), .S0(rom_addr0_r_n_3), 
           .S1(rom_addr0_r_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    FADD2B neg_rom_addr0_r_n_3 (.A0(rom_addr0_r_5_inv), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co2), .S0(rom_addr0_r_n_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    ROM64X1A triglut_1_0_25 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_12_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_25.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    FADD2B neg_rom_dout_s_n_1 (.A0(rom_dout_1_inv), .A1(rom_dout_2_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co0_1), .COUT(co1_1), .S0(rom_dout_s_n_1), 
           .S1(rom_dout_s_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    FADD2B neg_rom_dout_s_n_2 (.A0(rom_dout_3_inv), .A1(rom_dout_4_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co1_1), .COUT(co2_1), .S0(rom_dout_s_n_3), 
           .S1(rom_dout_s_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    FADD2B neg_rom_dout_s_n_3 (.A0(rom_dout_5_inv), .A1(rom_dout_6_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co2_1), .COUT(co3), .S0(rom_dout_s_n_5), 
           .S1(rom_dout_s_n_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    FADD2B neg_rom_dout_s_n_4 (.A0(rom_dout_7_inv), .A1(rom_dout_8_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co3), .COUT(co4), .S0(rom_dout_s_n_7), 
           .S1(rom_dout_s_n_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    FADD2B neg_rom_dout_s_n_5 (.A0(rom_dout_9_inv), .A1(rom_dout_10_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co4), .COUT(co5), .S0(rom_dout_s_n_9), 
           .S1(rom_dout_s_n_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    FADD2B neg_rom_dout_s_n_6 (.A0(rom_dout_11_inv), .A1(rom_dout_12_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co5), .S0(rom_dout_s_n_11), 
           .S1(rom_dout_s_n_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_30 (.A(rom_addr0_r_2), .Z(rom_addr0_r_2_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    FADD2B neg_rom_dout_c_n_0 (.A0(GND_net), .A1(rom_dout_13_inv), .B0(GND_net), 
           .B1(VCC_net), .CI(GND_net), .COUT(co0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    FADD2B neg_rom_dout_c_n_1 (.A0(rom_dout_14_inv), .A1(rom_dout_15_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co0_2), .COUT(co1_2), .S0(rom_dout_c_n_1), 
           .S1(rom_dout_c_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    FADD2B neg_rom_dout_c_n_2 (.A0(rom_dout_16_inv), .A1(rom_dout_17_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co1_2), .COUT(co2_2), .S0(rom_dout_c_n_3), 
           .S1(rom_dout_c_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    FADD2B neg_rom_dout_c_n_3 (.A0(rom_dout_18_inv), .A1(rom_dout_19_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co2_2), .COUT(co3_1), .S0(rom_dout_c_n_5), 
           .S1(rom_dout_c_n_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    FADD2B neg_rom_dout_c_n_4 (.A0(rom_dout_20_inv), .A1(rom_dout_21_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co3_1), .COUT(co4_1), .S0(rom_dout_c_n_7), 
           .S1(rom_dout_c_n_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    FADD2B neg_rom_dout_c_n_5 (.A0(rom_dout_22_inv), .A1(rom_dout_23_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co4_1), .COUT(co5_1), .S0(rom_dout_c_n_9), 
           .S1(rom_dout_c_n_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    FADD2B neg_rom_dout_c_n_6 (.A0(rom_dout_24_inv), .A1(rom_dout_25_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co5_1), .S0(rom_dout_c_n_11), 
           .S1(rom_dout_c_n_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_31 (.A(rom_addr0_r_3), .Z(rom_addr0_r_3_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_32 (.A(rom_addr0_r_4), .Z(rom_addr0_r_4_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_33 (.A(rom_addr0_r_5), .Z(rom_addr0_r_5_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_28 (.A(rom_addr0_r), .Z(rom_addr0_r_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    XOR2 XOR2_t1 (.A(mx_ctrl_r), .B(mx_ctrl_r_1), .Z(cosromoutsel_i)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(241[10:70])
    INV INV_27 (.A(rom_dout_12), .Z(rom_dout_12_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_26 (.A(rom_dout_11), .Z(rom_dout_11_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_25 (.A(rom_dout_10), .Z(rom_dout_10_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_24 (.A(rom_dout_9), .Z(rom_dout_9_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_23 (.A(rom_dout_8), .Z(rom_dout_8_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_22 (.A(rom_dout_7), .Z(rom_dout_7_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_21 (.A(rom_dout_6), .Z(rom_dout_6_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_20 (.A(rom_dout_5), .Z(rom_dout_5_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_19 (.A(rom_dout_4), .Z(rom_dout_4_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_18 (.A(rom_dout_3), .Z(rom_dout_3_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_17 (.A(rom_dout_2), .Z(rom_dout_2_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_16 (.A(rom_dout_1), .Z(rom_dout_1_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_15 (.A(rom_dout), .Z(rom_dout_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_14 (.A(rom_dout_25), .Z(rom_dout_25_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_13 (.A(rom_dout_24), .Z(rom_dout_24_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_12 (.A(rom_dout_23), .Z(rom_dout_23_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_11 (.A(rom_dout_22), .Z(rom_dout_22_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_10 (.A(rom_dout_21), .Z(rom_dout_21_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_9 (.A(rom_dout_20), .Z(rom_dout_20_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_8 (.A(rom_dout_19), .Z(rom_dout_19_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_7 (.A(rom_dout_18), .Z(rom_dout_18_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_6 (.A(rom_dout_17), .Z(rom_dout_17_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_5 (.A(rom_dout_16), .Z(rom_dout_16_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_4 (.A(rom_dout_15), .Z(rom_dout_15_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_3 (.A(rom_dout_14), .Z(rom_dout_14_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    INV INV_2 (.A(rom_dout_13), .Z(rom_dout_13_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    ROM16X1A LUT4_1 (.AD0(rom_addr0_r_9), .AD1(rom_addr0_r_8), .AD2(rom_addr0_r_7), 
            .AD3(rom_addr0_r_6), .DO0(func_or_inet)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam LUT4_1.initval = 16'b1111111111111110;
    ROM16X1A LUT4_0 (.AD0(GND_net), .AD1(rom_addr0_r_11), .AD2(rom_addr0_r_10), 
            .AD3(func_or_inet), .DO0(lx_ne0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam LUT4_0.initval = 16'b1111111111111110;
    INV INV_1 (.A(lx_ne0), .Z(lx_ne0_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    AND2 AND2_t0 (.A(mx_ctrl_r), .B(lx_ne0_inv), .Z(out_sel_i)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(305[10:64])
    FD1P3DX FF_62 (.D(\phase_accum[56] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(rom_addr0_r)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(309[13:86])
    defparam FF_62.GSR = "ENABLED";
    MUX21 muxb_56 (.D0(rom_addr0_r_1), .D1(rom_addr0_r_n_1), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_55 (.D0(rom_addr0_r_2), .D1(rom_addr0_r_n_2), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_54 (.D0(rom_addr0_r_3), .D1(rom_addr0_r_n_3), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_53 (.D0(rom_addr0_r_4), .D1(rom_addr0_r_n_4), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_52 (.D0(rom_addr0_r_5), .D1(rom_addr0_r_n_5), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    FD1P3DX FF_54 (.D(rom_dout_12_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(351[13] 352[25])
    defparam FF_54.GSR = "ENABLED";
    MUX21 muxb_50 (.D0(rom_dout_1), .D1(rom_dout_s_n_1), .SD(sinromoutsel), 
          .Z(rom_dout_s_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_49 (.D0(rom_dout_2), .D1(rom_dout_s_n_2), .SD(sinromoutsel), 
          .Z(rom_dout_s_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_48 (.D0(rom_dout_3), .D1(rom_dout_s_n_3), .SD(sinromoutsel), 
          .Z(rom_dout_s_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_47 (.D0(rom_dout_4), .D1(rom_dout_s_n_4), .SD(sinromoutsel), 
          .Z(rom_dout_s_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_46 (.D0(rom_dout_5), .D1(rom_dout_s_n_5), .SD(sinromoutsel), 
          .Z(rom_dout_s_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_45 (.D0(rom_dout_6), .D1(rom_dout_s_n_6), .SD(sinromoutsel), 
          .Z(rom_dout_s_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_44 (.D0(rom_dout_7), .D1(rom_dout_s_n_7), .SD(sinromoutsel), 
          .Z(rom_dout_s_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_43 (.D0(rom_dout_8), .D1(rom_dout_s_n_8), .SD(sinromoutsel), 
          .Z(rom_dout_s_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_42 (.D0(rom_dout_9), .D1(rom_dout_s_n_9), .SD(sinromoutsel), 
          .Z(rom_dout_s_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_41 (.D0(rom_dout_10), .D1(rom_dout_s_n_10), .SD(sinromoutsel), 
          .Z(rom_dout_s_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_40 (.D0(rom_dout_11), .D1(rom_dout_s_n_11), .SD(sinromoutsel), 
          .Z(rom_dout_s_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_39 (.D0(rom_dout_12), .D1(rom_dout_s_n_12), .SD(sinromoutsel), 
          .Z(rom_dout_s_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_37 (.D0(rom_dout_14), .D1(rom_dout_c_n_1), .SD(cosromoutsel), 
          .Z(rom_dout_c_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_36 (.D0(rom_dout_15), .D1(rom_dout_c_n_2), .SD(cosromoutsel), 
          .Z(rom_dout_c_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_35 (.D0(rom_dout_16), .D1(rom_dout_c_n_3), .SD(cosromoutsel), 
          .Z(rom_dout_c_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_34 (.D0(rom_dout_17), .D1(rom_dout_c_n_4), .SD(cosromoutsel), 
          .Z(rom_dout_c_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_33 (.D0(rom_dout_18), .D1(rom_dout_c_n_5), .SD(cosromoutsel), 
          .Z(rom_dout_c_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_32 (.D0(rom_dout_19), .D1(rom_dout_c_n_6), .SD(cosromoutsel), 
          .Z(rom_dout_c_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_31 (.D0(rom_dout_20), .D1(rom_dout_c_n_7), .SD(cosromoutsel), 
          .Z(rom_dout_c_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_30 (.D0(rom_dout_21), .D1(rom_dout_c_n_8), .SD(cosromoutsel), 
          .Z(rom_dout_c_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_29 (.D0(rom_dout_22), .D1(rom_dout_c_n_9), .SD(cosromoutsel), 
          .Z(rom_dout_c_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_28 (.D0(rom_dout_23), .D1(rom_dout_c_n_10), .SD(cosromoutsel), 
          .Z(rom_dout_c_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_27 (.D0(rom_dout_24), .D1(rom_dout_c_n_11), .SD(cosromoutsel), 
          .Z(rom_dout_c_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_26 (.D0(rom_dout_25), .D1(rom_dout_c_n_12), .SD(cosromoutsel), 
          .Z(rom_dout_c_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    FD1P3DX FF_26 (.D(out_sel_i), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(out_sel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(541[13:83])
    defparam FF_26.GSR = "ENABLED";
    MUX21 muxb_24 (.D0(rom_dout_s_1), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_23 (.D0(rom_dout_s_2), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_22 (.D0(rom_dout_s_3), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_21 (.D0(rom_dout_s_4), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_20 (.D0(rom_dout_s_5), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_19 (.D0(rom_dout_s_6), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_18 (.D0(rom_dout_s_7), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_17 (.D0(rom_dout_s_8), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_16 (.D0(rom_dout_s_9), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_15 (.D0(rom_dout_s_10), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_14 (.D0(rom_dout_s_11), .D1(VCC_net), .SD(out_sel), .Z(sinout_pre_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_13 (.D0(rom_dout_s_12), .D1(mx_ctrl_r_1), .SD(out_sel), 
          .Z(sinout_pre_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_11 (.D0(rom_dout_c_1), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_10 (.D0(rom_dout_c_2), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_9 (.D0(rom_dout_c_3), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_8 (.D0(rom_dout_c_4), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_7 (.D0(rom_dout_c_5), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_6 (.D0(rom_dout_c_6), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_5 (.D0(rom_dout_c_7), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_4 (.D0(rom_dout_c_8), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_3 (.D0(rom_dout_c_9), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_2 (.D0(rom_dout_c_10), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_1 (.D0(rom_dout_c_11), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    MUX21 muxb_0 (.D0(rom_dout_c_12), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    ROM64X1A triglut_1_0_24 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_11_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_24.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    ROM64X1A triglut_1_0_23 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_10_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_23.initval = 64'b1111111111111111111111111111111111111111110000000000000000000000;
    ROM64X1A triglut_1_0_22 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_9_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_22.initval = 64'b1111111111111111111111111111100000000000001111111111100000000000;
    ROM64X1A triglut_1_0_21 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_8_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_21.initval = 64'b1111111111111111111100000000011111110000001111110000011111000000;
    ROM64X1A triglut_1_0_20 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_7_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_20.initval = 64'b1111111111111100000011111000011110001110001110001110011100111000;
    ROM64X1A triglut_1_0_19 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_6_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_19.initval = 64'b1111111111000011100011100110011001001101101101001001011010110100;
    ROM64X1A triglut_1_0_18 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_5_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_18.initval = 64'b1111111000110011011010010101010100101001001001101100110001100110;
    ROM64X1A triglut_1_0_17 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_4_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_17.initval = 64'b1111100100101010110011000000000001110011011010110101010110101010;
    ROM64X1A triglut_1_0_16 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_3_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_16.initval = 64'b1110010110011100010101001111111101101010110011100000000011110000;
    ROM64X1A triglut_1_0_15 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_2_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_15.initval = 64'b1101000010100011001111010111110011001100010101100000000011001100;
    ROM64X1A triglut_1_0_14 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_1_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_14.initval = 64'b1111011011100010010110111011101001110011000000100111110010101010;
    ROM64X1A triglut_1_0_13 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_13.initval = 64'b1000100101001010011001010111111001010010011110001001001001111000;
    ROM64X1A triglut_1_0_12 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_25_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_12.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    ROM64X1A triglut_1_0_11 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_24_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_11.initval = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    ROM64X1A triglut_1_0_10 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_23_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_10.initval = 64'b0000000000000000000001111111111111111111111111111111111111111110;
    ROM64X1A triglut_1_0_9 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_22_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_9.initval = 64'b0000000000111111111110000000000000111111111111111111111111111110;
    ROM64X1A triglut_1_0_8 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_21_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_8.initval = 64'b0000011111000001111110000001111111000000000111111111111111111110;
    ROM64X1A triglut_1_0_7 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_20_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_7.initval = 64'b0011100111001110001110001110001111000011111000000111111111111110;
    ROM64X1A triglut_1_0_6 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_19_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_6.initval = 64'b0101101011010010010110110110010011001100111000111000011111111110;
    ROM64X1A triglut_1_0_5 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_18_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_5.initval = 64'b1100110001100110110010010010100101010101001011011001100011111110;
    ROM64X1A triglut_1_0_4 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_17_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_4.initval = 64'b1010101101010101101011011001110000000000011001101010100100111110;
    ROM64X1A triglut_1_0_3 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_16_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_3.initval = 64'b0001111000000000111001101010110111111110010101000111001101001110;
    ROM64X1A triglut_1_0_2 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_15_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_2.initval = 64'b0110011000000000110101000110011001111101011110011000101000010110;
    ROM64X1A triglut_1_0_1 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_14_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_1.initval = 64'b1010101001111100100000011001110010111011101101001000111011011110;
    ROM64X1A triglut_1_0_0 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_13_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    defparam triglut_1_0_0.initval = 64'b0011110010010010001111001001010011111101010011001010010100100010;
    FADD2B neg_rom_dout_s_n_0 (.A0(GND_net), .A1(rom_dout_inv), .B0(GND_net), 
           .B1(VCC_net), .CI(GND_net), .COUT(co0_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=138, LSE_RLINE=145 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(138[8] 145[2])
    
endmodule
//
// Verilog Description of module Mixer
//

module Mixer (\LOCosine[12] , MixerOutSin, osc_clk, DiffOut_c, MixerOutCos, 
            RFIn_c, GND_net, \LOCosine[10] , \LOCosine[11] , \LOCosine[8] , 
            \LOCosine[9] , \LOCosine[6] , \LOCosine[7] , \LOCosine[4] , 
            \LOCosine[5] , \LOCosine[2] , \LOCosine[3] , \LOCosine[1] , 
            \LOSine[12] , \LOSine[10] , \LOSine[11] , \LOSine[8] , \LOSine[9] , 
            \LOSine[6] , \LOSine[7] , \LOSine[4] , \LOSine[5] , \LOSine[2] , 
            \LOSine[3] , \LOSine[1] ) /* synthesis syn_module_defined=1 */ ;
    input \LOCosine[12] ;
    output [11:0]MixerOutSin;
    input osc_clk;
    output DiffOut_c;
    output [11:0]MixerOutCos;
    input RFIn_c;
    input GND_net;
    input \LOCosine[10] ;
    input \LOCosine[11] ;
    input \LOCosine[8] ;
    input \LOCosine[9] ;
    input \LOCosine[6] ;
    input \LOCosine[7] ;
    input \LOCosine[4] ;
    input \LOCosine[5] ;
    input \LOCosine[2] ;
    input \LOCosine[3] ;
    input \LOCosine[1] ;
    input \LOSine[12] ;
    input \LOSine[10] ;
    input \LOSine[11] ;
    input \LOSine[8] ;
    input \LOSine[9] ;
    input \LOSine[6] ;
    input \LOSine[7] ;
    input \LOSine[4] ;
    input \LOSine[5] ;
    input \LOSine[2] ;
    input \LOSine[3] ;
    input \LOSine[1] ;
    
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(71[8:15])
    wire [11:0]MixerOutCos_11__N_250;
    
    wire RFInR;
    wire [11:0]MixerOutCos_11__N_224;
    wire [11:0]MixerOutSin_11__N_212;
    
    wire n11347, n11346, n11345, n11344, n11343, n11342, n11309;
    wire [11:0]MixerOutSin_11__N_236;
    
    wire n11308, n11307, n11306, n11305, n11304;
    
    LUT4 MixerOutCos_11__I_0_i12_3_lut (.A(\LOCosine[12] ), .B(MixerOutCos_11__N_250[11]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i12_3_lut.init = 16'hcaca;
    FD1S3AX MixerOutSin_i0 (.D(MixerOutSin_11__N_212[0]), .CK(osc_clk), 
            .Q(MixerOutSin[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i0.GSR = "ENABLED";
    FD1S3AY RFInR_14 (.D(DiffOut_c), .CK(osc_clk), .Q(RFInR)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(23[10] 27[8])
    defparam RFInR_14.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i0 (.D(MixerOutCos_11__N_224[0]), .CK(osc_clk), 
            .Q(MixerOutCos[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i0.GSR = "ENABLED";
    FD1S3AY RFInR1_13 (.D(RFIn_c), .CK(osc_clk), .Q(DiffOut_c)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(23[10] 27[8])
    defparam RFInR1_13.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i1 (.D(MixerOutSin_11__N_212[1]), .CK(osc_clk), 
            .Q(MixerOutSin[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i1.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i2 (.D(MixerOutSin_11__N_212[2]), .CK(osc_clk), 
            .Q(MixerOutSin[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i2.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i3 (.D(MixerOutSin_11__N_212[3]), .CK(osc_clk), 
            .Q(MixerOutSin[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i3.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i4 (.D(MixerOutSin_11__N_212[4]), .CK(osc_clk), 
            .Q(MixerOutSin[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i4.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i5 (.D(MixerOutSin_11__N_212[5]), .CK(osc_clk), 
            .Q(MixerOutSin[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i5.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i6 (.D(MixerOutSin_11__N_212[6]), .CK(osc_clk), 
            .Q(MixerOutSin[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i6.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i7 (.D(MixerOutSin_11__N_212[7]), .CK(osc_clk), 
            .Q(MixerOutSin[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i7.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i8 (.D(MixerOutSin_11__N_212[8]), .CK(osc_clk), 
            .Q(MixerOutSin[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i8.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i9 (.D(MixerOutSin_11__N_212[9]), .CK(osc_clk), 
            .Q(MixerOutSin[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i9.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i10 (.D(MixerOutSin_11__N_212[10]), .CK(osc_clk), 
            .Q(MixerOutSin[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i10.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i11 (.D(MixerOutSin_11__N_212[11]), .CK(osc_clk), 
            .Q(MixerOutSin[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i11.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i1 (.D(MixerOutCos_11__N_224[1]), .CK(osc_clk), 
            .Q(MixerOutCos[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i1.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i2 (.D(MixerOutCos_11__N_224[2]), .CK(osc_clk), 
            .Q(MixerOutCos[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i2.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i3 (.D(MixerOutCos_11__N_224[3]), .CK(osc_clk), 
            .Q(MixerOutCos[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i3.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i4 (.D(MixerOutCos_11__N_224[4]), .CK(osc_clk), 
            .Q(MixerOutCos[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i4.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i5 (.D(MixerOutCos_11__N_224[5]), .CK(osc_clk), 
            .Q(MixerOutCos[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i5.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i6 (.D(MixerOutCos_11__N_224[6]), .CK(osc_clk), 
            .Q(MixerOutCos[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i6.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i7 (.D(MixerOutCos_11__N_224[7]), .CK(osc_clk), 
            .Q(MixerOutCos[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i7.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i8 (.D(MixerOutCos_11__N_224[8]), .CK(osc_clk), 
            .Q(MixerOutCos[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i8.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i9 (.D(MixerOutCos_11__N_224[9]), .CK(osc_clk), 
            .Q(MixerOutCos[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i9.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i10 (.D(MixerOutCos_11__N_224[10]), .CK(osc_clk), 
            .Q(MixerOutCos[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i10.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i11 (.D(MixerOutCos_11__N_224[11]), .CK(osc_clk), 
            .Q(MixerOutCos[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=157, LSE_RLINE=165 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i11.GSR = "ENABLED";
    CCU2D unary_minus_7_add_3_13 (.A0(\LOCosine[12] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11347), .S0(MixerOutCos_11__N_250[11]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(42[26:33])
    defparam unary_minus_7_add_3_13.INIT0 = 16'hf555;
    defparam unary_minus_7_add_3_13.INIT1 = 16'h0000;
    defparam unary_minus_7_add_3_13.INJECT1_0 = "NO";
    defparam unary_minus_7_add_3_13.INJECT1_1 = "NO";
    CCU2D unary_minus_7_add_3_11 (.A0(\LOCosine[10] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOCosine[11] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11346), .COUT(n11347), .S0(MixerOutCos_11__N_250[9]), 
          .S1(MixerOutCos_11__N_250[10]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(42[26:33])
    defparam unary_minus_7_add_3_11.INIT0 = 16'hf555;
    defparam unary_minus_7_add_3_11.INIT1 = 16'hf555;
    defparam unary_minus_7_add_3_11.INJECT1_0 = "NO";
    defparam unary_minus_7_add_3_11.INJECT1_1 = "NO";
    CCU2D unary_minus_7_add_3_9 (.A0(\LOCosine[8] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOCosine[9] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11345), .COUT(n11346), .S0(MixerOutCos_11__N_250[7]), 
          .S1(MixerOutCos_11__N_250[8]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(42[26:33])
    defparam unary_minus_7_add_3_9.INIT0 = 16'hf555;
    defparam unary_minus_7_add_3_9.INIT1 = 16'hf555;
    defparam unary_minus_7_add_3_9.INJECT1_0 = "NO";
    defparam unary_minus_7_add_3_9.INJECT1_1 = "NO";
    CCU2D unary_minus_7_add_3_7 (.A0(\LOCosine[6] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOCosine[7] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11344), .COUT(n11345), .S0(MixerOutCos_11__N_250[5]), 
          .S1(MixerOutCos_11__N_250[6]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(42[26:33])
    defparam unary_minus_7_add_3_7.INIT0 = 16'hf555;
    defparam unary_minus_7_add_3_7.INIT1 = 16'hf555;
    defparam unary_minus_7_add_3_7.INJECT1_0 = "NO";
    defparam unary_minus_7_add_3_7.INJECT1_1 = "NO";
    CCU2D unary_minus_7_add_3_5 (.A0(\LOCosine[4] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOCosine[5] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11343), .COUT(n11344), .S0(MixerOutCos_11__N_250[3]), 
          .S1(MixerOutCos_11__N_250[4]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(42[26:33])
    defparam unary_minus_7_add_3_5.INIT0 = 16'hf555;
    defparam unary_minus_7_add_3_5.INIT1 = 16'hf555;
    defparam unary_minus_7_add_3_5.INJECT1_0 = "NO";
    defparam unary_minus_7_add_3_5.INJECT1_1 = "NO";
    CCU2D unary_minus_7_add_3_3 (.A0(\LOCosine[2] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOCosine[3] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11342), .COUT(n11343), .S0(MixerOutCos_11__N_250[1]), 
          .S1(MixerOutCos_11__N_250[2]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(42[26:33])
    defparam unary_minus_7_add_3_3.INIT0 = 16'hf555;
    defparam unary_minus_7_add_3_3.INIT1 = 16'hf555;
    defparam unary_minus_7_add_3_3.INJECT1_0 = "NO";
    defparam unary_minus_7_add_3_3.INJECT1_1 = "NO";
    CCU2D unary_minus_7_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOCosine[1] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n11342), .S1(MixerOutCos_11__N_250[0]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(42[26:33])
    defparam unary_minus_7_add_3_1.INIT0 = 16'hF000;
    defparam unary_minus_7_add_3_1.INIT1 = 16'h0aaa;
    defparam unary_minus_7_add_3_1.INJECT1_0 = "NO";
    defparam unary_minus_7_add_3_1.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_13 (.A0(\LOSine[12] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11309), .S0(MixerOutSin_11__N_236[11]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(41[26:33])
    defparam unary_minus_6_add_3_13.INIT0 = 16'hf555;
    defparam unary_minus_6_add_3_13.INIT1 = 16'h0000;
    defparam unary_minus_6_add_3_13.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_13.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_11 (.A0(\LOSine[10] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOSine[11] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11308), .COUT(n11309), .S0(MixerOutSin_11__N_236[9]), 
          .S1(MixerOutSin_11__N_236[10]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(41[26:33])
    defparam unary_minus_6_add_3_11.INIT0 = 16'hf555;
    defparam unary_minus_6_add_3_11.INIT1 = 16'hf555;
    defparam unary_minus_6_add_3_11.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_11.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_9 (.A0(\LOSine[8] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOSine[9] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11307), .COUT(n11308), .S0(MixerOutSin_11__N_236[7]), 
          .S1(MixerOutSin_11__N_236[8]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(41[26:33])
    defparam unary_minus_6_add_3_9.INIT0 = 16'hf555;
    defparam unary_minus_6_add_3_9.INIT1 = 16'hf555;
    defparam unary_minus_6_add_3_9.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_9.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_7 (.A0(\LOSine[6] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOSine[7] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11306), .COUT(n11307), .S0(MixerOutSin_11__N_236[5]), 
          .S1(MixerOutSin_11__N_236[6]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(41[26:33])
    defparam unary_minus_6_add_3_7.INIT0 = 16'hf555;
    defparam unary_minus_6_add_3_7.INIT1 = 16'hf555;
    defparam unary_minus_6_add_3_7.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_7.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_5 (.A0(\LOSine[4] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOSine[5] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11305), .COUT(n11306), .S0(MixerOutSin_11__N_236[3]), 
          .S1(MixerOutSin_11__N_236[4]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(41[26:33])
    defparam unary_minus_6_add_3_5.INIT0 = 16'hf555;
    defparam unary_minus_6_add_3_5.INIT1 = 16'hf555;
    defparam unary_minus_6_add_3_5.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_5.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_3 (.A0(\LOSine[2] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOSine[3] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11304), .COUT(n11305), .S0(MixerOutSin_11__N_236[1]), 
          .S1(MixerOutSin_11__N_236[2]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(41[26:33])
    defparam unary_minus_6_add_3_3.INIT0 = 16'hf555;
    defparam unary_minus_6_add_3_3.INIT1 = 16'hf555;
    defparam unary_minus_6_add_3_3.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_3.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOSine[1] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n11304), .S1(MixerOutSin_11__N_236[0]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(41[26:33])
    defparam unary_minus_6_add_3_1.INIT0 = 16'hF000;
    defparam unary_minus_6_add_3_1.INIT1 = 16'h0aaa;
    defparam unary_minus_6_add_3_1.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_1.INJECT1_1 = "NO";
    LUT4 MixerOutSin_11__I_0_i1_3_lut (.A(\LOSine[1] ), .B(MixerOutSin_11__N_236[0]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i1_3_lut (.A(\LOCosine[1] ), .B(MixerOutCos_11__N_250[0]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i2_3_lut (.A(\LOSine[2] ), .B(MixerOutSin_11__N_236[1]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i3_3_lut (.A(\LOSine[3] ), .B(MixerOutSin_11__N_236[2]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i4_3_lut (.A(\LOSine[4] ), .B(MixerOutSin_11__N_236[3]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i5_3_lut (.A(\LOSine[5] ), .B(MixerOutSin_11__N_236[4]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i6_3_lut (.A(\LOSine[6] ), .B(MixerOutSin_11__N_236[5]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i7_3_lut (.A(\LOSine[7] ), .B(MixerOutSin_11__N_236[6]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i8_3_lut (.A(\LOSine[8] ), .B(MixerOutSin_11__N_236[7]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i9_3_lut (.A(\LOSine[9] ), .B(MixerOutSin_11__N_236[8]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i10_3_lut (.A(\LOSine[10] ), .B(MixerOutSin_11__N_236[9]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i11_3_lut (.A(\LOSine[11] ), .B(MixerOutSin_11__N_236[10]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i12_3_lut (.A(\LOSine[12] ), .B(MixerOutSin_11__N_236[11]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i2_3_lut (.A(\LOCosine[2] ), .B(MixerOutCos_11__N_250[1]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i3_3_lut (.A(\LOCosine[3] ), .B(MixerOutCos_11__N_250[2]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i4_3_lut (.A(\LOCosine[4] ), .B(MixerOutCos_11__N_250[3]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i5_3_lut (.A(\LOCosine[5] ), .B(MixerOutCos_11__N_250[4]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i6_3_lut (.A(\LOCosine[6] ), .B(MixerOutCos_11__N_250[5]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i7_3_lut (.A(\LOCosine[7] ), .B(MixerOutCos_11__N_250[6]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i8_3_lut (.A(\LOCosine[8] ), .B(MixerOutCos_11__N_250[7]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i9_3_lut (.A(\LOCosine[9] ), .B(MixerOutCos_11__N_250[8]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i10_3_lut (.A(\LOCosine[10] ), .B(MixerOutCos_11__N_250[9]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i11_3_lut (.A(\LOCosine[11] ), .B(MixerOutCos_11__N_250[10]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i11_3_lut.init = 16'hcaca;
    
endmodule
//
// Verilog Description of module nco_sig
//

module nco_sig (osc_clk, \phase_accum[56] , \phase_accum[57] , \phase_accum[58] , 
            \phase_accum[59] , \phase_accum[60] , \phase_accum[61] , \phase_accum[62] , 
            \phase_accum[63] , phase_inc_carrGen1, GND_net, sinGen_c) /* synthesis syn_module_defined=1 */ ;
    input osc_clk;
    output \phase_accum[56] ;
    output \phase_accum[57] ;
    output \phase_accum[58] ;
    output \phase_accum[59] ;
    output \phase_accum[60] ;
    output \phase_accum[61] ;
    output \phase_accum[62] ;
    output \phase_accum[63] ;
    input [63:0]phase_inc_carrGen1;
    input GND_net;
    output sinGen_c;
    
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(71[8:15])
    wire [63:0]phase_accum;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(29[19:30])
    wire [63:0]phase_accum_63__N_146;
    
    wire n10985, n10984, n10983, n10982, n10981, n10980, n10979, 
        n10978, n10977, n10976, n10975, n10974, n10973, n10972, 
        n10971, n10970, n10969, n10968, n10967, n10966, n10965, 
        n10964, n10963, n10962, n10961, n10960, n10959, n10958, 
        n10957, n10956, n10955;
    
    FD1S3AX phase_accum_i0 (.D(phase_accum_63__N_146[0]), .CK(osc_clk), 
            .Q(phase_accum[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i0.GSR = "ENABLED";
    FD1S3AX phase_accum_i1 (.D(phase_accum_63__N_146[1]), .CK(osc_clk), 
            .Q(phase_accum[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i1.GSR = "ENABLED";
    FD1S3AX phase_accum_i2 (.D(phase_accum_63__N_146[2]), .CK(osc_clk), 
            .Q(phase_accum[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i2.GSR = "ENABLED";
    FD1S3AX phase_accum_i3 (.D(phase_accum_63__N_146[3]), .CK(osc_clk), 
            .Q(phase_accum[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i3.GSR = "ENABLED";
    FD1S3AX phase_accum_i4 (.D(phase_accum_63__N_146[4]), .CK(osc_clk), 
            .Q(phase_accum[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i4.GSR = "ENABLED";
    FD1S3AX phase_accum_i5 (.D(phase_accum_63__N_146[5]), .CK(osc_clk), 
            .Q(phase_accum[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i5.GSR = "ENABLED";
    FD1S3AX phase_accum_i6 (.D(phase_accum_63__N_146[6]), .CK(osc_clk), 
            .Q(phase_accum[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i6.GSR = "ENABLED";
    FD1S3AX phase_accum_i7 (.D(phase_accum_63__N_146[7]), .CK(osc_clk), 
            .Q(phase_accum[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i7.GSR = "ENABLED";
    FD1S3AX phase_accum_i8 (.D(phase_accum_63__N_146[8]), .CK(osc_clk), 
            .Q(phase_accum[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i8.GSR = "ENABLED";
    FD1S3AX phase_accum_i9 (.D(phase_accum_63__N_146[9]), .CK(osc_clk), 
            .Q(phase_accum[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i9.GSR = "ENABLED";
    FD1S3AX phase_accum_i10 (.D(phase_accum_63__N_146[10]), .CK(osc_clk), 
            .Q(phase_accum[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i10.GSR = "ENABLED";
    FD1S3AX phase_accum_i11 (.D(phase_accum_63__N_146[11]), .CK(osc_clk), 
            .Q(phase_accum[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i11.GSR = "ENABLED";
    FD1S3AX phase_accum_i12 (.D(phase_accum_63__N_146[12]), .CK(osc_clk), 
            .Q(phase_accum[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i12.GSR = "ENABLED";
    FD1S3AX phase_accum_i13 (.D(phase_accum_63__N_146[13]), .CK(osc_clk), 
            .Q(phase_accum[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i13.GSR = "ENABLED";
    FD1S3AX phase_accum_i14 (.D(phase_accum_63__N_146[14]), .CK(osc_clk), 
            .Q(phase_accum[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i14.GSR = "ENABLED";
    FD1S3AX phase_accum_i15 (.D(phase_accum_63__N_146[15]), .CK(osc_clk), 
            .Q(phase_accum[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i15.GSR = "ENABLED";
    FD1S3AX phase_accum_i16 (.D(phase_accum_63__N_146[16]), .CK(osc_clk), 
            .Q(phase_accum[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i16.GSR = "ENABLED";
    FD1S3AX phase_accum_i17 (.D(phase_accum_63__N_146[17]), .CK(osc_clk), 
            .Q(phase_accum[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i17.GSR = "ENABLED";
    FD1S3AX phase_accum_i18 (.D(phase_accum_63__N_146[18]), .CK(osc_clk), 
            .Q(phase_accum[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i18.GSR = "ENABLED";
    FD1S3AX phase_accum_i19 (.D(phase_accum_63__N_146[19]), .CK(osc_clk), 
            .Q(phase_accum[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i19.GSR = "ENABLED";
    FD1S3AX phase_accum_i20 (.D(phase_accum_63__N_146[20]), .CK(osc_clk), 
            .Q(phase_accum[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i20.GSR = "ENABLED";
    FD1S3AX phase_accum_i21 (.D(phase_accum_63__N_146[21]), .CK(osc_clk), 
            .Q(phase_accum[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i21.GSR = "ENABLED";
    FD1S3AX phase_accum_i22 (.D(phase_accum_63__N_146[22]), .CK(osc_clk), 
            .Q(phase_accum[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i22.GSR = "ENABLED";
    FD1S3AX phase_accum_i23 (.D(phase_accum_63__N_146[23]), .CK(osc_clk), 
            .Q(phase_accum[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i23.GSR = "ENABLED";
    FD1S3AX phase_accum_i24 (.D(phase_accum_63__N_146[24]), .CK(osc_clk), 
            .Q(phase_accum[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i24.GSR = "ENABLED";
    FD1S3AX phase_accum_i25 (.D(phase_accum_63__N_146[25]), .CK(osc_clk), 
            .Q(phase_accum[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i25.GSR = "ENABLED";
    FD1S3AX phase_accum_i26 (.D(phase_accum_63__N_146[26]), .CK(osc_clk), 
            .Q(phase_accum[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i26.GSR = "ENABLED";
    FD1S3AX phase_accum_i27 (.D(phase_accum_63__N_146[27]), .CK(osc_clk), 
            .Q(phase_accum[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i27.GSR = "ENABLED";
    FD1S3AX phase_accum_i28 (.D(phase_accum_63__N_146[28]), .CK(osc_clk), 
            .Q(phase_accum[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i28.GSR = "ENABLED";
    FD1S3AX phase_accum_i29 (.D(phase_accum_63__N_146[29]), .CK(osc_clk), 
            .Q(phase_accum[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i29.GSR = "ENABLED";
    FD1S3AX phase_accum_i30 (.D(phase_accum_63__N_146[30]), .CK(osc_clk), 
            .Q(phase_accum[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i30.GSR = "ENABLED";
    FD1S3AX phase_accum_i31 (.D(phase_accum_63__N_146[31]), .CK(osc_clk), 
            .Q(phase_accum[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i31.GSR = "ENABLED";
    FD1S3AX phase_accum_i32 (.D(phase_accum_63__N_146[32]), .CK(osc_clk), 
            .Q(phase_accum[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i32.GSR = "ENABLED";
    FD1S3AX phase_accum_i33 (.D(phase_accum_63__N_146[33]), .CK(osc_clk), 
            .Q(phase_accum[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i33.GSR = "ENABLED";
    FD1S3AX phase_accum_i34 (.D(phase_accum_63__N_146[34]), .CK(osc_clk), 
            .Q(phase_accum[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i34.GSR = "ENABLED";
    FD1S3AX phase_accum_i35 (.D(phase_accum_63__N_146[35]), .CK(osc_clk), 
            .Q(phase_accum[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i35.GSR = "ENABLED";
    FD1S3AX phase_accum_i36 (.D(phase_accum_63__N_146[36]), .CK(osc_clk), 
            .Q(phase_accum[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i36.GSR = "ENABLED";
    FD1S3AX phase_accum_i37 (.D(phase_accum_63__N_146[37]), .CK(osc_clk), 
            .Q(phase_accum[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i37.GSR = "ENABLED";
    FD1S3AX phase_accum_i38 (.D(phase_accum_63__N_146[38]), .CK(osc_clk), 
            .Q(phase_accum[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i38.GSR = "ENABLED";
    FD1S3AX phase_accum_i39 (.D(phase_accum_63__N_146[39]), .CK(osc_clk), 
            .Q(phase_accum[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i39.GSR = "ENABLED";
    FD1S3AX phase_accum_i40 (.D(phase_accum_63__N_146[40]), .CK(osc_clk), 
            .Q(phase_accum[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i40.GSR = "ENABLED";
    FD1S3AX phase_accum_i41 (.D(phase_accum_63__N_146[41]), .CK(osc_clk), 
            .Q(phase_accum[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i41.GSR = "ENABLED";
    FD1S3AX phase_accum_i42 (.D(phase_accum_63__N_146[42]), .CK(osc_clk), 
            .Q(phase_accum[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i42.GSR = "ENABLED";
    FD1S3AX phase_accum_i43 (.D(phase_accum_63__N_146[43]), .CK(osc_clk), 
            .Q(phase_accum[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i43.GSR = "ENABLED";
    FD1S3AX phase_accum_i44 (.D(phase_accum_63__N_146[44]), .CK(osc_clk), 
            .Q(phase_accum[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i44.GSR = "ENABLED";
    FD1S3AX phase_accum_i45 (.D(phase_accum_63__N_146[45]), .CK(osc_clk), 
            .Q(phase_accum[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i45.GSR = "ENABLED";
    FD1S3AX phase_accum_i46 (.D(phase_accum_63__N_146[46]), .CK(osc_clk), 
            .Q(phase_accum[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i46.GSR = "ENABLED";
    FD1S3AX phase_accum_i47 (.D(phase_accum_63__N_146[47]), .CK(osc_clk), 
            .Q(phase_accum[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i47.GSR = "ENABLED";
    FD1S3AX phase_accum_i48 (.D(phase_accum_63__N_146[48]), .CK(osc_clk), 
            .Q(phase_accum[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i48.GSR = "ENABLED";
    FD1S3AX phase_accum_i49 (.D(phase_accum_63__N_146[49]), .CK(osc_clk), 
            .Q(phase_accum[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i49.GSR = "ENABLED";
    FD1S3AX phase_accum_i50 (.D(phase_accum_63__N_146[50]), .CK(osc_clk), 
            .Q(phase_accum[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i50.GSR = "ENABLED";
    FD1S3AX phase_accum_i51 (.D(phase_accum_63__N_146[51]), .CK(osc_clk), 
            .Q(phase_accum[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i51.GSR = "ENABLED";
    FD1S3AX phase_accum_i52 (.D(phase_accum_63__N_146[52]), .CK(osc_clk), 
            .Q(phase_accum[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i52.GSR = "ENABLED";
    FD1S3AX phase_accum_i53 (.D(phase_accum_63__N_146[53]), .CK(osc_clk), 
            .Q(phase_accum[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i53.GSR = "ENABLED";
    FD1S3AX phase_accum_i54 (.D(phase_accum_63__N_146[54]), .CK(osc_clk), 
            .Q(phase_accum[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i54.GSR = "ENABLED";
    FD1S3AX phase_accum_i55 (.D(phase_accum_63__N_146[55]), .CK(osc_clk), 
            .Q(phase_accum[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i55.GSR = "ENABLED";
    FD1S3AX phase_accum_i56 (.D(phase_accum_63__N_146[56]), .CK(osc_clk), 
            .Q(\phase_accum[56] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i56.GSR = "ENABLED";
    FD1S3AX phase_accum_i57 (.D(phase_accum_63__N_146[57]), .CK(osc_clk), 
            .Q(\phase_accum[57] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i57.GSR = "ENABLED";
    FD1S3AX phase_accum_i58 (.D(phase_accum_63__N_146[58]), .CK(osc_clk), 
            .Q(\phase_accum[58] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i58.GSR = "ENABLED";
    FD1S3AX phase_accum_i59 (.D(phase_accum_63__N_146[59]), .CK(osc_clk), 
            .Q(\phase_accum[59] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i59.GSR = "ENABLED";
    FD1S3AX phase_accum_i60 (.D(phase_accum_63__N_146[60]), .CK(osc_clk), 
            .Q(\phase_accum[60] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i60.GSR = "ENABLED";
    FD1S3AX phase_accum_i61 (.D(phase_accum_63__N_146[61]), .CK(osc_clk), 
            .Q(\phase_accum[61] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i61.GSR = "ENABLED";
    FD1S3AX phase_accum_i62 (.D(phase_accum_63__N_146[62]), .CK(osc_clk), 
            .Q(\phase_accum[62] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i62.GSR = "ENABLED";
    FD1S3AX phase_accum_i63 (.D(phase_accum_63__N_146[63]), .CK(osc_clk), 
            .Q(\phase_accum[63] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=148, LSE_RLINE=154 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i63.GSR = "ENABLED";
    CCU2D phase_accum_63__I_0_12_64 (.A0(\phase_accum[62] ), .B0(phase_inc_carrGen1[62]), 
          .C0(GND_net), .D0(GND_net), .A1(\phase_accum[63] ), .B1(phase_inc_carrGen1[63]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10985), .S0(phase_accum_63__N_146[62]), 
          .S1(phase_accum_63__N_146[63]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_64.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_64.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_64.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_64.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_62 (.A0(\phase_accum[60] ), .B0(phase_inc_carrGen1[60]), 
          .C0(GND_net), .D0(GND_net), .A1(\phase_accum[61] ), .B1(phase_inc_carrGen1[61]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10984), .COUT(n10985), .S0(phase_accum_63__N_146[60]), 
          .S1(phase_accum_63__N_146[61]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_62.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_62.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_62.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_62.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_60 (.A0(\phase_accum[58] ), .B0(phase_inc_carrGen1[58]), 
          .C0(GND_net), .D0(GND_net), .A1(\phase_accum[59] ), .B1(phase_inc_carrGen1[59]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10983), .COUT(n10984), .S0(phase_accum_63__N_146[58]), 
          .S1(phase_accum_63__N_146[59]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_60.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_60.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_60.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_60.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_58 (.A0(\phase_accum[56] ), .B0(phase_inc_carrGen1[56]), 
          .C0(GND_net), .D0(GND_net), .A1(\phase_accum[57] ), .B1(phase_inc_carrGen1[57]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10982), .COUT(n10983), .S0(phase_accum_63__N_146[56]), 
          .S1(phase_accum_63__N_146[57]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_58.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_58.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_58.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_58.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_56 (.A0(phase_accum[54]), .B0(phase_inc_carrGen1[54]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[55]), .B1(phase_inc_carrGen1[55]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10981), .COUT(n10982), .S0(phase_accum_63__N_146[54]), 
          .S1(phase_accum_63__N_146[55]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_56.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_56.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_56.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_56.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_54 (.A0(phase_accum[52]), .B0(phase_inc_carrGen1[52]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[53]), .B1(phase_inc_carrGen1[53]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10980), .COUT(n10981), .S0(phase_accum_63__N_146[52]), 
          .S1(phase_accum_63__N_146[53]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_54.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_54.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_54.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_54.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_52 (.A0(phase_accum[50]), .B0(phase_inc_carrGen1[50]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[51]), .B1(phase_inc_carrGen1[51]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10979), .COUT(n10980), .S0(phase_accum_63__N_146[50]), 
          .S1(phase_accum_63__N_146[51]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_52.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_52.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_52.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_52.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_50 (.A0(phase_accum[48]), .B0(phase_inc_carrGen1[48]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[49]), .B1(phase_inc_carrGen1[49]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10978), .COUT(n10979), .S0(phase_accum_63__N_146[48]), 
          .S1(phase_accum_63__N_146[49]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_50.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_50.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_50.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_50.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_48 (.A0(phase_accum[46]), .B0(phase_inc_carrGen1[46]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[47]), .B1(phase_inc_carrGen1[47]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10977), .COUT(n10978), .S0(phase_accum_63__N_146[46]), 
          .S1(phase_accum_63__N_146[47]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_48.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_48.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_48.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_48.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_46 (.A0(phase_accum[44]), .B0(phase_inc_carrGen1[44]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[45]), .B1(phase_inc_carrGen1[45]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10976), .COUT(n10977), .S0(phase_accum_63__N_146[44]), 
          .S1(phase_accum_63__N_146[45]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_46.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_46.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_46.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_46.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_44 (.A0(phase_accum[42]), .B0(phase_inc_carrGen1[42]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[43]), .B1(phase_inc_carrGen1[43]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10975), .COUT(n10976), .S0(phase_accum_63__N_146[42]), 
          .S1(phase_accum_63__N_146[43]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_44.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_44.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_44.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_44.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_42 (.A0(phase_accum[40]), .B0(phase_inc_carrGen1[40]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[41]), .B1(phase_inc_carrGen1[41]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10974), .COUT(n10975), .S0(phase_accum_63__N_146[40]), 
          .S1(phase_accum_63__N_146[41]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_42.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_42.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_42.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_42.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_40 (.A0(phase_accum[38]), .B0(phase_inc_carrGen1[38]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[39]), .B1(phase_inc_carrGen1[39]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10973), .COUT(n10974), .S0(phase_accum_63__N_146[38]), 
          .S1(phase_accum_63__N_146[39]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_40.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_40.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_40.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_40.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_38 (.A0(phase_accum[36]), .B0(phase_inc_carrGen1[36]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[37]), .B1(phase_inc_carrGen1[37]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10972), .COUT(n10973), .S0(phase_accum_63__N_146[36]), 
          .S1(phase_accum_63__N_146[37]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_38.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_38.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_38.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_38.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_36 (.A0(phase_accum[34]), .B0(phase_inc_carrGen1[34]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[35]), .B1(phase_inc_carrGen1[35]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10971), .COUT(n10972), .S0(phase_accum_63__N_146[34]), 
          .S1(phase_accum_63__N_146[35]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_36.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_36.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_36.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_36.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_34 (.A0(phase_accum[32]), .B0(phase_inc_carrGen1[32]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[33]), .B1(phase_inc_carrGen1[33]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10970), .COUT(n10971), .S0(phase_accum_63__N_146[32]), 
          .S1(phase_accum_63__N_146[33]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_34.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_34.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_34.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_34.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_32 (.A0(phase_accum[30]), .B0(phase_inc_carrGen1[30]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[31]), .B1(phase_inc_carrGen1[31]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10969), .COUT(n10970), .S0(phase_accum_63__N_146[30]), 
          .S1(phase_accum_63__N_146[31]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_32.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_32.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_32.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_32.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_30 (.A0(phase_accum[28]), .B0(phase_inc_carrGen1[28]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[29]), .B1(phase_inc_carrGen1[29]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10968), .COUT(n10969), .S0(phase_accum_63__N_146[28]), 
          .S1(phase_accum_63__N_146[29]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_30.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_30.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_30.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_30.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_28 (.A0(phase_accum[26]), .B0(phase_inc_carrGen1[26]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[27]), .B1(phase_inc_carrGen1[27]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10967), .COUT(n10968), .S0(phase_accum_63__N_146[26]), 
          .S1(phase_accum_63__N_146[27]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_28.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_28.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_28.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_28.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_26 (.A0(phase_accum[24]), .B0(phase_inc_carrGen1[24]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[25]), .B1(phase_inc_carrGen1[25]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10966), .COUT(n10967), .S0(phase_accum_63__N_146[24]), 
          .S1(phase_accum_63__N_146[25]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_26.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_26.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_26.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_26.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_24 (.A0(phase_accum[22]), .B0(phase_inc_carrGen1[22]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[23]), .B1(phase_inc_carrGen1[23]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10965), .COUT(n10966), .S0(phase_accum_63__N_146[22]), 
          .S1(phase_accum_63__N_146[23]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_24.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_24.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_24.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_24.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_22 (.A0(phase_accum[20]), .B0(phase_inc_carrGen1[20]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[21]), .B1(phase_inc_carrGen1[21]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10964), .COUT(n10965), .S0(phase_accum_63__N_146[20]), 
          .S1(phase_accum_63__N_146[21]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_22.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_22.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_22.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_22.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_20 (.A0(phase_accum[18]), .B0(phase_inc_carrGen1[18]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[19]), .B1(phase_inc_carrGen1[19]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10963), .COUT(n10964), .S0(phase_accum_63__N_146[18]), 
          .S1(phase_accum_63__N_146[19]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_20.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_20.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_20.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_20.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_18 (.A0(phase_accum[16]), .B0(phase_inc_carrGen1[16]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[17]), .B1(phase_inc_carrGen1[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10962), .COUT(n10963), .S0(phase_accum_63__N_146[16]), 
          .S1(phase_accum_63__N_146[17]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_18.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_18.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_18.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_18.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_16 (.A0(phase_accum[14]), .B0(phase_inc_carrGen1[14]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[15]), .B1(phase_inc_carrGen1[15]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10961), .COUT(n10962), .S0(phase_accum_63__N_146[14]), 
          .S1(phase_accum_63__N_146[15]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_16.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_16.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_16.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_16.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_14 (.A0(phase_accum[12]), .B0(phase_inc_carrGen1[12]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[13]), .B1(phase_inc_carrGen1[13]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10960), .COUT(n10961), .S0(phase_accum_63__N_146[12]), 
          .S1(phase_accum_63__N_146[13]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_14.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_14.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_14.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_14.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_12 (.A0(phase_accum[10]), .B0(phase_inc_carrGen1[10]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[11]), .B1(phase_inc_carrGen1[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10959), .COUT(n10960), .S0(phase_accum_63__N_146[10]), 
          .S1(phase_accum_63__N_146[11]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_12.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_12.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_12.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_12.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_10 (.A0(phase_accum[8]), .B0(phase_inc_carrGen1[8]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[9]), .B1(phase_inc_carrGen1[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10958), .COUT(n10959), .S0(phase_accum_63__N_146[8]), 
          .S1(phase_accum_63__N_146[9]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_10.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_10.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_10.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_10.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_8 (.A0(phase_accum[6]), .B0(phase_inc_carrGen1[6]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[7]), .B1(phase_inc_carrGen1[7]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10957), .COUT(n10958), .S0(phase_accum_63__N_146[6]), 
          .S1(phase_accum_63__N_146[7]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_8.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_8.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_8.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_8.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_6 (.A0(phase_accum[4]), .B0(phase_inc_carrGen1[4]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[5]), .B1(phase_inc_carrGen1[5]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10956), .COUT(n10957), .S0(phase_accum_63__N_146[4]), 
          .S1(phase_accum_63__N_146[5]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_6.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_6.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_6.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_6.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_4 (.A0(phase_accum[2]), .B0(phase_inc_carrGen1[2]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[3]), .B1(phase_inc_carrGen1[3]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10955), .COUT(n10956), .S0(phase_accum_63__N_146[2]), 
          .S1(phase_accum_63__N_146[3]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_4.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_4.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_4.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_4.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_2 (.A0(phase_accum[0]), .B0(phase_inc_carrGen1[0]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[1]), .B1(phase_inc_carrGen1[1]), 
          .C1(GND_net), .D1(GND_net), .COUT(n10955), .S1(phase_accum_63__N_146[1]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_2.INIT0 = 16'h7000;
    defparam phase_accum_63__I_0_12_2.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_2.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_2.INJECT1_1 = "NO";
    LUT4 phase_accum_63__I_0_13_1_lut (.A(\phase_accum[63] ), .Z(sinGen_c)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(32[18:56])
    defparam phase_accum_63__I_0_13_1_lut.init = 16'h5555;
    LUT4 i4905_2_lut (.A(phase_accum[0]), .B(phase_inc_carrGen1[0]), .Z(phase_accum_63__N_146[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4905_2_lut.init = 16'h6666;
    
endmodule
//
// Verilog Description of module \CIC(width=72,decimation_ratio=4096) 
//

module \CIC(width=72,decimation_ratio=4096)  (osc_clk, MixerOutSin, GND_net, 
            CIC1_out_clkSin, \CICGain[1] , \CICGain[0] , \CIC1_outSin[0] , 
            n63, \d_out_11__N_1819[2] , n64, \d_out_11__N_1819[3] , 
            n65, \d_out_11__N_1819[4] , n66, \d_out_11__N_1819[5] , 
            n67, \d_out_11__N_1819[6] , n68, \d_out_11__N_1819[7] , 
            \d10[68] , \d_out_11__N_1819[8] , n70, \d_out_11__N_1819[9] , 
            \d10[71] , \d_out_11__N_1819[11] , \d10[65] , \d10[66] , 
            \d10[63] , \d10[64] , \d10[61] , \d10[62] , n61, \d10[59] , 
            n62, \d10[60] , \CIC1_outSin[1] , \CIC1_outSin[2] , \CIC1_outSin[3] , 
            \CIC1_outSin[4] , \CIC1_outSin[5] , MYLED_c_0, MYLED_c_1, 
            MYLED_c_2, MYLED_c_3, MYLED_c_4, MYLED_c_5, \d10[67] , 
            \d10[69] , \d10[70] , \d_out_11__N_1819[10] ) /* synthesis syn_module_defined=1 */ ;
    input osc_clk;
    input [11:0]MixerOutSin;
    input GND_net;
    output CIC1_out_clkSin;
    input \CICGain[1] ;
    input \CICGain[0] ;
    output \CIC1_outSin[0] ;
    input n63;
    output \d_out_11__N_1819[2] ;
    input n64;
    output \d_out_11__N_1819[3] ;
    input n65;
    output \d_out_11__N_1819[4] ;
    input n66;
    output \d_out_11__N_1819[5] ;
    input n67;
    output \d_out_11__N_1819[6] ;
    input n68;
    output \d_out_11__N_1819[7] ;
    input \d10[68] ;
    output \d_out_11__N_1819[8] ;
    input n70;
    output \d_out_11__N_1819[9] ;
    input \d10[71] ;
    output \d_out_11__N_1819[11] ;
    input \d10[65] ;
    input \d10[66] ;
    input \d10[63] ;
    input \d10[64] ;
    input \d10[61] ;
    input \d10[62] ;
    input n61;
    input \d10[59] ;
    input n62;
    input \d10[60] ;
    output \CIC1_outSin[1] ;
    output \CIC1_outSin[2] ;
    output \CIC1_outSin[3] ;
    output \CIC1_outSin[4] ;
    output \CIC1_outSin[5] ;
    output MYLED_c_0;
    output MYLED_c_1;
    output MYLED_c_2;
    output MYLED_c_3;
    output MYLED_c_4;
    output MYLED_c_5;
    input \d10[67] ;
    input \d10[69] ;
    input \d10[70] ;
    output \d_out_11__N_1819[10] ;
    
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(71[8:15])
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(82[6:21])
    wire [71:0]d_d_tmp;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(30[33:40])
    
    wire osc_clk_enable_75;
    wire [71:0]d_tmp;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(30[26:31])
    
    wire n12263;
    wire [71:0]d1;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(35[26:28])
    
    wire n4276;
    wire [35:0]n4277;
    wire [71:0]d1_71__N_418;
    
    wire n12264, osc_clk_enable_1458;
    wire [71:0]d5;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(39[26:28])
    wire [71:0]d2;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(36[26:28])
    wire [71:0]d2_71__N_490;
    
    wire n11839;
    wire [71:0]d9;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(46[26:28])
    wire [71:0]d_d9;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(46[30:34])
    wire [35:0]n5949;
    
    wire n11840;
    wire [71:0]d3;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(37[26:28])
    wire [71:0]d3_71__N_562;
    wire [71:0]d4;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(38[26:28])
    wire [71:0]d4_71__N_634;
    wire [71:0]d5_71__N_706;
    wire [71:0]d6;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(43[26:28])
    wire [71:0]d6_71__N_1459;
    wire [71:0]d_d6;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(43[30:34])
    
    wire n11831, n11832, d_clk_tmp, n8356, v_comb;
    wire [71:0]d7;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(44[26:28])
    wire [71:0]d7_71__N_1531;
    wire [35:0]n5987;
    
    wire n5948;
    wire [71:0]d10_71__N_1747;
    
    wire n63_c, n131;
    wire [71:0]d_out_11__N_1819;
    
    wire n64_c, n132;
    wire [71:0]d_d7;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(44[30:34])
    wire [71:0]d8;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(45[26:28])
    wire [71:0]d8_71__N_1603;
    wire [71:0]d_d8;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(45[30:34])
    wire [71:0]d9_71__N_1675;
    wire [15:0]count;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(50[14:19])
    wire [15:0]count_15__N_1442;
    
    wire n65_c, n133, n66_c, n134;
    wire [71:0]d10;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(47[26:29])
    
    wire n62_c, n13488, n135, n68_c, n136, n137, n70_c, n138, 
        n11628, n11629, n140, n12262, n12261, n12260, n12259, 
        n12258, n12257, n12256, n12255, n12254, n12253, osc_clk_enable_547, 
        n11627, n131_adj_2488, n13401, n11626, n11625, n11624, n132_adj_2491, 
        n13127, n133_adj_2494, n134_adj_2497, n135_adj_2499, n136_adj_2502, 
        n137_adj_2504, n140_adj_2508, n138_adj_2509, n11880;
    wire [35:0]n5797;
    
    wire n11879, n11878, n11877, n11876, n11875, n11874, n11873, 
        n11872, n11871, n11870, n11869, n11868, osc_clk_enable_147, 
        n11830, n11829, n11828, n11827, n11826, n11825, n11824, 
        n11823, n11822, n11821, n11838, n11820, n11819, n11818, 
        n11817, n11816, n11867, n11866, n11815, n11865, n11814, 
        n11864, n11863, n11813, osc_clk_enable_297, n11861, n5796, 
        n11860, n11859, n11858, n11857, n11856, n11855, n11854, 
        n11812, n11853, n11811, n11852, n11851, n11850, n11849, 
        n11848, n11847, n11846, n11845, n11810, n11809, n11808, 
        n11807, n11806, osc_clk_enable_247, n12248;
    wire [35:0]n4429;
    
    wire n11805, n61_adj_2521, n11837, n11836, n8376;
    wire [15:0]n375;
    
    wire d_clk_tmp_N_1831, n13125, n13, n13113, n13505, n12247, 
        n12246, n12245, n12244, n12243, n12242, n12241, n12240, 
        n12239, n12238, n12237, n12236, n12235, n12234, osc_clk_enable_197, 
        osc_clk_enable_347, osc_clk_enable_397, osc_clk_enable_447, osc_clk_enable_497, 
        osc_clk_enable_597, osc_clk_enable_647, osc_clk_enable_697, n12233, 
        n12232, n12229, n4428, n12228, n12227, n12226, n12225, 
        n12224, n12223, n12222, n12221, n12220, n31, n12219, n12218, 
        n12217, n12216, n12215, n12214, n12213, n12212, n11844, 
        n11835, n11834, n11833, n12207;
    wire [35:0]n4581;
    
    wire n12206, n11427;
    wire [35:0]n6861;
    
    wire n11426, n11425, n11424, n11423, n11422, n11421, n11420, 
        n11419, n11418, n11417, n11416, n11415, n11414, n11413, 
        n11412, n11411, n11410, n11408, n6860, n11407, n11406, 
        n11405, n11404, n11403, n11402, n11401, n11400, n11399, 
        n11398, n11397, n11396, n11395, n11394, n11393, n11392, 
        n11391, n11387;
    wire [35:0]n7013;
    
    wire n11386, n11385, n11384, n11383, n11382, n11381, n11380, 
        n11379, n11378, n11377, n11376, n11375, n11374, n11373, 
        n11372, n11371, n11370, n11368, n7012, n11367, n11366, 
        n11365, n11364, n11363, n11362, n11361, n11360, n11359, 
        n11358, n11357, n11356, n11355, n11354, n11353, n11352, 
        n11351, n11262, n4124, n11261, n11260, n11259, n11258, 
        n11257, n11256, n11255, n11254, n11253, n11252, n11251, 
        n11250, n11249, n11248, n11247, n11246, n11245, n11223, 
        n11222, n11221, n11220, n11219, n11218, n11217, n11216, 
        n11215, n11214, n11213, n11212, n11211, n11210, n11209, 
        n11208, n11207, n11206, n11099, n11098, n11097, n11096, 
        n11095, n11094, n11093, n11092, n11072, n4884, n11071, 
        n11070, n11069, n11068, n11067, n11066, n11065, n11064, 
        n11063, n11062, n11061, n11060, n11059, n11058, n11057, 
        n11056, n11055, n11053, n4732, n11052, n11051, n11050, 
        n11049, n11048, n11047, n11046, n11045, n11044, n11043, 
        n11042, n11041, n11040, n11039, n11038, n11037, n11036, 
        n11034, n4580, n11033, n11032, n11031, n11030, n11029, 
        n11028, n11027, n11026, n11025, n11024, n11023, n11022, 
        n11021, n11020, n11019, n11018, n11017, n11015, n11014, 
        n11013, n11012, n11011, n11010, n11009, n11008, n11007, 
        n11006, n11005, n11004, n11003, n11002, n11001, n11000, 
        n10999, n10998, n10953, n10952, n10951, n10950, n10949, 
        n10948, n10947, n10946, n10945, n10944, n10943, n10942, 
        n10941, n10940, n10939, n10938, n10937, n10936, n12424, 
        n12423, n12422, n11777, n11776, n11775, n11774, n11773, 
        n11772, n11771, n11770, n11769, n11768, n11767, n11766, 
        n11765, n11764, n11763, n11762, n11761, n11760, n11641, 
        n11640, n11639, n11638, n11637, n11636, n11635, n11634, 
        n11633, n11632, n11631, n11630, n12421, n12420, n12419, 
        n12418, n7, n12793, n12417, n12416, n12415, n12414, n12413, 
        n12412, n12411, n12410, n12409, n12408, n12407, n12205, 
        n12204, n12203, n12202, n12201, n12200, n12199, n12198, 
        n12197, n12196, n12195, n12194, n12193, n12192, n12191, 
        n12188, n12187, n12186, n12185, n12184, n12183, n12182, 
        n12181, n12180, n12179, n12178, n12177, n12176, n12175, 
        n12174, n12173, n12172, n12171, n12166;
    wire [35:0]n4733;
    
    wire n12165, n12164, n12163, n12162, n12161, n12160, n12159, 
        n12158, n12157, n12156, n12155, n12154, n12153, n12152, 
        n12151, n12150, n13391, n13395, n13394, n13398, n13397, 
        n13400, n12147, n12146, n12330;
    wire [35:0]n4125;
    
    wire n12329, n12145, n12328, n12327, n12326, n12144, n12143, 
        n12325, n12324, n12323, n12142, n12322, n12321, n12320, 
        n12141, n12140, n12319, n12318, n12317, n12316, n12315, 
        n12314, n21, n19, n15, n16, n12313, n12311, n12310, 
        n12309, n12308, n12307, n12306, n12305, n12304, n12303, 
        n12139, n12302, n12301, n12300, n12299, n12298, n12297, 
        n12138, n12296, n12295, n12294, n12289, n12137, n12288, 
        n12287, n12286, n12285, n12284, n12283, n12282, n12281, 
        n12280, n12279, n12278, n12277, n12276, n12275, n12136, 
        n12135, n13392, n12134, n12133, n12132, n12131, n12130, 
        n12125;
    wire [35:0]n4885;
    
    wire n12124, n12123, n12122, n12121, n12120, n12119, n12118, 
        n12117, n12116, n12115, n12114, n12113, n12112, n12111, 
        n12110, n12109, n12274, n12273, n12106, n12105, n12104, 
        n12103, n12102, n12101, n12100, n12099, n12098, n12097, 
        n12096, n12095, n12094, n12093, n12092, n12091, n12090, 
        n12089, n12270, n12269, n12268, n12267, n12266, n12265;
    
    FD1P3AX d_d_tmp_i0_i0 (.D(d_tmp[0]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i0.GSR = "ENABLED";
    CCU2D add_1045_23 (.A0(d1[56]), .B0(n4276), .C0(n4277[20]), .D0(MixerOutSin[11]), 
          .A1(d1[57]), .B1(n4276), .C1(n4277[21]), .D1(MixerOutSin[11]), 
          .CIN(n12263), .COUT(n12264), .S0(d1_71__N_418[56]), .S1(d1_71__N_418[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1045_23.INIT0 = 16'h74b8;
    defparam add_1045_23.INIT1 = 16'h74b8;
    defparam add_1045_23.INJECT1_0 = "NO";
    defparam add_1045_23.INJECT1_1 = "NO";
    FD1P3AX d_tmp_i0_i10 (.D(d5[10]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i9 (.D(d5[9]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i9.GSR = "ENABLED";
    FD1S3AX d2_i0 (.D(d2_71__N_490[0]), .CK(osc_clk), .Q(d2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i0.GSR = "ENABLED";
    CCU2D add_1099_35 (.A0(d9[69]), .B0(d_d9[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[70]), .B1(d_d9[70]), .C1(GND_net), .D1(GND_net), .CIN(n11839), 
          .COUT(n11840), .S0(n5949[33]), .S1(n5949[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1099_35.INIT0 = 16'h5999;
    defparam add_1099_35.INIT1 = 16'h5999;
    defparam add_1099_35.INJECT1_0 = "NO";
    defparam add_1099_35.INJECT1_1 = "NO";
    FD1S3AX d3_i0 (.D(d3_71__N_562[0]), .CK(osc_clk), .Q(d3[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i0.GSR = "ENABLED";
    FD1S3AX d4_i0 (.D(d4_71__N_634[0]), .CK(osc_clk), .Q(d4[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i0.GSR = "ENABLED";
    FD1S3AX d5_i0 (.D(d5_71__N_706[0]), .CK(osc_clk), .Q(d5[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i0.GSR = "ENABLED";
    FD1P3AX d6_i0_i0 (.D(d6_71__N_1459[0]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i0 (.D(d6[0]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i0.GSR = "ENABLED";
    CCU2D add_1099_19 (.A0(d9[53]), .B0(d_d9[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[54]), .B1(d_d9[54]), .C1(GND_net), .D1(GND_net), .CIN(n11831), 
          .COUT(n11832));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1099_19.INIT0 = 16'h5999;
    defparam add_1099_19.INIT1 = 16'h5999;
    defparam add_1099_19.INJECT1_0 = "NO";
    defparam add_1099_19.INJECT1_1 = "NO";
    FD1S3JX d_clk_tmp_65 (.D(n8356), .CK(osc_clk), .PD(osc_clk_enable_1458), 
            .Q(d_clk_tmp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_clk_tmp_65.GSR = "ENABLED";
    FD1S3AX v_comb_66 (.D(osc_clk_enable_1458), .CK(osc_clk), .Q(v_comb)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66.GSR = "ENABLED";
    FD1S3AX d_clk_67 (.D(d_clk_tmp), .CK(osc_clk), .Q(CIC1_out_clkSin)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_clk_67.GSR = "ENABLED";
    FD1P3AX d7_i0_i0 (.D(d7_71__N_1531[0]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i0.GSR = "ENABLED";
    LUT4 mux_1237_i2_3_lut (.A(n5949[21]), .B(n5987[21]), .C(n5948), .Z(d10_71__N_1747[57])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1237_i2_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i203_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63_c), .D(n131), .Z(d_out_11__N_1819[2])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i203_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i204_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64_c), .D(n132), .Z(d_out_11__N_1819[3])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i204_3_lut_4_lut.init = 16'hfe10;
    FD1P3AX d_d7_i0_i0 (.D(d7[0]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d8_i0_i0 (.D(d8_71__N_1603[0]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i0 (.D(d8[0]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d9_i0_i0 (.D(d9_71__N_1675[0]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i0 (.D(d9[0]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_out_i0_i0 (.D(d_out_11__N_1819[0]), .SP(osc_clk_enable_75), 
            .CK(osc_clk), .Q(\CIC1_outSin[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i0.GSR = "ENABLED";
    FD1S3AX d1_i0 (.D(d1_71__N_418[0]), .CK(osc_clk), .Q(d1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i0.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i8 (.D(d5[8]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i8.GSR = "ENABLED";
    FD1S3IX count__i0 (.D(count_15__N_1442[0]), .CK(osc_clk), .CD(osc_clk_enable_1458), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i0.GSR = "ENABLED";
    LUT4 shift_right_31_i205_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65_c), .D(n133), .Z(d_out_11__N_1819[4])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i205_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i206_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66_c), .D(n134), .Z(d_out_11__N_1819[5])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i206_3_lut_4_lut.init = 16'hfe10;
    FD1P3AX d_tmp_i0_i7 (.D(d5[7]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i7.GSR = "ENABLED";
    LUT4 shift_right_31_i62_3_lut (.A(d10[61]), .B(d10[62]), .C(\CICGain[0] ), 
         .Z(n62_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i62_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i207_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n13488), .D(n135), .Z(d_out_11__N_1819[6])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i207_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i208_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n68_c), .D(n136), .Z(d_out_11__N_1819[7])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i208_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1237_i3_3_lut (.A(n5949[22]), .B(n5987[22]), .C(n5948), .Z(d10_71__N_1747[58])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1237_i3_3_lut.init = 16'hcaca;
    FD1P3AX d_tmp_i0_i6 (.D(d5[6]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i5 (.D(d5[5]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i5.GSR = "ENABLED";
    LUT4 shift_right_31_i141_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n137), .D(d10[68]), .Z(d_out_11__N_1819[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i141_3_lut_4_lut.init = 16'hf1e0;
    LUT4 shift_right_31_i210_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n70_c), .D(n138), .Z(d_out_11__N_1819[9])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i210_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i63_3_lut (.A(d10[62]), .B(d10[63]), .C(\CICGain[0] ), 
         .Z(n63_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i63_3_lut.init = 16'hcaca;
    FD1P3AX d_tmp_i0_i4 (.D(d5[4]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i4.GSR = "ENABLED";
    LUT4 mux_1237_i4_3_lut (.A(n5949[23]), .B(n5987[23]), .C(n5948), .Z(d10_71__N_1747[59])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1237_i4_3_lut.init = 16'hcaca;
    CCU2D add_1098_11 (.A0(d9[9]), .B0(d_d9[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[10]), .B1(d_d9[10]), .C1(GND_net), .D1(GND_net), .CIN(n11628), 
          .COUT(n11629));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1098_11.INIT0 = 16'h5999;
    defparam add_1098_11.INIT1 = 16'h5999;
    defparam add_1098_11.INJECT1_0 = "NO";
    defparam add_1098_11.INJECT1_1 = "NO";
    LUT4 shift_right_31_i212_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(d10[71]), .D(n140), .Z(d_out_11__N_1819[11])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i212_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_1045_21 (.A0(d1[54]), .B0(n4276), .C0(n4277[18]), .D0(MixerOutSin[11]), 
          .A1(d1[55]), .B1(n4276), .C1(n4277[19]), .D1(MixerOutSin[11]), 
          .CIN(n12262), .COUT(n12263), .S0(d1_71__N_418[54]), .S1(d1_71__N_418[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1045_21.INIT0 = 16'h74b8;
    defparam add_1045_21.INIT1 = 16'h74b8;
    defparam add_1045_21.INJECT1_0 = "NO";
    defparam add_1045_21.INJECT1_1 = "NO";
    CCU2D add_1045_19 (.A0(d1[52]), .B0(n4276), .C0(n4277[16]), .D0(MixerOutSin[11]), 
          .A1(d1[53]), .B1(n4276), .C1(n4277[17]), .D1(MixerOutSin[11]), 
          .CIN(n12261), .COUT(n12262), .S0(d1_71__N_418[52]), .S1(d1_71__N_418[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1045_19.INIT0 = 16'h74b8;
    defparam add_1045_19.INIT1 = 16'h74b8;
    defparam add_1045_19.INJECT1_0 = "NO";
    defparam add_1045_19.INJECT1_1 = "NO";
    CCU2D add_1045_17 (.A0(d1[50]), .B0(n4276), .C0(n4277[14]), .D0(MixerOutSin[11]), 
          .A1(d1[51]), .B1(n4276), .C1(n4277[15]), .D1(MixerOutSin[11]), 
          .CIN(n12260), .COUT(n12261), .S0(d1_71__N_418[50]), .S1(d1_71__N_418[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1045_17.INIT0 = 16'h74b8;
    defparam add_1045_17.INIT1 = 16'h74b8;
    defparam add_1045_17.INJECT1_0 = "NO";
    defparam add_1045_17.INJECT1_1 = "NO";
    CCU2D add_1045_15 (.A0(d1[48]), .B0(n4276), .C0(n4277[12]), .D0(MixerOutSin[11]), 
          .A1(d1[49]), .B1(n4276), .C1(n4277[13]), .D1(MixerOutSin[11]), 
          .CIN(n12259), .COUT(n12260), .S0(d1_71__N_418[48]), .S1(d1_71__N_418[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1045_15.INIT0 = 16'h74b8;
    defparam add_1045_15.INIT1 = 16'h74b8;
    defparam add_1045_15.INJECT1_0 = "NO";
    defparam add_1045_15.INJECT1_1 = "NO";
    CCU2D add_1045_13 (.A0(d1[46]), .B0(n4276), .C0(n4277[10]), .D0(MixerOutSin[11]), 
          .A1(d1[47]), .B1(n4276), .C1(n4277[11]), .D1(MixerOutSin[11]), 
          .CIN(n12258), .COUT(n12259), .S0(d1_71__N_418[46]), .S1(d1_71__N_418[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1045_13.INIT0 = 16'h74b8;
    defparam add_1045_13.INIT1 = 16'h74b8;
    defparam add_1045_13.INJECT1_0 = "NO";
    defparam add_1045_13.INJECT1_1 = "NO";
    CCU2D add_1045_11 (.A0(d1[44]), .B0(n4276), .C0(n4277[8]), .D0(MixerOutSin[11]), 
          .A1(d1[45]), .B1(n4276), .C1(n4277[9]), .D1(MixerOutSin[11]), 
          .CIN(n12257), .COUT(n12258), .S0(d1_71__N_418[44]), .S1(d1_71__N_418[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1045_11.INIT0 = 16'h74b8;
    defparam add_1045_11.INIT1 = 16'h74b8;
    defparam add_1045_11.INJECT1_0 = "NO";
    defparam add_1045_11.INJECT1_1 = "NO";
    CCU2D add_1045_9 (.A0(d1[42]), .B0(n4276), .C0(n4277[6]), .D0(MixerOutSin[11]), 
          .A1(d1[43]), .B1(n4276), .C1(n4277[7]), .D1(MixerOutSin[11]), 
          .CIN(n12256), .COUT(n12257), .S0(d1_71__N_418[42]), .S1(d1_71__N_418[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1045_9.INIT0 = 16'h74b8;
    defparam add_1045_9.INIT1 = 16'h74b8;
    defparam add_1045_9.INJECT1_0 = "NO";
    defparam add_1045_9.INJECT1_1 = "NO";
    CCU2D add_1045_7 (.A0(d1[40]), .B0(n4276), .C0(n4277[4]), .D0(MixerOutSin[11]), 
          .A1(d1[41]), .B1(n4276), .C1(n4277[5]), .D1(MixerOutSin[11]), 
          .CIN(n12255), .COUT(n12256), .S0(d1_71__N_418[40]), .S1(d1_71__N_418[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1045_7.INIT0 = 16'h74b8;
    defparam add_1045_7.INIT1 = 16'h74b8;
    defparam add_1045_7.INJECT1_0 = "NO";
    defparam add_1045_7.INJECT1_1 = "NO";
    CCU2D add_1045_5 (.A0(d1[38]), .B0(n4276), .C0(n4277[2]), .D0(MixerOutSin[11]), 
          .A1(d1[39]), .B1(n4276), .C1(n4277[3]), .D1(MixerOutSin[11]), 
          .CIN(n12254), .COUT(n12255), .S0(d1_71__N_418[38]), .S1(d1_71__N_418[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1045_5.INIT0 = 16'h74b8;
    defparam add_1045_5.INIT1 = 16'h74b8;
    defparam add_1045_5.INJECT1_0 = "NO";
    defparam add_1045_5.INJECT1_1 = "NO";
    CCU2D add_1045_3 (.A0(d1[36]), .B0(n4276), .C0(n4277[0]), .D0(MixerOutSin[11]), 
          .A1(d1[37]), .B1(n4276), .C1(n4277[1]), .D1(MixerOutSin[11]), 
          .CIN(n12253), .COUT(n12254), .S0(d1_71__N_418[36]), .S1(d1_71__N_418[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1045_3.INIT0 = 16'h74b8;
    defparam add_1045_3.INIT1 = 16'h74b8;
    defparam add_1045_3.INJECT1_0 = "NO";
    defparam add_1045_3.INJECT1_1 = "NO";
    CCU2D add_1045_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n4276), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n12253));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1045_1.INIT0 = 16'hF000;
    defparam add_1045_1.INIT1 = 16'h0555;
    defparam add_1045_1.INJECT1_0 = "NO";
    defparam add_1045_1.INJECT1_1 = "NO";
    FD1S3AX v_comb_66_rep_91 (.D(osc_clk_enable_1458), .CK(osc_clk), .Q(osc_clk_enable_547)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_91.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i3 (.D(d5[3]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i3.GSR = "ENABLED";
    CCU2D add_1098_9 (.A0(d9[7]), .B0(d_d9[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[8]), .B1(d_d9[8]), .C1(GND_net), .D1(GND_net), .CIN(n11627), 
          .COUT(n11628));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1098_9.INIT0 = 16'h5999;
    defparam add_1098_9.INIT1 = 16'h5999;
    defparam add_1098_9.INJECT1_0 = "NO";
    defparam add_1098_9.INJECT1_1 = "NO";
    LUT4 shift_right_31_i203_3_lut_4_lut_adj_25 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63), .D(n131_adj_2488), .Z(\d_out_11__N_1819[2] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i203_3_lut_4_lut_adj_25.init = 16'hfe10;
    LUT4 i11_3_lut_4_lut_then_3_lut_3_lut (.A(d10[67]), .B(\CICGain[0] ), 
         .C(d10[68]), .Z(n13401)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam i11_3_lut_4_lut_then_3_lut_3_lut.init = 16'hb8b8;
    LUT4 mux_1237_i5_3_lut (.A(n5949[24]), .B(n5987[24]), .C(n5948), .Z(d10_71__N_1747[60])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1237_i5_3_lut.init = 16'hcaca;
    CCU2D add_1098_7 (.A0(d9[5]), .B0(d_d9[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[6]), .B1(d_d9[6]), .C1(GND_net), .D1(GND_net), .CIN(n11626), 
          .COUT(n11627));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1098_7.INIT0 = 16'h5999;
    defparam add_1098_7.INIT1 = 16'h5999;
    defparam add_1098_7.INJECT1_0 = "NO";
    defparam add_1098_7.INJECT1_1 = "NO";
    CCU2D add_1098_5 (.A0(d9[3]), .B0(d_d9[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[4]), .B1(d_d9[4]), .C1(GND_net), .D1(GND_net), .CIN(n11625), 
          .COUT(n11626));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1098_5.INIT0 = 16'h5999;
    defparam add_1098_5.INIT1 = 16'h5999;
    defparam add_1098_5.INJECT1_0 = "NO";
    defparam add_1098_5.INJECT1_1 = "NO";
    CCU2D add_1098_3 (.A0(d9[1]), .B0(d_d9[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[2]), .B1(d_d9[2]), .C1(GND_net), .D1(GND_net), .CIN(n11624), 
          .COUT(n11625));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1098_3.INIT0 = 16'h5999;
    defparam add_1098_3.INIT1 = 16'h5999;
    defparam add_1098_3.INJECT1_0 = "NO";
    defparam add_1098_3.INJECT1_1 = "NO";
    CCU2D add_1098_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d9[0]), .B1(d_d9[0]), .C1(GND_net), .D1(GND_net), .COUT(n11624));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1098_1.INIT0 = 16'h0000;
    defparam add_1098_1.INIT1 = 16'h5999;
    defparam add_1098_1.INJECT1_0 = "NO";
    defparam add_1098_1.INJECT1_1 = "NO";
    LUT4 shift_right_31_i204_3_lut_4_lut_adj_26 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64), .D(n132_adj_2491), .Z(\d_out_11__N_1819[3] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i204_3_lut_4_lut_adj_26.init = 16'hfe10;
    FD1P3AX d_tmp_i0_i2 (.D(d5[2]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i2.GSR = "ENABLED";
    LUT4 i5659_4_lut (.A(count[5]), .B(count[4]), .C(count[9]), .D(count[7]), 
         .Z(n13127)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5659_4_lut.init = 16'h8000;
    LUT4 shift_right_31_i205_3_lut_4_lut_adj_27 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65), .D(n133_adj_2494), .Z(\d_out_11__N_1819[4] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i205_3_lut_4_lut_adj_27.init = 16'hfe10;
    LUT4 shift_right_31_i206_3_lut_4_lut_adj_28 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66), .D(n134_adj_2497), .Z(\d_out_11__N_1819[5] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i206_3_lut_4_lut_adj_28.init = 16'hfe10;
    LUT4 shift_right_31_i207_3_lut_4_lut_adj_29 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n67), .D(n135_adj_2499), .Z(\d_out_11__N_1819[6] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i207_3_lut_4_lut_adj_29.init = 16'hfe10;
    LUT4 shift_right_31_i208_3_lut_4_lut_adj_30 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n68), .D(n136_adj_2502), .Z(\d_out_11__N_1819[7] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i208_3_lut_4_lut_adj_30.init = 16'hfe10;
    LUT4 shift_right_31_i141_3_lut_4_lut_adj_31 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n137_adj_2504), .D(\d10[68] ), .Z(\d_out_11__N_1819[8] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i141_3_lut_4_lut_adj_31.init = 16'hf1e0;
    LUT4 shift_right_31_i140_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n70), .D(\d10[68] ), .Z(n140_adj_2508)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i140_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i210_3_lut_4_lut_adj_32 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n70), .D(n138_adj_2509), .Z(\d_out_11__N_1819[9] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i210_3_lut_4_lut_adj_32.init = 16'hfe10;
    LUT4 shift_right_31_i64_3_lut (.A(d10[63]), .B(d10[64]), .C(\CICGain[0] ), 
         .Z(n64_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i64_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i212_3_lut_4_lut_adj_33 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(\d10[71] ), .D(n140_adj_2508), .Z(\d_out_11__N_1819[11] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i212_3_lut_4_lut_adj_33.init = 16'hfe10;
    LUT4 shift_right_31_i137_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n67), .D(\d10[65] ), .Z(n137_adj_2504)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i137_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i138_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n68), .D(\d10[66] ), .Z(n138_adj_2509)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i138_3_lut_4_lut.init = 16'hf960;
    FD1P3AX d_tmp_i0_i1 (.D(d5[1]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i11 (.D(d5[11]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i22 (.D(d5[22]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i22.GSR = "ENABLED";
    LUT4 shift_right_31_i65_3_lut (.A(d10[64]), .B(d10[65]), .C(\CICGain[0] ), 
         .Z(n65_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i65_3_lut.init = 16'hcaca;
    LUT4 mux_1237_i6_3_lut (.A(n5949[25]), .B(n5987[25]), .C(n5948), .Z(d10_71__N_1747[61])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1237_i6_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i135_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65), .D(\d10[63] ), .Z(n135_adj_2499)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i135_3_lut_4_lut.init = 16'hf960;
    CCU2D add_1094_37 (.A0(d8[71]), .B0(d_d8[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11880), 
          .S0(n5797[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1094_37.INIT0 = 16'h5999;
    defparam add_1094_37.INIT1 = 16'h0000;
    defparam add_1094_37.INJECT1_0 = "NO";
    defparam add_1094_37.INJECT1_1 = "NO";
    CCU2D add_1094_35 (.A0(d8[69]), .B0(d_d8[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[70]), .B1(d_d8[70]), .C1(GND_net), .D1(GND_net), .CIN(n11879), 
          .COUT(n11880), .S0(n5797[33]), .S1(n5797[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1094_35.INIT0 = 16'h5999;
    defparam add_1094_35.INIT1 = 16'h5999;
    defparam add_1094_35.INJECT1_0 = "NO";
    defparam add_1094_35.INJECT1_1 = "NO";
    CCU2D add_1094_33 (.A0(d8[67]), .B0(d_d8[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[68]), .B1(d_d8[68]), .C1(GND_net), .D1(GND_net), .CIN(n11878), 
          .COUT(n11879), .S0(n5797[31]), .S1(n5797[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1094_33.INIT0 = 16'h5999;
    defparam add_1094_33.INIT1 = 16'h5999;
    defparam add_1094_33.INJECT1_0 = "NO";
    defparam add_1094_33.INJECT1_1 = "NO";
    CCU2D add_1094_31 (.A0(d8[65]), .B0(d_d8[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[66]), .B1(d_d8[66]), .C1(GND_net), .D1(GND_net), .CIN(n11877), 
          .COUT(n11878), .S0(n5797[29]), .S1(n5797[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1094_31.INIT0 = 16'h5999;
    defparam add_1094_31.INIT1 = 16'h5999;
    defparam add_1094_31.INJECT1_0 = "NO";
    defparam add_1094_31.INJECT1_1 = "NO";
    CCU2D add_1094_29 (.A0(d8[63]), .B0(d_d8[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[64]), .B1(d_d8[64]), .C1(GND_net), .D1(GND_net), .CIN(n11876), 
          .COUT(n11877), .S0(n5797[27]), .S1(n5797[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1094_29.INIT0 = 16'h5999;
    defparam add_1094_29.INIT1 = 16'h5999;
    defparam add_1094_29.INJECT1_0 = "NO";
    defparam add_1094_29.INJECT1_1 = "NO";
    CCU2D add_1094_27 (.A0(d8[61]), .B0(d_d8[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[62]), .B1(d_d8[62]), .C1(GND_net), .D1(GND_net), .CIN(n11875), 
          .COUT(n11876), .S0(n5797[25]), .S1(n5797[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1094_27.INIT0 = 16'h5999;
    defparam add_1094_27.INIT1 = 16'h5999;
    defparam add_1094_27.INJECT1_0 = "NO";
    defparam add_1094_27.INJECT1_1 = "NO";
    CCU2D add_1094_25 (.A0(d8[59]), .B0(d_d8[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[60]), .B1(d_d8[60]), .C1(GND_net), .D1(GND_net), .CIN(n11874), 
          .COUT(n11875), .S0(n5797[23]), .S1(n5797[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1094_25.INIT0 = 16'h5999;
    defparam add_1094_25.INIT1 = 16'h5999;
    defparam add_1094_25.INJECT1_0 = "NO";
    defparam add_1094_25.INJECT1_1 = "NO";
    CCU2D add_1094_23 (.A0(d8[57]), .B0(d_d8[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[58]), .B1(d_d8[58]), .C1(GND_net), .D1(GND_net), .CIN(n11873), 
          .COUT(n11874), .S0(n5797[21]), .S1(n5797[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1094_23.INIT0 = 16'h5999;
    defparam add_1094_23.INIT1 = 16'h5999;
    defparam add_1094_23.INJECT1_0 = "NO";
    defparam add_1094_23.INJECT1_1 = "NO";
    CCU2D add_1094_21 (.A0(d8[55]), .B0(d_d8[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[56]), .B1(d_d8[56]), .C1(GND_net), .D1(GND_net), .CIN(n11872), 
          .COUT(n11873), .S0(n5797[19]), .S1(n5797[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1094_21.INIT0 = 16'h5999;
    defparam add_1094_21.INIT1 = 16'h5999;
    defparam add_1094_21.INJECT1_0 = "NO";
    defparam add_1094_21.INJECT1_1 = "NO";
    CCU2D add_1094_19 (.A0(d8[53]), .B0(d_d8[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[54]), .B1(d_d8[54]), .C1(GND_net), .D1(GND_net), .CIN(n11871), 
          .COUT(n11872), .S0(n5797[17]), .S1(n5797[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1094_19.INIT0 = 16'h5999;
    defparam add_1094_19.INIT1 = 16'h5999;
    defparam add_1094_19.INJECT1_0 = "NO";
    defparam add_1094_19.INJECT1_1 = "NO";
    CCU2D add_1094_17 (.A0(d8[51]), .B0(d_d8[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[52]), .B1(d_d8[52]), .C1(GND_net), .D1(GND_net), .CIN(n11870), 
          .COUT(n11871), .S0(n5797[15]), .S1(n5797[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1094_17.INIT0 = 16'h5999;
    defparam add_1094_17.INIT1 = 16'h5999;
    defparam add_1094_17.INJECT1_0 = "NO";
    defparam add_1094_17.INJECT1_1 = "NO";
    CCU2D add_1094_15 (.A0(d8[49]), .B0(d_d8[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[50]), .B1(d_d8[50]), .C1(GND_net), .D1(GND_net), .CIN(n11869), 
          .COUT(n11870), .S0(n5797[13]), .S1(n5797[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1094_15.INIT0 = 16'h5999;
    defparam add_1094_15.INIT1 = 16'h5999;
    defparam add_1094_15.INJECT1_0 = "NO";
    defparam add_1094_15.INJECT1_1 = "NO";
    CCU2D add_1094_13 (.A0(d8[47]), .B0(d_d8[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[48]), .B1(d_d8[48]), .C1(GND_net), .D1(GND_net), .CIN(n11868), 
          .COUT(n11869), .S0(n5797[11]), .S1(n5797[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1094_13.INIT0 = 16'h5999;
    defparam add_1094_13.INIT1 = 16'h5999;
    defparam add_1094_13.INJECT1_0 = "NO";
    defparam add_1094_13.INJECT1_1 = "NO";
    LUT4 mux_1237_i7_3_lut (.A(n5949[26]), .B(n5987[26]), .C(n5948), .Z(d10_71__N_1747[62])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1237_i7_3_lut.init = 16'hcaca;
    FD1P3AX d_d_tmp_i0_i71 (.D(d_tmp[71]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i70 (.D(d_tmp[70]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i69 (.D(d_tmp[69]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i68 (.D(d_tmp[68]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i67 (.D(d_tmp[67]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i66 (.D(d_tmp[66]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i65 (.D(d_tmp[65]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i64 (.D(d_tmp[64]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i63 (.D(d_tmp[63]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i62 (.D(d_tmp[62]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i61 (.D(d_tmp[61]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i60 (.D(d_tmp[60]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i59 (.D(d_tmp[59]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i58 (.D(d_tmp[58]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i57 (.D(d_tmp[57]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i56 (.D(d_tmp[56]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i55 (.D(d_tmp[55]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i54 (.D(d_tmp[54]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i53 (.D(d_tmp[53]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i52 (.D(d_tmp[52]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i51 (.D(d_tmp[51]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i50 (.D(d_tmp[50]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i49 (.D(d_tmp[49]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i48 (.D(d_tmp[48]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i47 (.D(d_tmp[47]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i46 (.D(d_tmp[46]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i45 (.D(d_tmp[45]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i44 (.D(d_tmp[44]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i43 (.D(d_tmp[43]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i42 (.D(d_tmp[42]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i41 (.D(d_tmp[41]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i40 (.D(d_tmp[40]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i39 (.D(d_tmp[39]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i32 (.D(d_tmp[32]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i31 (.D(d_tmp[31]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i30 (.D(d_tmp[30]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i29 (.D(d_tmp[29]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i28 (.D(d_tmp[28]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i27 (.D(d_tmp[27]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i26 (.D(d_tmp[26]), .SP(osc_clk_enable_75), .CK(osc_clk), 
            .Q(d_d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i33 (.D(d_tmp[33]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i34 (.D(d_tmp[34]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i34.GSR = "ENABLED";
    LUT4 shift_right_31_i136_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66), .D(\d10[64] ), .Z(n136_adj_2502)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i136_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i133_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63), .D(\d10[61] ), .Z(n133_adj_2494)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i133_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i134_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64), .D(\d10[62] ), .Z(n134_adj_2497)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i134_3_lut_4_lut.init = 16'hf960;
    CCU2D add_1099_17 (.A0(d9[51]), .B0(d_d9[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[52]), .B1(d_d9[52]), .C1(GND_net), .D1(GND_net), .CIN(n11830), 
          .COUT(n11831));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1099_17.INIT0 = 16'h5999;
    defparam add_1099_17.INIT1 = 16'h5999;
    defparam add_1099_17.INJECT1_0 = "NO";
    defparam add_1099_17.INJECT1_1 = "NO";
    CCU2D add_1099_15 (.A0(d9[49]), .B0(d_d9[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[50]), .B1(d_d9[50]), .C1(GND_net), .D1(GND_net), .CIN(n11829), 
          .COUT(n11830));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1099_15.INIT0 = 16'h5999;
    defparam add_1099_15.INIT1 = 16'h5999;
    defparam add_1099_15.INJECT1_0 = "NO";
    defparam add_1099_15.INJECT1_1 = "NO";
    FD1P3AX d_d_tmp_i0_i35 (.D(d_tmp[35]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i35.GSR = "ENABLED";
    CCU2D add_1099_13 (.A0(d9[47]), .B0(d_d9[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[48]), .B1(d_d9[48]), .C1(GND_net), .D1(GND_net), .CIN(n11828), 
          .COUT(n11829));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1099_13.INIT0 = 16'h5999;
    defparam add_1099_13.INIT1 = 16'h5999;
    defparam add_1099_13.INJECT1_0 = "NO";
    defparam add_1099_13.INJECT1_1 = "NO";
    CCU2D add_1099_11 (.A0(d9[45]), .B0(d_d9[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[46]), .B1(d_d9[46]), .C1(GND_net), .D1(GND_net), .CIN(n11827), 
          .COUT(n11828));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1099_11.INIT0 = 16'h5999;
    defparam add_1099_11.INIT1 = 16'h5999;
    defparam add_1099_11.INJECT1_0 = "NO";
    defparam add_1099_11.INJECT1_1 = "NO";
    CCU2D add_1099_9 (.A0(d9[43]), .B0(d_d9[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[44]), .B1(d_d9[44]), .C1(GND_net), .D1(GND_net), .CIN(n11826), 
          .COUT(n11827));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1099_9.INIT0 = 16'h5999;
    defparam add_1099_9.INIT1 = 16'h5999;
    defparam add_1099_9.INJECT1_0 = "NO";
    defparam add_1099_9.INJECT1_1 = "NO";
    CCU2D add_1099_7 (.A0(d9[41]), .B0(d_d9[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[42]), .B1(d_d9[42]), .C1(GND_net), .D1(GND_net), .CIN(n11825), 
          .COUT(n11826));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1099_7.INIT0 = 16'h5999;
    defparam add_1099_7.INIT1 = 16'h5999;
    defparam add_1099_7.INJECT1_0 = "NO";
    defparam add_1099_7.INJECT1_1 = "NO";
    CCU2D add_1099_5 (.A0(d9[39]), .B0(d_d9[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[40]), .B1(d_d9[40]), .C1(GND_net), .D1(GND_net), .CIN(n11824), 
          .COUT(n11825));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1099_5.INIT0 = 16'h5999;
    defparam add_1099_5.INIT1 = 16'h5999;
    defparam add_1099_5.INJECT1_0 = "NO";
    defparam add_1099_5.INJECT1_1 = "NO";
    CCU2D add_1099_3 (.A0(d9[37]), .B0(d_d9[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[38]), .B1(d_d9[38]), .C1(GND_net), .D1(GND_net), .CIN(n11823), 
          .COUT(n11824));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1099_3.INIT0 = 16'h5999;
    defparam add_1099_3.INIT1 = 16'h5999;
    defparam add_1099_3.INJECT1_0 = "NO";
    defparam add_1099_3.INJECT1_1 = "NO";
    CCU2D add_1099_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d9[36]), .B1(d_d9[36]), .C1(GND_net), .D1(GND_net), .COUT(n11823));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1099_1.INIT0 = 16'hF000;
    defparam add_1099_1.INIT1 = 16'h5999;
    defparam add_1099_1.INJECT1_0 = "NO";
    defparam add_1099_1.INJECT1_1 = "NO";
    CCU2D add_1100_37 (.A0(d9[71]), .B0(d_d9[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11822), 
          .S0(n5987[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1100_37.INIT0 = 16'h5999;
    defparam add_1100_37.INIT1 = 16'h0000;
    defparam add_1100_37.INJECT1_0 = "NO";
    defparam add_1100_37.INJECT1_1 = "NO";
    CCU2D add_1100_35 (.A0(d9[69]), .B0(d_d9[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[70]), .B1(d_d9[70]), .C1(GND_net), .D1(GND_net), .CIN(n11821), 
          .COUT(n11822), .S0(n5987[33]), .S1(n5987[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1100_35.INIT0 = 16'h5999;
    defparam add_1100_35.INIT1 = 16'h5999;
    defparam add_1100_35.INJECT1_0 = "NO";
    defparam add_1100_35.INJECT1_1 = "NO";
    CCU2D add_1099_33 (.A0(d9[67]), .B0(d_d9[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[68]), .B1(d_d9[68]), .C1(GND_net), .D1(GND_net), .CIN(n11838), 
          .COUT(n11839), .S0(n5949[31]), .S1(n5949[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1099_33.INIT0 = 16'h5999;
    defparam add_1099_33.INIT1 = 16'h5999;
    defparam add_1099_33.INJECT1_0 = "NO";
    defparam add_1099_33.INJECT1_1 = "NO";
    LUT4 mux_1237_i8_3_lut (.A(n5949[27]), .B(n5987[27]), .C(n5948), .Z(d10_71__N_1747[63])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1237_i8_3_lut.init = 16'hcaca;
    CCU2D add_1100_33 (.A0(d9[67]), .B0(d_d9[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[68]), .B1(d_d9[68]), .C1(GND_net), .D1(GND_net), .CIN(n11820), 
          .COUT(n11821), .S0(n5987[31]), .S1(n5987[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1100_33.INIT0 = 16'h5999;
    defparam add_1100_33.INIT1 = 16'h5999;
    defparam add_1100_33.INJECT1_0 = "NO";
    defparam add_1100_33.INJECT1_1 = "NO";
    CCU2D add_1100_31 (.A0(d9[65]), .B0(d_d9[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[66]), .B1(d_d9[66]), .C1(GND_net), .D1(GND_net), .CIN(n11819), 
          .COUT(n11820), .S0(n5987[29]), .S1(n5987[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1100_31.INIT0 = 16'h5999;
    defparam add_1100_31.INIT1 = 16'h5999;
    defparam add_1100_31.INJECT1_0 = "NO";
    defparam add_1100_31.INJECT1_1 = "NO";
    CCU2D add_1100_29 (.A0(d9[63]), .B0(d_d9[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[64]), .B1(d_d9[64]), .C1(GND_net), .D1(GND_net), .CIN(n11818), 
          .COUT(n11819), .S0(n5987[27]), .S1(n5987[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1100_29.INIT0 = 16'h5999;
    defparam add_1100_29.INIT1 = 16'h5999;
    defparam add_1100_29.INJECT1_0 = "NO";
    defparam add_1100_29.INJECT1_1 = "NO";
    CCU2D add_1100_27 (.A0(d9[61]), .B0(d_d9[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[62]), .B1(d_d9[62]), .C1(GND_net), .D1(GND_net), .CIN(n11817), 
          .COUT(n11818), .S0(n5987[25]), .S1(n5987[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1100_27.INIT0 = 16'h5999;
    defparam add_1100_27.INIT1 = 16'h5999;
    defparam add_1100_27.INJECT1_0 = "NO";
    defparam add_1100_27.INJECT1_1 = "NO";
    CCU2D add_1100_25 (.A0(d9[59]), .B0(d_d9[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[60]), .B1(d_d9[60]), .C1(GND_net), .D1(GND_net), .CIN(n11816), 
          .COUT(n11817), .S0(n5987[23]), .S1(n5987[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1100_25.INIT0 = 16'h5999;
    defparam add_1100_25.INIT1 = 16'h5999;
    defparam add_1100_25.INJECT1_0 = "NO";
    defparam add_1100_25.INJECT1_1 = "NO";
    LUT4 shift_right_31_i131_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n61), .D(\d10[59] ), .Z(n131_adj_2488)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i131_3_lut_4_lut.init = 16'hf960;
    CCU2D add_1094_11 (.A0(d8[45]), .B0(d_d8[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[46]), .B1(d_d8[46]), .C1(GND_net), .D1(GND_net), .CIN(n11867), 
          .COUT(n11868), .S0(n5797[9]), .S1(n5797[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1094_11.INIT0 = 16'h5999;
    defparam add_1094_11.INIT1 = 16'h5999;
    defparam add_1094_11.INJECT1_0 = "NO";
    defparam add_1094_11.INJECT1_1 = "NO";
    CCU2D add_1094_9 (.A0(d8[43]), .B0(d_d8[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[44]), .B1(d_d8[44]), .C1(GND_net), .D1(GND_net), .CIN(n11866), 
          .COUT(n11867), .S0(n5797[7]), .S1(n5797[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1094_9.INIT0 = 16'h5999;
    defparam add_1094_9.INIT1 = 16'h5999;
    defparam add_1094_9.INJECT1_0 = "NO";
    defparam add_1094_9.INJECT1_1 = "NO";
    CCU2D add_1100_23 (.A0(d9[57]), .B0(d_d9[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[58]), .B1(d_d9[58]), .C1(GND_net), .D1(GND_net), .CIN(n11815), 
          .COUT(n11816), .S0(n5987[21]), .S1(n5987[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1100_23.INIT0 = 16'h5999;
    defparam add_1100_23.INIT1 = 16'h5999;
    defparam add_1100_23.INJECT1_0 = "NO";
    defparam add_1100_23.INJECT1_1 = "NO";
    LUT4 shift_right_31_i132_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n62), .D(\d10[60] ), .Z(n132_adj_2491)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i132_3_lut_4_lut.init = 16'hf960;
    CCU2D add_1094_7 (.A0(d8[41]), .B0(d_d8[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[42]), .B1(d_d8[42]), .C1(GND_net), .D1(GND_net), .CIN(n11865), 
          .COUT(n11866), .S0(n5797[5]), .S1(n5797[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1094_7.INIT0 = 16'h5999;
    defparam add_1094_7.INIT1 = 16'h5999;
    defparam add_1094_7.INJECT1_0 = "NO";
    defparam add_1094_7.INJECT1_1 = "NO";
    CCU2D add_1100_21 (.A0(d9[55]), .B0(d_d9[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[56]), .B1(d_d9[56]), .C1(GND_net), .D1(GND_net), .CIN(n11814), 
          .COUT(n11815));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1100_21.INIT0 = 16'h5999;
    defparam add_1100_21.INIT1 = 16'h5999;
    defparam add_1100_21.INJECT1_0 = "NO";
    defparam add_1100_21.INJECT1_1 = "NO";
    FD1P3AX d_d_tmp_i0_i36 (.D(d_tmp[36]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i36.GSR = "ENABLED";
    CCU2D add_1094_5 (.A0(d8[39]), .B0(d_d8[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[40]), .B1(d_d8[40]), .C1(GND_net), .D1(GND_net), .CIN(n11864), 
          .COUT(n11865), .S0(n5797[3]), .S1(n5797[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1094_5.INIT0 = 16'h5999;
    defparam add_1094_5.INIT1 = 16'h5999;
    defparam add_1094_5.INJECT1_0 = "NO";
    defparam add_1094_5.INJECT1_1 = "NO";
    CCU2D add_1094_3 (.A0(d8[37]), .B0(d_d8[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[38]), .B1(d_d8[38]), .C1(GND_net), .D1(GND_net), .CIN(n11863), 
          .COUT(n11864), .S0(n5797[1]), .S1(n5797[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1094_3.INIT0 = 16'h5999;
    defparam add_1094_3.INIT1 = 16'h5999;
    defparam add_1094_3.INJECT1_0 = "NO";
    defparam add_1094_3.INJECT1_1 = "NO";
    CCU2D add_1094_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d8[36]), .B1(d_d8[36]), .C1(GND_net), .D1(GND_net), .COUT(n11863), 
          .S1(n5797[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1094_1.INIT0 = 16'hF000;
    defparam add_1094_1.INIT1 = 16'h5999;
    defparam add_1094_1.INJECT1_0 = "NO";
    defparam add_1094_1.INJECT1_1 = "NO";
    LUT4 shift_right_31_i140_3_lut_4_lut_adj_34 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n70_c), .D(d10[68]), .Z(n140)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i140_3_lut_4_lut_adj_34.init = 16'hf960;
    LUT4 mux_1237_i9_3_lut (.A(n5949[28]), .B(n5987[28]), .C(n5948), .Z(d10_71__N_1747[64])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1237_i9_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i138_3_lut_4_lut_adj_35 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n68_c), .D(d10[66]), .Z(n138)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i138_3_lut_4_lut_adj_35.init = 16'hf960;
    CCU2D add_1100_19 (.A0(d9[53]), .B0(d_d9[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[54]), .B1(d_d9[54]), .C1(GND_net), .D1(GND_net), .CIN(n11813), 
          .COUT(n11814));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1100_19.INIT0 = 16'h5999;
    defparam add_1100_19.INIT1 = 16'h5999;
    defparam add_1100_19.INJECT1_0 = "NO";
    defparam add_1100_19.INJECT1_1 = "NO";
    LUT4 mux_1237_i10_3_lut (.A(n5949[29]), .B(n5987[29]), .C(n5948), 
         .Z(d10_71__N_1747[65])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1237_i10_3_lut.init = 16'hcaca;
    FD1S3AX v_comb_66_rep_86 (.D(osc_clk_enable_1458), .CK(osc_clk), .Q(osc_clk_enable_297)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_86.GSR = "ENABLED";
    CCU2D add_1095_37 (.A0(d_d8[70]), .B0(n5796), .C0(n5797[34]), .D0(d8[70]), 
          .A1(d_d8[71]), .B1(n5796), .C1(n5797[35]), .D1(d8[71]), .CIN(n11861), 
          .S0(d9_71__N_1675[70]), .S1(d9_71__N_1675[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1095_37.INIT0 = 16'hb874;
    defparam add_1095_37.INIT1 = 16'hb874;
    defparam add_1095_37.INJECT1_0 = "NO";
    defparam add_1095_37.INJECT1_1 = "NO";
    CCU2D add_1095_35 (.A0(d_d8[68]), .B0(n5796), .C0(n5797[32]), .D0(d8[68]), 
          .A1(d_d8[69]), .B1(n5796), .C1(n5797[33]), .D1(d8[69]), .CIN(n11860), 
          .COUT(n11861), .S0(d9_71__N_1675[68]), .S1(d9_71__N_1675[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1095_35.INIT0 = 16'hb874;
    defparam add_1095_35.INIT1 = 16'hb874;
    defparam add_1095_35.INJECT1_0 = "NO";
    defparam add_1095_35.INJECT1_1 = "NO";
    CCU2D add_1095_33 (.A0(d_d8[66]), .B0(n5796), .C0(n5797[30]), .D0(d8[66]), 
          .A1(d_d8[67]), .B1(n5796), .C1(n5797[31]), .D1(d8[67]), .CIN(n11859), 
          .COUT(n11860), .S0(d9_71__N_1675[66]), .S1(d9_71__N_1675[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1095_33.INIT0 = 16'hb874;
    defparam add_1095_33.INIT1 = 16'hb874;
    defparam add_1095_33.INJECT1_0 = "NO";
    defparam add_1095_33.INJECT1_1 = "NO";
    CCU2D add_1095_31 (.A0(d_d8[64]), .B0(n5796), .C0(n5797[28]), .D0(d8[64]), 
          .A1(d_d8[65]), .B1(n5796), .C1(n5797[29]), .D1(d8[65]), .CIN(n11858), 
          .COUT(n11859), .S0(d9_71__N_1675[64]), .S1(d9_71__N_1675[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1095_31.INIT0 = 16'hb874;
    defparam add_1095_31.INIT1 = 16'hb874;
    defparam add_1095_31.INJECT1_0 = "NO";
    defparam add_1095_31.INJECT1_1 = "NO";
    CCU2D add_1095_29 (.A0(d_d8[62]), .B0(n5796), .C0(n5797[26]), .D0(d8[62]), 
          .A1(d_d8[63]), .B1(n5796), .C1(n5797[27]), .D1(d8[63]), .CIN(n11857), 
          .COUT(n11858), .S0(d9_71__N_1675[62]), .S1(d9_71__N_1675[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1095_29.INIT0 = 16'hb874;
    defparam add_1095_29.INIT1 = 16'hb874;
    defparam add_1095_29.INJECT1_0 = "NO";
    defparam add_1095_29.INJECT1_1 = "NO";
    CCU2D add_1095_27 (.A0(d_d8[60]), .B0(n5796), .C0(n5797[24]), .D0(d8[60]), 
          .A1(d_d8[61]), .B1(n5796), .C1(n5797[25]), .D1(d8[61]), .CIN(n11856), 
          .COUT(n11857), .S0(d9_71__N_1675[60]), .S1(d9_71__N_1675[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1095_27.INIT0 = 16'hb874;
    defparam add_1095_27.INIT1 = 16'hb874;
    defparam add_1095_27.INJECT1_0 = "NO";
    defparam add_1095_27.INJECT1_1 = "NO";
    CCU2D add_1095_25 (.A0(d_d8[58]), .B0(n5796), .C0(n5797[22]), .D0(d8[58]), 
          .A1(d_d8[59]), .B1(n5796), .C1(n5797[23]), .D1(d8[59]), .CIN(n11855), 
          .COUT(n11856), .S0(d9_71__N_1675[58]), .S1(d9_71__N_1675[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1095_25.INIT0 = 16'hb874;
    defparam add_1095_25.INIT1 = 16'hb874;
    defparam add_1095_25.INJECT1_0 = "NO";
    defparam add_1095_25.INJECT1_1 = "NO";
    CCU2D add_1095_23 (.A0(d_d8[56]), .B0(n5796), .C0(n5797[20]), .D0(d8[56]), 
          .A1(d_d8[57]), .B1(n5796), .C1(n5797[21]), .D1(d8[57]), .CIN(n11854), 
          .COUT(n11855), .S0(d9_71__N_1675[56]), .S1(d9_71__N_1675[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1095_23.INIT0 = 16'hb874;
    defparam add_1095_23.INIT1 = 16'hb874;
    defparam add_1095_23.INJECT1_0 = "NO";
    defparam add_1095_23.INJECT1_1 = "NO";
    CCU2D add_1100_17 (.A0(d9[51]), .B0(d_d9[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[52]), .B1(d_d9[52]), .C1(GND_net), .D1(GND_net), .CIN(n11812), 
          .COUT(n11813));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1100_17.INIT0 = 16'h5999;
    defparam add_1100_17.INIT1 = 16'h5999;
    defparam add_1100_17.INJECT1_0 = "NO";
    defparam add_1100_17.INJECT1_1 = "NO";
    CCU2D add_1095_21 (.A0(d_d8[54]), .B0(n5796), .C0(n5797[18]), .D0(d8[54]), 
          .A1(d_d8[55]), .B1(n5796), .C1(n5797[19]), .D1(d8[55]), .CIN(n11853), 
          .COUT(n11854), .S0(d9_71__N_1675[54]), .S1(d9_71__N_1675[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1095_21.INIT0 = 16'hb874;
    defparam add_1095_21.INIT1 = 16'hb874;
    defparam add_1095_21.INJECT1_0 = "NO";
    defparam add_1095_21.INJECT1_1 = "NO";
    CCU2D add_1100_15 (.A0(d9[49]), .B0(d_d9[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[50]), .B1(d_d9[50]), .C1(GND_net), .D1(GND_net), .CIN(n11811), 
          .COUT(n11812));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1100_15.INIT0 = 16'h5999;
    defparam add_1100_15.INIT1 = 16'h5999;
    defparam add_1100_15.INJECT1_0 = "NO";
    defparam add_1100_15.INJECT1_1 = "NO";
    CCU2D add_1095_19 (.A0(d_d8[52]), .B0(n5796), .C0(n5797[16]), .D0(d8[52]), 
          .A1(d_d8[53]), .B1(n5796), .C1(n5797[17]), .D1(d8[53]), .CIN(n11852), 
          .COUT(n11853), .S0(d9_71__N_1675[52]), .S1(d9_71__N_1675[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1095_19.INIT0 = 16'hb874;
    defparam add_1095_19.INIT1 = 16'hb874;
    defparam add_1095_19.INJECT1_0 = "NO";
    defparam add_1095_19.INJECT1_1 = "NO";
    CCU2D add_1095_17 (.A0(d_d8[50]), .B0(n5796), .C0(n5797[14]), .D0(d8[50]), 
          .A1(d_d8[51]), .B1(n5796), .C1(n5797[15]), .D1(d8[51]), .CIN(n11851), 
          .COUT(n11852), .S0(d9_71__N_1675[50]), .S1(d9_71__N_1675[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1095_17.INIT0 = 16'hb874;
    defparam add_1095_17.INIT1 = 16'hb874;
    defparam add_1095_17.INJECT1_0 = "NO";
    defparam add_1095_17.INJECT1_1 = "NO";
    CCU2D add_1095_15 (.A0(d_d8[48]), .B0(n5796), .C0(n5797[12]), .D0(d8[48]), 
          .A1(d_d8[49]), .B1(n5796), .C1(n5797[13]), .D1(d8[49]), .CIN(n11850), 
          .COUT(n11851), .S0(d9_71__N_1675[48]), .S1(d9_71__N_1675[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1095_15.INIT0 = 16'hb874;
    defparam add_1095_15.INIT1 = 16'hb874;
    defparam add_1095_15.INJECT1_0 = "NO";
    defparam add_1095_15.INJECT1_1 = "NO";
    CCU2D add_1095_13 (.A0(d_d8[46]), .B0(n5796), .C0(n5797[10]), .D0(d8[46]), 
          .A1(d_d8[47]), .B1(n5796), .C1(n5797[11]), .D1(d8[47]), .CIN(n11849), 
          .COUT(n11850), .S0(d9_71__N_1675[46]), .S1(d9_71__N_1675[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1095_13.INIT0 = 16'hb874;
    defparam add_1095_13.INIT1 = 16'hb874;
    defparam add_1095_13.INJECT1_0 = "NO";
    defparam add_1095_13.INJECT1_1 = "NO";
    CCU2D add_1095_11 (.A0(d_d8[44]), .B0(n5796), .C0(n5797[8]), .D0(d8[44]), 
          .A1(d_d8[45]), .B1(n5796), .C1(n5797[9]), .D1(d8[45]), .CIN(n11848), 
          .COUT(n11849), .S0(d9_71__N_1675[44]), .S1(d9_71__N_1675[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1095_11.INIT0 = 16'hb874;
    defparam add_1095_11.INIT1 = 16'hb874;
    defparam add_1095_11.INJECT1_0 = "NO";
    defparam add_1095_11.INJECT1_1 = "NO";
    CCU2D add_1095_9 (.A0(d_d8[42]), .B0(n5796), .C0(n5797[6]), .D0(d8[42]), 
          .A1(d_d8[43]), .B1(n5796), .C1(n5797[7]), .D1(d8[43]), .CIN(n11847), 
          .COUT(n11848), .S0(d9_71__N_1675[42]), .S1(d9_71__N_1675[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1095_9.INIT0 = 16'hb874;
    defparam add_1095_9.INIT1 = 16'hb874;
    defparam add_1095_9.INJECT1_0 = "NO";
    defparam add_1095_9.INJECT1_1 = "NO";
    CCU2D add_1095_7 (.A0(d_d8[40]), .B0(n5796), .C0(n5797[4]), .D0(d8[40]), 
          .A1(d_d8[41]), .B1(n5796), .C1(n5797[5]), .D1(d8[41]), .CIN(n11846), 
          .COUT(n11847), .S0(d9_71__N_1675[40]), .S1(d9_71__N_1675[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1095_7.INIT0 = 16'hb874;
    defparam add_1095_7.INIT1 = 16'hb874;
    defparam add_1095_7.INJECT1_0 = "NO";
    defparam add_1095_7.INJECT1_1 = "NO";
    CCU2D add_1095_5 (.A0(d_d8[38]), .B0(n5796), .C0(n5797[2]), .D0(d8[38]), 
          .A1(d_d8[39]), .B1(n5796), .C1(n5797[3]), .D1(d8[39]), .CIN(n11845), 
          .COUT(n11846), .S0(d9_71__N_1675[38]), .S1(d9_71__N_1675[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1095_5.INIT0 = 16'hb874;
    defparam add_1095_5.INIT1 = 16'hb874;
    defparam add_1095_5.INJECT1_0 = "NO";
    defparam add_1095_5.INJECT1_1 = "NO";
    CCU2D add_1100_13 (.A0(d9[47]), .B0(d_d9[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[48]), .B1(d_d9[48]), .C1(GND_net), .D1(GND_net), .CIN(n11810), 
          .COUT(n11811));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1100_13.INIT0 = 16'h5999;
    defparam add_1100_13.INIT1 = 16'h5999;
    defparam add_1100_13.INJECT1_0 = "NO";
    defparam add_1100_13.INJECT1_1 = "NO";
    CCU2D add_1100_11 (.A0(d9[45]), .B0(d_d9[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[46]), .B1(d_d9[46]), .C1(GND_net), .D1(GND_net), .CIN(n11809), 
          .COUT(n11810));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1100_11.INIT0 = 16'h5999;
    defparam add_1100_11.INIT1 = 16'h5999;
    defparam add_1100_11.INJECT1_0 = "NO";
    defparam add_1100_11.INJECT1_1 = "NO";
    LUT4 mux_1237_i11_3_lut (.A(n5949[30]), .B(n5987[30]), .C(n5948), 
         .Z(d10_71__N_1747[66])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1237_i11_3_lut.init = 16'hcaca;
    CCU2D add_1100_9 (.A0(d9[43]), .B0(d_d9[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[44]), .B1(d_d9[44]), .C1(GND_net), .D1(GND_net), .CIN(n11808), 
          .COUT(n11809));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1100_9.INIT0 = 16'h5999;
    defparam add_1100_9.INIT1 = 16'h5999;
    defparam add_1100_9.INJECT1_0 = "NO";
    defparam add_1100_9.INJECT1_1 = "NO";
    LUT4 mux_1237_i12_3_lut (.A(n5949[31]), .B(n5987[31]), .C(n5948), 
         .Z(d10_71__N_1747[67])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1237_i12_3_lut.init = 16'hcaca;
    CCU2D add_1100_7 (.A0(d9[41]), .B0(d_d9[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[42]), .B1(d_d9[42]), .C1(GND_net), .D1(GND_net), .CIN(n11807), 
          .COUT(n11808));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1100_7.INIT0 = 16'h5999;
    defparam add_1100_7.INIT1 = 16'h5999;
    defparam add_1100_7.INJECT1_0 = "NO";
    defparam add_1100_7.INJECT1_1 = "NO";
    CCU2D add_1100_5 (.A0(d9[39]), .B0(d_d9[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[40]), .B1(d_d9[40]), .C1(GND_net), .D1(GND_net), .CIN(n11806), 
          .COUT(n11807));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1100_5.INIT0 = 16'h5999;
    defparam add_1100_5.INIT1 = 16'h5999;
    defparam add_1100_5.INJECT1_0 = "NO";
    defparam add_1100_5.INJECT1_1 = "NO";
    FD1S3AX v_comb_66_rep_85 (.D(osc_clk_enable_1458), .CK(osc_clk), .Q(osc_clk_enable_247)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_85.GSR = "ENABLED";
    LUT4 mux_1237_i13_3_lut (.A(n5949[32]), .B(n5987[32]), .C(n5948), 
         .Z(d10_71__N_1747[68])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1237_i13_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i137_3_lut_4_lut_adj_36 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n13488), .D(d10[65]), .Z(n137)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i137_3_lut_4_lut_adj_36.init = 16'hf960;
    FD1P3AX d_d_tmp_i0_i37 (.D(d_tmp[37]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i38 (.D(d_tmp[38]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i38.GSR = "ENABLED";
    CCU2D add_1049_36 (.A0(d1[70]), .B0(d2[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[71]), .B1(d2[71]), .C1(GND_net), .D1(GND_net), .CIN(n12248), 
          .S0(n4429[34]), .S1(n4429[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1049_36.INIT0 = 16'h5666;
    defparam add_1049_36.INIT1 = 16'h5666;
    defparam add_1049_36.INJECT1_0 = "NO";
    defparam add_1049_36.INJECT1_1 = "NO";
    LUT4 mux_1237_i14_3_lut (.A(n5949[33]), .B(n5987[33]), .C(n5948), 
         .Z(d10_71__N_1747[69])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1237_i14_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i66_3_lut (.A(d10[65]), .B(d10[66]), .C(\CICGain[0] ), 
         .Z(n66_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i66_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i133_3_lut_4_lut_adj_37 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63_c), .D(d10[61]), .Z(n133)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i133_3_lut_4_lut_adj_37.init = 16'hf960;
    CCU2D add_1100_3 (.A0(d9[37]), .B0(d_d9[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[38]), .B1(d_d9[38]), .C1(GND_net), .D1(GND_net), .CIN(n11805), 
          .COUT(n11806));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1100_3.INIT0 = 16'h5999;
    defparam add_1100_3.INIT1 = 16'h5999;
    defparam add_1100_3.INJECT1_0 = "NO";
    defparam add_1100_3.INJECT1_1 = "NO";
    CCU2D add_1100_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d9[36]), .B1(d_d9[36]), .C1(GND_net), .D1(GND_net), .COUT(n11805));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1100_1.INIT0 = 16'h0000;
    defparam add_1100_1.INIT1 = 16'h5999;
    defparam add_1100_1.INJECT1_0 = "NO";
    defparam add_1100_1.INJECT1_1 = "NO";
    LUT4 shift_right_31_i61_3_lut (.A(d10[60]), .B(d10[61]), .C(\CICGain[0] ), 
         .Z(n61_adj_2521)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i61_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i136_3_lut_4_lut_adj_38 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66_c), .D(d10[64]), .Z(n136)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i136_3_lut_4_lut_adj_38.init = 16'hf960;
    LUT4 shift_right_31_i132_3_lut_4_lut_adj_39 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n62_c), .D(d10[60]), .Z(n132)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i132_3_lut_4_lut_adj_39.init = 16'hf960;
    FD1P3AX d_tmp_i0_i21 (.D(d5[21]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i25 (.D(d_tmp[25]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i24 (.D(d_tmp[24]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i23 (.D(d_tmp[23]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i22 (.D(d_tmp[22]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i22.GSR = "ENABLED";
    CCU2D add_1099_31 (.A0(d9[65]), .B0(d_d9[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[66]), .B1(d_d9[66]), .C1(GND_net), .D1(GND_net), .CIN(n11837), 
          .COUT(n11838), .S0(n5949[29]), .S1(n5949[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1099_31.INIT0 = 16'h5999;
    defparam add_1099_31.INIT1 = 16'h5999;
    defparam add_1099_31.INJECT1_0 = "NO";
    defparam add_1099_31.INJECT1_1 = "NO";
    FD1P3AX d_d_tmp_i0_i21 (.D(d_tmp[21]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i20 (.D(d_tmp[20]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i19 (.D(d_tmp[19]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i18 (.D(d_tmp[18]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i17 (.D(d_tmp[17]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i16 (.D(d_tmp[16]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i15 (.D(d_tmp[15]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i14 (.D(d_tmp[14]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i13 (.D(d_tmp[13]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i12 (.D(d_tmp[12]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i11 (.D(d_tmp[11]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i11.GSR = "ENABLED";
    CCU2D add_1099_29 (.A0(d9[63]), .B0(d_d9[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[64]), .B1(d_d9[64]), .C1(GND_net), .D1(GND_net), .CIN(n11836), 
          .COUT(n11837), .S0(n5949[27]), .S1(n5949[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1099_29.INIT0 = 16'h5999;
    defparam add_1099_29.INIT1 = 16'h5999;
    defparam add_1099_29.INJECT1_0 = "NO";
    defparam add_1099_29.INJECT1_1 = "NO";
    LUT4 mux_1237_i15_3_lut (.A(n5949[34]), .B(n5987[34]), .C(n5948), 
         .Z(d10_71__N_1747[70])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1237_i15_3_lut.init = 16'hcaca;
    FD1S3IX count__i1 (.D(n375[1]), .CK(osc_clk), .CD(n8376), .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i1.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i10 (.D(d_tmp[10]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i9 (.D(d_tmp[9]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i8 (.D(d_tmp[8]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i7 (.D(d_tmp[7]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i6 (.D(d_tmp[6]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i6.GSR = "ENABLED";
    LUT4 shift_right_31_i135_3_lut_4_lut_adj_40 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65_c), .D(d10[63]), .Z(n135)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i135_3_lut_4_lut_adj_40.init = 16'hf960;
    LUT4 mux_1237_i16_3_lut (.A(n5949[35]), .B(n5987[35]), .C(n5948), 
         .Z(d10_71__N_1747[71])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1237_i16_3_lut.init = 16'hcaca;
    FD1P3AX d_d_tmp_i0_i5 (.D(d_tmp[5]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i4 (.D(d_tmp[4]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i3 (.D(d_tmp[3]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i2 (.D(d_tmp[2]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i1 (.D(d_tmp[1]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d_d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i71 (.D(d5[71]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i70 (.D(d5[70]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i69 (.D(d5[69]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i68 (.D(d5[68]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i67 (.D(d5[67]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i66 (.D(d5[66]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i65 (.D(d5[65]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i64 (.D(d5[64]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i63 (.D(d5[63]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i62 (.D(d5[62]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i61 (.D(d5[61]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i60 (.D(d5[60]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i59 (.D(d5[59]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i58 (.D(d5[58]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i57 (.D(d5[57]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i56 (.D(d5[56]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i55 (.D(d5[55]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i54 (.D(d5[54]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i53 (.D(d5[53]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i52 (.D(d5[52]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i51 (.D(d5[51]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i50 (.D(d5[50]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i49 (.D(d5[49]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i48 (.D(d5[48]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i47 (.D(d5[47]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i46 (.D(d5[46]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i45 (.D(d5[45]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i44 (.D(d5[44]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i43 (.D(d5[43]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i42 (.D(d5[42]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i41 (.D(d5[41]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i40 (.D(d5[40]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i39 (.D(d5[39]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i38 (.D(d5[38]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i37 (.D(d5[37]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i36 (.D(d5[36]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i35 (.D(d5[35]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i34 (.D(d5[34]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i33 (.D(d5[33]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i32 (.D(d5[32]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i31 (.D(d5[31]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i30 (.D(d5[30]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i29 (.D(d5[29]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i28 (.D(d5[28]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i27 (.D(d5[27]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i26 (.D(d5[26]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i25 (.D(d5[25]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i24 (.D(d5[24]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i20 (.D(d5[20]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i19 (.D(d5[19]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i23 (.D(d5[23]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i23.GSR = "ENABLED";
    LUT4 i5704_4_lut_rep_95 (.A(n13125), .B(n13), .C(n13127), .D(n13113), 
         .Z(n13505)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i5704_4_lut_rep_95.init = 16'h2000;
    FD1P3AX d_tmp_i0_i18 (.D(d5[18]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i18.GSR = "ENABLED";
    LUT4 i5704_4_lut_rep_96 (.A(n13125), .B(n13), .C(n13127), .D(n13113), 
         .Z(osc_clk_enable_1458)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i5704_4_lut_rep_96.init = 16'h2000;
    FD1P3AX d_tmp_i0_i17 (.D(d5[17]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i17.GSR = "ENABLED";
    LUT4 i5645_2_lut (.A(count[10]), .B(count[2]), .Z(n13113)) /* synthesis lut_function=(A (B)) */ ;
    defparam i5645_2_lut.init = 16'h8888;
    FD1P3AX d_tmp_i0_i16 (.D(d5[16]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i16.GSR = "ENABLED";
    LUT4 shift_right_31_i68_3_lut (.A(d10[67]), .B(d10[68]), .C(\CICGain[0] ), 
         .Z(n68_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i68_3_lut.init = 16'hcaca;
    FD1P3AX d_tmp_i0_i15 (.D(d5[15]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i14 (.D(d5[14]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i14.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_83 (.D(osc_clk_enable_1458), .CK(osc_clk), .Q(osc_clk_enable_147)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_83.GSR = "ENABLED";
    LUT4 i4904_2_lut (.A(MixerOutSin[0]), .B(d1[0]), .Z(d1_71__N_418[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4904_2_lut.init = 16'h6666;
    FD1P3AX d_tmp_i0_i13 (.D(d5[13]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i13.GSR = "ENABLED";
    LUT4 shift_right_31_i134_3_lut_4_lut_adj_41 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64_c), .D(d10[62]), .Z(n134)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i134_3_lut_4_lut_adj_41.init = 16'hf960;
    FD1P3AX d_tmp_i0_i12 (.D(d5[12]), .SP(d_clk_tmp_N_1831), .CK(osc_clk), 
            .Q(d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i12.GSR = "ENABLED";
    FD1S3AX d2_i1 (.D(d2_71__N_490[1]), .CK(osc_clk), .Q(d2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i1.GSR = "ENABLED";
    CCU2D add_1049_34 (.A0(d1[68]), .B0(d2[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[69]), .B1(d2[69]), .C1(GND_net), .D1(GND_net), .CIN(n12247), 
          .COUT(n12248), .S0(n4429[32]), .S1(n4429[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1049_34.INIT0 = 16'h5666;
    defparam add_1049_34.INIT1 = 16'h5666;
    defparam add_1049_34.INJECT1_0 = "NO";
    defparam add_1049_34.INJECT1_1 = "NO";
    CCU2D add_1049_32 (.A0(d1[66]), .B0(d2[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[67]), .B1(d2[67]), .C1(GND_net), .D1(GND_net), .CIN(n12246), 
          .COUT(n12247), .S0(n4429[30]), .S1(n4429[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1049_32.INIT0 = 16'h5666;
    defparam add_1049_32.INIT1 = 16'h5666;
    defparam add_1049_32.INJECT1_0 = "NO";
    defparam add_1049_32.INJECT1_1 = "NO";
    CCU2D add_1049_30 (.A0(d1[64]), .B0(d2[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[65]), .B1(d2[65]), .C1(GND_net), .D1(GND_net), .CIN(n12245), 
          .COUT(n12246), .S0(n4429[28]), .S1(n4429[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1049_30.INIT0 = 16'h5666;
    defparam add_1049_30.INIT1 = 16'h5666;
    defparam add_1049_30.INJECT1_0 = "NO";
    defparam add_1049_30.INJECT1_1 = "NO";
    CCU2D add_1049_28 (.A0(d1[62]), .B0(d2[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[63]), .B1(d2[63]), .C1(GND_net), .D1(GND_net), .CIN(n12244), 
          .COUT(n12245), .S0(n4429[26]), .S1(n4429[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1049_28.INIT0 = 16'h5666;
    defparam add_1049_28.INIT1 = 16'h5666;
    defparam add_1049_28.INJECT1_0 = "NO";
    defparam add_1049_28.INJECT1_1 = "NO";
    CCU2D add_1049_26 (.A0(d1[60]), .B0(d2[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[61]), .B1(d2[61]), .C1(GND_net), .D1(GND_net), .CIN(n12243), 
          .COUT(n12244), .S0(n4429[24]), .S1(n4429[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1049_26.INIT0 = 16'h5666;
    defparam add_1049_26.INIT1 = 16'h5666;
    defparam add_1049_26.INJECT1_0 = "NO";
    defparam add_1049_26.INJECT1_1 = "NO";
    CCU2D add_1049_24 (.A0(d1[58]), .B0(d2[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[59]), .B1(d2[59]), .C1(GND_net), .D1(GND_net), .CIN(n12242), 
          .COUT(n12243), .S0(n4429[22]), .S1(n4429[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1049_24.INIT0 = 16'h5666;
    defparam add_1049_24.INIT1 = 16'h5666;
    defparam add_1049_24.INJECT1_0 = "NO";
    defparam add_1049_24.INJECT1_1 = "NO";
    CCU2D add_1049_22 (.A0(d1[56]), .B0(d2[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[57]), .B1(d2[57]), .C1(GND_net), .D1(GND_net), .CIN(n12241), 
          .COUT(n12242), .S0(n4429[20]), .S1(n4429[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1049_22.INIT0 = 16'h5666;
    defparam add_1049_22.INIT1 = 16'h5666;
    defparam add_1049_22.INJECT1_0 = "NO";
    defparam add_1049_22.INJECT1_1 = "NO";
    CCU2D add_1049_20 (.A0(d1[54]), .B0(d2[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[55]), .B1(d2[55]), .C1(GND_net), .D1(GND_net), .CIN(n12240), 
          .COUT(n12241), .S0(n4429[18]), .S1(n4429[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1049_20.INIT0 = 16'h5666;
    defparam add_1049_20.INIT1 = 16'h5666;
    defparam add_1049_20.INJECT1_0 = "NO";
    defparam add_1049_20.INJECT1_1 = "NO";
    CCU2D add_1049_18 (.A0(d1[52]), .B0(d2[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[53]), .B1(d2[53]), .C1(GND_net), .D1(GND_net), .CIN(n12239), 
          .COUT(n12240), .S0(n4429[16]), .S1(n4429[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1049_18.INIT0 = 16'h5666;
    defparam add_1049_18.INIT1 = 16'h5666;
    defparam add_1049_18.INJECT1_0 = "NO";
    defparam add_1049_18.INJECT1_1 = "NO";
    CCU2D add_1049_16 (.A0(d1[50]), .B0(d2[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[51]), .B1(d2[51]), .C1(GND_net), .D1(GND_net), .CIN(n12238), 
          .COUT(n12239), .S0(n4429[14]), .S1(n4429[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1049_16.INIT0 = 16'h5666;
    defparam add_1049_16.INIT1 = 16'h5666;
    defparam add_1049_16.INJECT1_0 = "NO";
    defparam add_1049_16.INJECT1_1 = "NO";
    CCU2D add_1049_14 (.A0(d1[48]), .B0(d2[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[49]), .B1(d2[49]), .C1(GND_net), .D1(GND_net), .CIN(n12237), 
          .COUT(n12238), .S0(n4429[12]), .S1(n4429[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1049_14.INIT0 = 16'h5666;
    defparam add_1049_14.INIT1 = 16'h5666;
    defparam add_1049_14.INJECT1_0 = "NO";
    defparam add_1049_14.INJECT1_1 = "NO";
    CCU2D add_1049_12 (.A0(d1[46]), .B0(d2[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[47]), .B1(d2[47]), .C1(GND_net), .D1(GND_net), .CIN(n12236), 
          .COUT(n12237), .S0(n4429[10]), .S1(n4429[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1049_12.INIT0 = 16'h5666;
    defparam add_1049_12.INIT1 = 16'h5666;
    defparam add_1049_12.INJECT1_0 = "NO";
    defparam add_1049_12.INJECT1_1 = "NO";
    CCU2D add_1049_10 (.A0(d1[44]), .B0(d2[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[45]), .B1(d2[45]), .C1(GND_net), .D1(GND_net), .CIN(n12235), 
          .COUT(n12236), .S0(n4429[8]), .S1(n4429[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1049_10.INIT0 = 16'h5666;
    defparam add_1049_10.INIT1 = 16'h5666;
    defparam add_1049_10.INJECT1_0 = "NO";
    defparam add_1049_10.INJECT1_1 = "NO";
    CCU2D add_1049_8 (.A0(d1[42]), .B0(d2[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[43]), .B1(d2[43]), .C1(GND_net), .D1(GND_net), .CIN(n12234), 
          .COUT(n12235), .S0(n4429[6]), .S1(n4429[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1049_8.INIT0 = 16'h5666;
    defparam add_1049_8.INIT1 = 16'h5666;
    defparam add_1049_8.INJECT1_0 = "NO";
    defparam add_1049_8.INJECT1_1 = "NO";
    FD1S3AX d2_i2 (.D(d2_71__N_490[2]), .CK(osc_clk), .Q(d2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i2.GSR = "ENABLED";
    FD1S3AX d2_i3 (.D(d2_71__N_490[3]), .CK(osc_clk), .Q(d2[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i3.GSR = "ENABLED";
    FD1S3AX d2_i4 (.D(d2_71__N_490[4]), .CK(osc_clk), .Q(d2[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i4.GSR = "ENABLED";
    FD1S3AX d2_i5 (.D(d2_71__N_490[5]), .CK(osc_clk), .Q(d2[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i5.GSR = "ENABLED";
    FD1S3AX d2_i6 (.D(d2_71__N_490[6]), .CK(osc_clk), .Q(d2[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i6.GSR = "ENABLED";
    FD1S3AX d2_i7 (.D(d2_71__N_490[7]), .CK(osc_clk), .Q(d2[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i7.GSR = "ENABLED";
    FD1S3AX d2_i8 (.D(d2_71__N_490[8]), .CK(osc_clk), .Q(d2[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i8.GSR = "ENABLED";
    FD1S3AX d2_i9 (.D(d2_71__N_490[9]), .CK(osc_clk), .Q(d2[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i9.GSR = "ENABLED";
    FD1S3AX d2_i10 (.D(d2_71__N_490[10]), .CK(osc_clk), .Q(d2[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i10.GSR = "ENABLED";
    FD1S3AX d2_i11 (.D(d2_71__N_490[11]), .CK(osc_clk), .Q(d2[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i11.GSR = "ENABLED";
    FD1S3AX d2_i12 (.D(d2_71__N_490[12]), .CK(osc_clk), .Q(d2[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i12.GSR = "ENABLED";
    FD1S3AX d2_i13 (.D(d2_71__N_490[13]), .CK(osc_clk), .Q(d2[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i13.GSR = "ENABLED";
    FD1S3AX d2_i14 (.D(d2_71__N_490[14]), .CK(osc_clk), .Q(d2[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i14.GSR = "ENABLED";
    FD1S3AX d2_i15 (.D(d2_71__N_490[15]), .CK(osc_clk), .Q(d2[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i15.GSR = "ENABLED";
    FD1S3AX d2_i16 (.D(d2_71__N_490[16]), .CK(osc_clk), .Q(d2[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i16.GSR = "ENABLED";
    FD1S3AX d2_i17 (.D(d2_71__N_490[17]), .CK(osc_clk), .Q(d2[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i17.GSR = "ENABLED";
    FD1S3AX d2_i18 (.D(d2_71__N_490[18]), .CK(osc_clk), .Q(d2[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i18.GSR = "ENABLED";
    FD1S3AX d2_i19 (.D(d2_71__N_490[19]), .CK(osc_clk), .Q(d2[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i19.GSR = "ENABLED";
    FD1S3AX d2_i20 (.D(d2_71__N_490[20]), .CK(osc_clk), .Q(d2[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i20.GSR = "ENABLED";
    FD1S3AX d2_i21 (.D(d2_71__N_490[21]), .CK(osc_clk), .Q(d2[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i21.GSR = "ENABLED";
    FD1S3AX d2_i22 (.D(d2_71__N_490[22]), .CK(osc_clk), .Q(d2[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i22.GSR = "ENABLED";
    FD1S3AX d2_i23 (.D(d2_71__N_490[23]), .CK(osc_clk), .Q(d2[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i23.GSR = "ENABLED";
    FD1S3AX d2_i24 (.D(d2_71__N_490[24]), .CK(osc_clk), .Q(d2[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i24.GSR = "ENABLED";
    FD1S3AX d2_i25 (.D(d2_71__N_490[25]), .CK(osc_clk), .Q(d2[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i25.GSR = "ENABLED";
    FD1S3AX d2_i26 (.D(d2_71__N_490[26]), .CK(osc_clk), .Q(d2[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i26.GSR = "ENABLED";
    FD1S3AX d2_i27 (.D(d2_71__N_490[27]), .CK(osc_clk), .Q(d2[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i27.GSR = "ENABLED";
    FD1S3AX d2_i28 (.D(d2_71__N_490[28]), .CK(osc_clk), .Q(d2[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i28.GSR = "ENABLED";
    FD1S3AX d2_i29 (.D(d2_71__N_490[29]), .CK(osc_clk), .Q(d2[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i29.GSR = "ENABLED";
    FD1S3AX d2_i30 (.D(d2_71__N_490[30]), .CK(osc_clk), .Q(d2[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i30.GSR = "ENABLED";
    FD1S3AX d2_i31 (.D(d2_71__N_490[31]), .CK(osc_clk), .Q(d2[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i31.GSR = "ENABLED";
    FD1S3AX d2_i32 (.D(d2_71__N_490[32]), .CK(osc_clk), .Q(d2[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i32.GSR = "ENABLED";
    FD1S3AX d2_i33 (.D(d2_71__N_490[33]), .CK(osc_clk), .Q(d2[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i33.GSR = "ENABLED";
    FD1S3AX d2_i34 (.D(d2_71__N_490[34]), .CK(osc_clk), .Q(d2[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i34.GSR = "ENABLED";
    FD1S3AX d2_i35 (.D(d2_71__N_490[35]), .CK(osc_clk), .Q(d2[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i35.GSR = "ENABLED";
    FD1S3AX d2_i36 (.D(d2_71__N_490[36]), .CK(osc_clk), .Q(d2[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i36.GSR = "ENABLED";
    FD1S3AX d2_i37 (.D(d2_71__N_490[37]), .CK(osc_clk), .Q(d2[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i37.GSR = "ENABLED";
    FD1S3AX d2_i38 (.D(d2_71__N_490[38]), .CK(osc_clk), .Q(d2[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i38.GSR = "ENABLED";
    FD1S3AX d2_i39 (.D(d2_71__N_490[39]), .CK(osc_clk), .Q(d2[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i39.GSR = "ENABLED";
    FD1S3AX d2_i40 (.D(d2_71__N_490[40]), .CK(osc_clk), .Q(d2[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i40.GSR = "ENABLED";
    FD1S3AX d2_i41 (.D(d2_71__N_490[41]), .CK(osc_clk), .Q(d2[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i41.GSR = "ENABLED";
    FD1S3AX d2_i42 (.D(d2_71__N_490[42]), .CK(osc_clk), .Q(d2[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i42.GSR = "ENABLED";
    FD1S3AX d2_i43 (.D(d2_71__N_490[43]), .CK(osc_clk), .Q(d2[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i43.GSR = "ENABLED";
    FD1S3AX d2_i44 (.D(d2_71__N_490[44]), .CK(osc_clk), .Q(d2[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i44.GSR = "ENABLED";
    FD1S3AX d2_i45 (.D(d2_71__N_490[45]), .CK(osc_clk), .Q(d2[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i45.GSR = "ENABLED";
    FD1S3AX d2_i46 (.D(d2_71__N_490[46]), .CK(osc_clk), .Q(d2[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i46.GSR = "ENABLED";
    FD1S3AX d2_i47 (.D(d2_71__N_490[47]), .CK(osc_clk), .Q(d2[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i47.GSR = "ENABLED";
    FD1S3AX d2_i48 (.D(d2_71__N_490[48]), .CK(osc_clk), .Q(d2[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i48.GSR = "ENABLED";
    FD1S3AX d2_i49 (.D(d2_71__N_490[49]), .CK(osc_clk), .Q(d2[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i49.GSR = "ENABLED";
    FD1S3AX d2_i50 (.D(d2_71__N_490[50]), .CK(osc_clk), .Q(d2[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i50.GSR = "ENABLED";
    FD1S3AX d2_i51 (.D(d2_71__N_490[51]), .CK(osc_clk), .Q(d2[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i51.GSR = "ENABLED";
    FD1S3AX d2_i52 (.D(d2_71__N_490[52]), .CK(osc_clk), .Q(d2[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i52.GSR = "ENABLED";
    FD1S3AX d2_i53 (.D(d2_71__N_490[53]), .CK(osc_clk), .Q(d2[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i53.GSR = "ENABLED";
    FD1S3AX d2_i54 (.D(d2_71__N_490[54]), .CK(osc_clk), .Q(d2[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i54.GSR = "ENABLED";
    FD1S3AX d2_i55 (.D(d2_71__N_490[55]), .CK(osc_clk), .Q(d2[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i55.GSR = "ENABLED";
    FD1S3AX d2_i56 (.D(d2_71__N_490[56]), .CK(osc_clk), .Q(d2[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i56.GSR = "ENABLED";
    FD1S3AX d2_i57 (.D(d2_71__N_490[57]), .CK(osc_clk), .Q(d2[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i57.GSR = "ENABLED";
    FD1S3AX d2_i58 (.D(d2_71__N_490[58]), .CK(osc_clk), .Q(d2[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i58.GSR = "ENABLED";
    FD1S3AX d2_i59 (.D(d2_71__N_490[59]), .CK(osc_clk), .Q(d2[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i59.GSR = "ENABLED";
    FD1S3AX d2_i60 (.D(d2_71__N_490[60]), .CK(osc_clk), .Q(d2[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i60.GSR = "ENABLED";
    FD1S3AX d2_i61 (.D(d2_71__N_490[61]), .CK(osc_clk), .Q(d2[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i61.GSR = "ENABLED";
    FD1S3AX d2_i62 (.D(d2_71__N_490[62]), .CK(osc_clk), .Q(d2[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i62.GSR = "ENABLED";
    FD1S3AX d2_i63 (.D(d2_71__N_490[63]), .CK(osc_clk), .Q(d2[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i63.GSR = "ENABLED";
    FD1S3AX d2_i64 (.D(d2_71__N_490[64]), .CK(osc_clk), .Q(d2[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i64.GSR = "ENABLED";
    FD1S3AX d2_i65 (.D(d2_71__N_490[65]), .CK(osc_clk), .Q(d2[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i65.GSR = "ENABLED";
    FD1S3AX d2_i66 (.D(d2_71__N_490[66]), .CK(osc_clk), .Q(d2[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i66.GSR = "ENABLED";
    FD1S3AX d2_i67 (.D(d2_71__N_490[67]), .CK(osc_clk), .Q(d2[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i67.GSR = "ENABLED";
    FD1S3AX d2_i68 (.D(d2_71__N_490[68]), .CK(osc_clk), .Q(d2[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i68.GSR = "ENABLED";
    FD1S3AX d2_i69 (.D(d2_71__N_490[69]), .CK(osc_clk), .Q(d2[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i69.GSR = "ENABLED";
    FD1S3AX d2_i70 (.D(d2_71__N_490[70]), .CK(osc_clk), .Q(d2[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i70.GSR = "ENABLED";
    FD1S3AX d2_i71 (.D(d2_71__N_490[71]), .CK(osc_clk), .Q(d2[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i71.GSR = "ENABLED";
    FD1S3AX d3_i1 (.D(d3_71__N_562[1]), .CK(osc_clk), .Q(d3[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i1.GSR = "ENABLED";
    FD1S3AX d3_i2 (.D(d3_71__N_562[2]), .CK(osc_clk), .Q(d3[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i2.GSR = "ENABLED";
    FD1S3AX d3_i3 (.D(d3_71__N_562[3]), .CK(osc_clk), .Q(d3[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i3.GSR = "ENABLED";
    FD1S3AX d3_i4 (.D(d3_71__N_562[4]), .CK(osc_clk), .Q(d3[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i4.GSR = "ENABLED";
    FD1S3AX d3_i5 (.D(d3_71__N_562[5]), .CK(osc_clk), .Q(d3[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i5.GSR = "ENABLED";
    FD1S3AX d3_i6 (.D(d3_71__N_562[6]), .CK(osc_clk), .Q(d3[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i6.GSR = "ENABLED";
    FD1S3AX d3_i7 (.D(d3_71__N_562[7]), .CK(osc_clk), .Q(d3[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i7.GSR = "ENABLED";
    FD1S3AX d3_i8 (.D(d3_71__N_562[8]), .CK(osc_clk), .Q(d3[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i8.GSR = "ENABLED";
    FD1S3AX d3_i9 (.D(d3_71__N_562[9]), .CK(osc_clk), .Q(d3[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i9.GSR = "ENABLED";
    FD1S3AX d3_i10 (.D(d3_71__N_562[10]), .CK(osc_clk), .Q(d3[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i10.GSR = "ENABLED";
    FD1S3AX d3_i11 (.D(d3_71__N_562[11]), .CK(osc_clk), .Q(d3[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i11.GSR = "ENABLED";
    FD1S3AX d3_i12 (.D(d3_71__N_562[12]), .CK(osc_clk), .Q(d3[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i12.GSR = "ENABLED";
    FD1S3AX d3_i13 (.D(d3_71__N_562[13]), .CK(osc_clk), .Q(d3[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i13.GSR = "ENABLED";
    FD1S3AX d3_i14 (.D(d3_71__N_562[14]), .CK(osc_clk), .Q(d3[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i14.GSR = "ENABLED";
    FD1S3AX d3_i15 (.D(d3_71__N_562[15]), .CK(osc_clk), .Q(d3[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i15.GSR = "ENABLED";
    FD1S3AX d3_i16 (.D(d3_71__N_562[16]), .CK(osc_clk), .Q(d3[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i16.GSR = "ENABLED";
    FD1S3AX d3_i17 (.D(d3_71__N_562[17]), .CK(osc_clk), .Q(d3[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i17.GSR = "ENABLED";
    FD1S3AX d3_i18 (.D(d3_71__N_562[18]), .CK(osc_clk), .Q(d3[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i18.GSR = "ENABLED";
    FD1S3AX d3_i19 (.D(d3_71__N_562[19]), .CK(osc_clk), .Q(d3[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i19.GSR = "ENABLED";
    FD1S3AX d3_i20 (.D(d3_71__N_562[20]), .CK(osc_clk), .Q(d3[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i20.GSR = "ENABLED";
    FD1S3AX d3_i21 (.D(d3_71__N_562[21]), .CK(osc_clk), .Q(d3[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i21.GSR = "ENABLED";
    FD1S3AX d3_i22 (.D(d3_71__N_562[22]), .CK(osc_clk), .Q(d3[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i22.GSR = "ENABLED";
    FD1S3AX d3_i23 (.D(d3_71__N_562[23]), .CK(osc_clk), .Q(d3[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i23.GSR = "ENABLED";
    FD1S3AX d3_i24 (.D(d3_71__N_562[24]), .CK(osc_clk), .Q(d3[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i24.GSR = "ENABLED";
    FD1S3AX d3_i25 (.D(d3_71__N_562[25]), .CK(osc_clk), .Q(d3[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i25.GSR = "ENABLED";
    FD1S3AX d3_i26 (.D(d3_71__N_562[26]), .CK(osc_clk), .Q(d3[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i26.GSR = "ENABLED";
    FD1S3AX d3_i27 (.D(d3_71__N_562[27]), .CK(osc_clk), .Q(d3[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i27.GSR = "ENABLED";
    FD1S3AX d3_i28 (.D(d3_71__N_562[28]), .CK(osc_clk), .Q(d3[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i28.GSR = "ENABLED";
    FD1S3AX d3_i29 (.D(d3_71__N_562[29]), .CK(osc_clk), .Q(d3[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i29.GSR = "ENABLED";
    FD1S3AX d3_i30 (.D(d3_71__N_562[30]), .CK(osc_clk), .Q(d3[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i30.GSR = "ENABLED";
    FD1S3AX d3_i31 (.D(d3_71__N_562[31]), .CK(osc_clk), .Q(d3[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i31.GSR = "ENABLED";
    FD1S3AX d3_i32 (.D(d3_71__N_562[32]), .CK(osc_clk), .Q(d3[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i32.GSR = "ENABLED";
    FD1S3AX d3_i33 (.D(d3_71__N_562[33]), .CK(osc_clk), .Q(d3[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i33.GSR = "ENABLED";
    FD1S3AX d3_i34 (.D(d3_71__N_562[34]), .CK(osc_clk), .Q(d3[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i34.GSR = "ENABLED";
    FD1S3AX d3_i35 (.D(d3_71__N_562[35]), .CK(osc_clk), .Q(d3[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i35.GSR = "ENABLED";
    FD1S3AX d3_i36 (.D(d3_71__N_562[36]), .CK(osc_clk), .Q(d3[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i36.GSR = "ENABLED";
    FD1S3AX d3_i37 (.D(d3_71__N_562[37]), .CK(osc_clk), .Q(d3[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i37.GSR = "ENABLED";
    FD1S3AX d3_i38 (.D(d3_71__N_562[38]), .CK(osc_clk), .Q(d3[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i38.GSR = "ENABLED";
    FD1S3AX d3_i39 (.D(d3_71__N_562[39]), .CK(osc_clk), .Q(d3[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i39.GSR = "ENABLED";
    FD1S3AX d3_i40 (.D(d3_71__N_562[40]), .CK(osc_clk), .Q(d3[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i40.GSR = "ENABLED";
    FD1S3AX d3_i41 (.D(d3_71__N_562[41]), .CK(osc_clk), .Q(d3[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i41.GSR = "ENABLED";
    FD1S3AX d3_i42 (.D(d3_71__N_562[42]), .CK(osc_clk), .Q(d3[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i42.GSR = "ENABLED";
    FD1S3AX d3_i43 (.D(d3_71__N_562[43]), .CK(osc_clk), .Q(d3[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i43.GSR = "ENABLED";
    FD1S3AX d3_i44 (.D(d3_71__N_562[44]), .CK(osc_clk), .Q(d3[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i44.GSR = "ENABLED";
    FD1S3AX d3_i45 (.D(d3_71__N_562[45]), .CK(osc_clk), .Q(d3[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i45.GSR = "ENABLED";
    FD1S3AX d3_i46 (.D(d3_71__N_562[46]), .CK(osc_clk), .Q(d3[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i46.GSR = "ENABLED";
    FD1S3AX d3_i47 (.D(d3_71__N_562[47]), .CK(osc_clk), .Q(d3[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i47.GSR = "ENABLED";
    FD1S3AX d3_i48 (.D(d3_71__N_562[48]), .CK(osc_clk), .Q(d3[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i48.GSR = "ENABLED";
    FD1S3AX d3_i49 (.D(d3_71__N_562[49]), .CK(osc_clk), .Q(d3[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i49.GSR = "ENABLED";
    FD1S3AX d3_i50 (.D(d3_71__N_562[50]), .CK(osc_clk), .Q(d3[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i50.GSR = "ENABLED";
    FD1S3AX d3_i51 (.D(d3_71__N_562[51]), .CK(osc_clk), .Q(d3[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i51.GSR = "ENABLED";
    FD1S3AX d3_i52 (.D(d3_71__N_562[52]), .CK(osc_clk), .Q(d3[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i52.GSR = "ENABLED";
    FD1S3AX d3_i53 (.D(d3_71__N_562[53]), .CK(osc_clk), .Q(d3[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i53.GSR = "ENABLED";
    FD1S3AX d3_i54 (.D(d3_71__N_562[54]), .CK(osc_clk), .Q(d3[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i54.GSR = "ENABLED";
    FD1S3AX d3_i55 (.D(d3_71__N_562[55]), .CK(osc_clk), .Q(d3[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i55.GSR = "ENABLED";
    FD1S3AX d3_i56 (.D(d3_71__N_562[56]), .CK(osc_clk), .Q(d3[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i56.GSR = "ENABLED";
    FD1S3AX d3_i57 (.D(d3_71__N_562[57]), .CK(osc_clk), .Q(d3[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i57.GSR = "ENABLED";
    FD1S3AX d3_i58 (.D(d3_71__N_562[58]), .CK(osc_clk), .Q(d3[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i58.GSR = "ENABLED";
    FD1S3AX d3_i59 (.D(d3_71__N_562[59]), .CK(osc_clk), .Q(d3[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i59.GSR = "ENABLED";
    FD1S3AX d3_i60 (.D(d3_71__N_562[60]), .CK(osc_clk), .Q(d3[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i60.GSR = "ENABLED";
    FD1S3AX d3_i61 (.D(d3_71__N_562[61]), .CK(osc_clk), .Q(d3[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i61.GSR = "ENABLED";
    FD1S3AX d3_i62 (.D(d3_71__N_562[62]), .CK(osc_clk), .Q(d3[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i62.GSR = "ENABLED";
    FD1S3AX d3_i63 (.D(d3_71__N_562[63]), .CK(osc_clk), .Q(d3[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i63.GSR = "ENABLED";
    FD1S3AX d3_i64 (.D(d3_71__N_562[64]), .CK(osc_clk), .Q(d3[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i64.GSR = "ENABLED";
    FD1S3AX d3_i65 (.D(d3_71__N_562[65]), .CK(osc_clk), .Q(d3[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i65.GSR = "ENABLED";
    FD1S3AX d3_i66 (.D(d3_71__N_562[66]), .CK(osc_clk), .Q(d3[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i66.GSR = "ENABLED";
    FD1S3AX d3_i67 (.D(d3_71__N_562[67]), .CK(osc_clk), .Q(d3[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i67.GSR = "ENABLED";
    FD1S3AX d3_i68 (.D(d3_71__N_562[68]), .CK(osc_clk), .Q(d3[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i68.GSR = "ENABLED";
    FD1S3AX d3_i69 (.D(d3_71__N_562[69]), .CK(osc_clk), .Q(d3[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i69.GSR = "ENABLED";
    FD1S3AX d3_i70 (.D(d3_71__N_562[70]), .CK(osc_clk), .Q(d3[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i70.GSR = "ENABLED";
    FD1S3AX d3_i71 (.D(d3_71__N_562[71]), .CK(osc_clk), .Q(d3[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i71.GSR = "ENABLED";
    FD1S3AX d4_i1 (.D(d4_71__N_634[1]), .CK(osc_clk), .Q(d4[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i1.GSR = "ENABLED";
    FD1S3AX d4_i2 (.D(d4_71__N_634[2]), .CK(osc_clk), .Q(d4[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i2.GSR = "ENABLED";
    FD1S3AX d4_i3 (.D(d4_71__N_634[3]), .CK(osc_clk), .Q(d4[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i3.GSR = "ENABLED";
    FD1S3AX d4_i4 (.D(d4_71__N_634[4]), .CK(osc_clk), .Q(d4[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i4.GSR = "ENABLED";
    FD1S3AX d4_i5 (.D(d4_71__N_634[5]), .CK(osc_clk), .Q(d4[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i5.GSR = "ENABLED";
    FD1S3AX d4_i6 (.D(d4_71__N_634[6]), .CK(osc_clk), .Q(d4[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i6.GSR = "ENABLED";
    FD1S3AX d4_i7 (.D(d4_71__N_634[7]), .CK(osc_clk), .Q(d4[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i7.GSR = "ENABLED";
    FD1S3AX d4_i8 (.D(d4_71__N_634[8]), .CK(osc_clk), .Q(d4[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i8.GSR = "ENABLED";
    FD1S3AX d4_i9 (.D(d4_71__N_634[9]), .CK(osc_clk), .Q(d4[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i9.GSR = "ENABLED";
    FD1S3AX d4_i10 (.D(d4_71__N_634[10]), .CK(osc_clk), .Q(d4[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i10.GSR = "ENABLED";
    FD1S3AX d4_i11 (.D(d4_71__N_634[11]), .CK(osc_clk), .Q(d4[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i11.GSR = "ENABLED";
    FD1S3AX d4_i12 (.D(d4_71__N_634[12]), .CK(osc_clk), .Q(d4[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i12.GSR = "ENABLED";
    FD1S3AX d4_i13 (.D(d4_71__N_634[13]), .CK(osc_clk), .Q(d4[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i13.GSR = "ENABLED";
    FD1S3AX d4_i14 (.D(d4_71__N_634[14]), .CK(osc_clk), .Q(d4[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i14.GSR = "ENABLED";
    FD1S3AX d4_i15 (.D(d4_71__N_634[15]), .CK(osc_clk), .Q(d4[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i15.GSR = "ENABLED";
    FD1S3AX d4_i16 (.D(d4_71__N_634[16]), .CK(osc_clk), .Q(d4[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i16.GSR = "ENABLED";
    FD1S3AX d4_i17 (.D(d4_71__N_634[17]), .CK(osc_clk), .Q(d4[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i17.GSR = "ENABLED";
    FD1S3AX d4_i18 (.D(d4_71__N_634[18]), .CK(osc_clk), .Q(d4[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i18.GSR = "ENABLED";
    FD1S3AX d4_i19 (.D(d4_71__N_634[19]), .CK(osc_clk), .Q(d4[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i19.GSR = "ENABLED";
    FD1S3AX d4_i20 (.D(d4_71__N_634[20]), .CK(osc_clk), .Q(d4[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i20.GSR = "ENABLED";
    FD1S3AX d4_i21 (.D(d4_71__N_634[21]), .CK(osc_clk), .Q(d4[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i21.GSR = "ENABLED";
    FD1S3AX d4_i22 (.D(d4_71__N_634[22]), .CK(osc_clk), .Q(d4[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i22.GSR = "ENABLED";
    FD1S3AX d4_i23 (.D(d4_71__N_634[23]), .CK(osc_clk), .Q(d4[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i23.GSR = "ENABLED";
    FD1S3AX d4_i24 (.D(d4_71__N_634[24]), .CK(osc_clk), .Q(d4[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i24.GSR = "ENABLED";
    FD1S3AX d4_i25 (.D(d4_71__N_634[25]), .CK(osc_clk), .Q(d4[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i25.GSR = "ENABLED";
    FD1S3AX d4_i26 (.D(d4_71__N_634[26]), .CK(osc_clk), .Q(d4[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i26.GSR = "ENABLED";
    FD1S3AX d4_i27 (.D(d4_71__N_634[27]), .CK(osc_clk), .Q(d4[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i27.GSR = "ENABLED";
    FD1S3AX d4_i28 (.D(d4_71__N_634[28]), .CK(osc_clk), .Q(d4[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i28.GSR = "ENABLED";
    FD1S3AX d4_i29 (.D(d4_71__N_634[29]), .CK(osc_clk), .Q(d4[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i29.GSR = "ENABLED";
    FD1S3AX d4_i30 (.D(d4_71__N_634[30]), .CK(osc_clk), .Q(d4[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i30.GSR = "ENABLED";
    FD1S3AX d4_i31 (.D(d4_71__N_634[31]), .CK(osc_clk), .Q(d4[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i31.GSR = "ENABLED";
    FD1S3AX d4_i32 (.D(d4_71__N_634[32]), .CK(osc_clk), .Q(d4[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i32.GSR = "ENABLED";
    FD1S3AX d4_i33 (.D(d4_71__N_634[33]), .CK(osc_clk), .Q(d4[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i33.GSR = "ENABLED";
    FD1S3AX d4_i34 (.D(d4_71__N_634[34]), .CK(osc_clk), .Q(d4[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i34.GSR = "ENABLED";
    FD1S3AX d4_i35 (.D(d4_71__N_634[35]), .CK(osc_clk), .Q(d4[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i35.GSR = "ENABLED";
    FD1S3AX d4_i36 (.D(d4_71__N_634[36]), .CK(osc_clk), .Q(d4[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i36.GSR = "ENABLED";
    FD1S3AX d4_i37 (.D(d4_71__N_634[37]), .CK(osc_clk), .Q(d4[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i37.GSR = "ENABLED";
    FD1S3AX d4_i38 (.D(d4_71__N_634[38]), .CK(osc_clk), .Q(d4[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i38.GSR = "ENABLED";
    FD1S3AX d4_i39 (.D(d4_71__N_634[39]), .CK(osc_clk), .Q(d4[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i39.GSR = "ENABLED";
    FD1S3AX d4_i40 (.D(d4_71__N_634[40]), .CK(osc_clk), .Q(d4[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i40.GSR = "ENABLED";
    FD1S3AX d4_i41 (.D(d4_71__N_634[41]), .CK(osc_clk), .Q(d4[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i41.GSR = "ENABLED";
    FD1S3AX d4_i42 (.D(d4_71__N_634[42]), .CK(osc_clk), .Q(d4[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i42.GSR = "ENABLED";
    FD1S3AX d4_i43 (.D(d4_71__N_634[43]), .CK(osc_clk), .Q(d4[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i43.GSR = "ENABLED";
    FD1S3AX d4_i44 (.D(d4_71__N_634[44]), .CK(osc_clk), .Q(d4[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i44.GSR = "ENABLED";
    FD1S3AX d4_i45 (.D(d4_71__N_634[45]), .CK(osc_clk), .Q(d4[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i45.GSR = "ENABLED";
    FD1S3AX d4_i46 (.D(d4_71__N_634[46]), .CK(osc_clk), .Q(d4[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i46.GSR = "ENABLED";
    FD1S3AX d4_i47 (.D(d4_71__N_634[47]), .CK(osc_clk), .Q(d4[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i47.GSR = "ENABLED";
    FD1S3AX d4_i48 (.D(d4_71__N_634[48]), .CK(osc_clk), .Q(d4[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i48.GSR = "ENABLED";
    FD1S3AX d4_i49 (.D(d4_71__N_634[49]), .CK(osc_clk), .Q(d4[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i49.GSR = "ENABLED";
    FD1S3AX d4_i50 (.D(d4_71__N_634[50]), .CK(osc_clk), .Q(d4[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i50.GSR = "ENABLED";
    FD1S3AX d4_i51 (.D(d4_71__N_634[51]), .CK(osc_clk), .Q(d4[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i51.GSR = "ENABLED";
    FD1S3AX d4_i52 (.D(d4_71__N_634[52]), .CK(osc_clk), .Q(d4[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i52.GSR = "ENABLED";
    FD1S3AX d4_i53 (.D(d4_71__N_634[53]), .CK(osc_clk), .Q(d4[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i53.GSR = "ENABLED";
    FD1S3AX d4_i54 (.D(d4_71__N_634[54]), .CK(osc_clk), .Q(d4[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i54.GSR = "ENABLED";
    FD1S3AX d4_i55 (.D(d4_71__N_634[55]), .CK(osc_clk), .Q(d4[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i55.GSR = "ENABLED";
    FD1S3AX d4_i56 (.D(d4_71__N_634[56]), .CK(osc_clk), .Q(d4[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i56.GSR = "ENABLED";
    FD1S3AX d4_i57 (.D(d4_71__N_634[57]), .CK(osc_clk), .Q(d4[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i57.GSR = "ENABLED";
    FD1S3AX d4_i58 (.D(d4_71__N_634[58]), .CK(osc_clk), .Q(d4[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i58.GSR = "ENABLED";
    FD1S3AX d4_i59 (.D(d4_71__N_634[59]), .CK(osc_clk), .Q(d4[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i59.GSR = "ENABLED";
    FD1S3AX d4_i60 (.D(d4_71__N_634[60]), .CK(osc_clk), .Q(d4[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i60.GSR = "ENABLED";
    FD1S3AX d4_i61 (.D(d4_71__N_634[61]), .CK(osc_clk), .Q(d4[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i61.GSR = "ENABLED";
    FD1S3AX d4_i62 (.D(d4_71__N_634[62]), .CK(osc_clk), .Q(d4[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i62.GSR = "ENABLED";
    FD1S3AX d4_i63 (.D(d4_71__N_634[63]), .CK(osc_clk), .Q(d4[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i63.GSR = "ENABLED";
    FD1S3AX d4_i64 (.D(d4_71__N_634[64]), .CK(osc_clk), .Q(d4[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i64.GSR = "ENABLED";
    FD1S3AX d4_i65 (.D(d4_71__N_634[65]), .CK(osc_clk), .Q(d4[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i65.GSR = "ENABLED";
    FD1S3AX d4_i66 (.D(d4_71__N_634[66]), .CK(osc_clk), .Q(d4[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i66.GSR = "ENABLED";
    FD1S3AX d4_i67 (.D(d4_71__N_634[67]), .CK(osc_clk), .Q(d4[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i67.GSR = "ENABLED";
    FD1S3AX d4_i68 (.D(d4_71__N_634[68]), .CK(osc_clk), .Q(d4[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i68.GSR = "ENABLED";
    FD1S3AX d4_i69 (.D(d4_71__N_634[69]), .CK(osc_clk), .Q(d4[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i69.GSR = "ENABLED";
    FD1S3AX d4_i70 (.D(d4_71__N_634[70]), .CK(osc_clk), .Q(d4[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i70.GSR = "ENABLED";
    FD1S3AX d4_i71 (.D(d4_71__N_634[71]), .CK(osc_clk), .Q(d4[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i71.GSR = "ENABLED";
    FD1S3AX d5_i1 (.D(d5_71__N_706[1]), .CK(osc_clk), .Q(d5[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i1.GSR = "ENABLED";
    FD1S3AX d5_i2 (.D(d5_71__N_706[2]), .CK(osc_clk), .Q(d5[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i2.GSR = "ENABLED";
    FD1S3AX d5_i3 (.D(d5_71__N_706[3]), .CK(osc_clk), .Q(d5[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i3.GSR = "ENABLED";
    FD1S3AX d5_i4 (.D(d5_71__N_706[4]), .CK(osc_clk), .Q(d5[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i4.GSR = "ENABLED";
    FD1S3AX d5_i5 (.D(d5_71__N_706[5]), .CK(osc_clk), .Q(d5[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i5.GSR = "ENABLED";
    FD1S3AX d5_i6 (.D(d5_71__N_706[6]), .CK(osc_clk), .Q(d5[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i6.GSR = "ENABLED";
    FD1S3AX d5_i7 (.D(d5_71__N_706[7]), .CK(osc_clk), .Q(d5[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i7.GSR = "ENABLED";
    FD1S3AX d5_i8 (.D(d5_71__N_706[8]), .CK(osc_clk), .Q(d5[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i8.GSR = "ENABLED";
    FD1S3AX d5_i9 (.D(d5_71__N_706[9]), .CK(osc_clk), .Q(d5[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i9.GSR = "ENABLED";
    FD1S3AX d5_i10 (.D(d5_71__N_706[10]), .CK(osc_clk), .Q(d5[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i10.GSR = "ENABLED";
    FD1S3AX d5_i11 (.D(d5_71__N_706[11]), .CK(osc_clk), .Q(d5[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i11.GSR = "ENABLED";
    FD1S3AX d5_i12 (.D(d5_71__N_706[12]), .CK(osc_clk), .Q(d5[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i12.GSR = "ENABLED";
    FD1S3AX d5_i13 (.D(d5_71__N_706[13]), .CK(osc_clk), .Q(d5[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i13.GSR = "ENABLED";
    FD1S3AX d5_i14 (.D(d5_71__N_706[14]), .CK(osc_clk), .Q(d5[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i14.GSR = "ENABLED";
    FD1S3AX d5_i15 (.D(d5_71__N_706[15]), .CK(osc_clk), .Q(d5[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i15.GSR = "ENABLED";
    FD1S3AX d5_i16 (.D(d5_71__N_706[16]), .CK(osc_clk), .Q(d5[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i16.GSR = "ENABLED";
    FD1S3AX d5_i17 (.D(d5_71__N_706[17]), .CK(osc_clk), .Q(d5[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i17.GSR = "ENABLED";
    FD1S3AX d5_i18 (.D(d5_71__N_706[18]), .CK(osc_clk), .Q(d5[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i18.GSR = "ENABLED";
    FD1S3AX d5_i19 (.D(d5_71__N_706[19]), .CK(osc_clk), .Q(d5[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i19.GSR = "ENABLED";
    FD1S3AX d5_i20 (.D(d5_71__N_706[20]), .CK(osc_clk), .Q(d5[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i20.GSR = "ENABLED";
    FD1S3AX d5_i21 (.D(d5_71__N_706[21]), .CK(osc_clk), .Q(d5[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i21.GSR = "ENABLED";
    FD1S3AX d5_i22 (.D(d5_71__N_706[22]), .CK(osc_clk), .Q(d5[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i22.GSR = "ENABLED";
    FD1S3AX d5_i23 (.D(d5_71__N_706[23]), .CK(osc_clk), .Q(d5[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i23.GSR = "ENABLED";
    FD1S3AX d5_i24 (.D(d5_71__N_706[24]), .CK(osc_clk), .Q(d5[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i24.GSR = "ENABLED";
    FD1S3AX d5_i25 (.D(d5_71__N_706[25]), .CK(osc_clk), .Q(d5[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i25.GSR = "ENABLED";
    FD1S3AX d5_i26 (.D(d5_71__N_706[26]), .CK(osc_clk), .Q(d5[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i26.GSR = "ENABLED";
    FD1S3AX d5_i27 (.D(d5_71__N_706[27]), .CK(osc_clk), .Q(d5[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i27.GSR = "ENABLED";
    FD1S3AX d5_i28 (.D(d5_71__N_706[28]), .CK(osc_clk), .Q(d5[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i28.GSR = "ENABLED";
    FD1S3AX d5_i29 (.D(d5_71__N_706[29]), .CK(osc_clk), .Q(d5[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i29.GSR = "ENABLED";
    FD1S3AX d5_i30 (.D(d5_71__N_706[30]), .CK(osc_clk), .Q(d5[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i30.GSR = "ENABLED";
    FD1S3AX d5_i31 (.D(d5_71__N_706[31]), .CK(osc_clk), .Q(d5[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i31.GSR = "ENABLED";
    FD1S3AX d5_i32 (.D(d5_71__N_706[32]), .CK(osc_clk), .Q(d5[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i32.GSR = "ENABLED";
    FD1S3AX d5_i33 (.D(d5_71__N_706[33]), .CK(osc_clk), .Q(d5[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i33.GSR = "ENABLED";
    FD1S3AX d5_i34 (.D(d5_71__N_706[34]), .CK(osc_clk), .Q(d5[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i34.GSR = "ENABLED";
    FD1S3AX d5_i35 (.D(d5_71__N_706[35]), .CK(osc_clk), .Q(d5[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i35.GSR = "ENABLED";
    FD1S3AX d5_i36 (.D(d5_71__N_706[36]), .CK(osc_clk), .Q(d5[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i36.GSR = "ENABLED";
    FD1S3AX d5_i37 (.D(d5_71__N_706[37]), .CK(osc_clk), .Q(d5[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i37.GSR = "ENABLED";
    FD1S3AX d5_i38 (.D(d5_71__N_706[38]), .CK(osc_clk), .Q(d5[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i38.GSR = "ENABLED";
    FD1S3AX d5_i39 (.D(d5_71__N_706[39]), .CK(osc_clk), .Q(d5[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i39.GSR = "ENABLED";
    FD1S3AX d5_i40 (.D(d5_71__N_706[40]), .CK(osc_clk), .Q(d5[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i40.GSR = "ENABLED";
    FD1S3AX d5_i41 (.D(d5_71__N_706[41]), .CK(osc_clk), .Q(d5[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i41.GSR = "ENABLED";
    FD1S3AX d5_i42 (.D(d5_71__N_706[42]), .CK(osc_clk), .Q(d5[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i42.GSR = "ENABLED";
    FD1S3AX d5_i43 (.D(d5_71__N_706[43]), .CK(osc_clk), .Q(d5[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i43.GSR = "ENABLED";
    FD1S3AX d5_i44 (.D(d5_71__N_706[44]), .CK(osc_clk), .Q(d5[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i44.GSR = "ENABLED";
    FD1S3AX d5_i45 (.D(d5_71__N_706[45]), .CK(osc_clk), .Q(d5[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i45.GSR = "ENABLED";
    FD1S3AX d5_i46 (.D(d5_71__N_706[46]), .CK(osc_clk), .Q(d5[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i46.GSR = "ENABLED";
    FD1S3AX d5_i47 (.D(d5_71__N_706[47]), .CK(osc_clk), .Q(d5[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i47.GSR = "ENABLED";
    FD1S3AX d5_i48 (.D(d5_71__N_706[48]), .CK(osc_clk), .Q(d5[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i48.GSR = "ENABLED";
    FD1S3AX d5_i49 (.D(d5_71__N_706[49]), .CK(osc_clk), .Q(d5[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i49.GSR = "ENABLED";
    FD1S3AX d5_i50 (.D(d5_71__N_706[50]), .CK(osc_clk), .Q(d5[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i50.GSR = "ENABLED";
    FD1S3AX d5_i51 (.D(d5_71__N_706[51]), .CK(osc_clk), .Q(d5[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i51.GSR = "ENABLED";
    FD1S3AX d5_i52 (.D(d5_71__N_706[52]), .CK(osc_clk), .Q(d5[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i52.GSR = "ENABLED";
    FD1S3AX d5_i53 (.D(d5_71__N_706[53]), .CK(osc_clk), .Q(d5[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i53.GSR = "ENABLED";
    FD1S3AX d5_i54 (.D(d5_71__N_706[54]), .CK(osc_clk), .Q(d5[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i54.GSR = "ENABLED";
    FD1S3AX d5_i55 (.D(d5_71__N_706[55]), .CK(osc_clk), .Q(d5[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i55.GSR = "ENABLED";
    FD1S3AX d5_i56 (.D(d5_71__N_706[56]), .CK(osc_clk), .Q(d5[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i56.GSR = "ENABLED";
    FD1S3AX d5_i57 (.D(d5_71__N_706[57]), .CK(osc_clk), .Q(d5[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i57.GSR = "ENABLED";
    FD1S3AX d5_i58 (.D(d5_71__N_706[58]), .CK(osc_clk), .Q(d5[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i58.GSR = "ENABLED";
    FD1S3AX d5_i59 (.D(d5_71__N_706[59]), .CK(osc_clk), .Q(d5[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i59.GSR = "ENABLED";
    FD1S3AX d5_i60 (.D(d5_71__N_706[60]), .CK(osc_clk), .Q(d5[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i60.GSR = "ENABLED";
    FD1S3AX d5_i61 (.D(d5_71__N_706[61]), .CK(osc_clk), .Q(d5[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i61.GSR = "ENABLED";
    FD1S3AX d5_i62 (.D(d5_71__N_706[62]), .CK(osc_clk), .Q(d5[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i62.GSR = "ENABLED";
    FD1S3AX d5_i63 (.D(d5_71__N_706[63]), .CK(osc_clk), .Q(d5[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i63.GSR = "ENABLED";
    FD1S3AX d5_i64 (.D(d5_71__N_706[64]), .CK(osc_clk), .Q(d5[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i64.GSR = "ENABLED";
    FD1S3AX d5_i65 (.D(d5_71__N_706[65]), .CK(osc_clk), .Q(d5[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i65.GSR = "ENABLED";
    FD1S3AX d5_i66 (.D(d5_71__N_706[66]), .CK(osc_clk), .Q(d5[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i66.GSR = "ENABLED";
    FD1S3AX d5_i67 (.D(d5_71__N_706[67]), .CK(osc_clk), .Q(d5[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i67.GSR = "ENABLED";
    FD1S3AX d5_i68 (.D(d5_71__N_706[68]), .CK(osc_clk), .Q(d5[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i68.GSR = "ENABLED";
    FD1S3AX d5_i69 (.D(d5_71__N_706[69]), .CK(osc_clk), .Q(d5[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i69.GSR = "ENABLED";
    FD1S3AX d5_i70 (.D(d5_71__N_706[70]), .CK(osc_clk), .Q(d5[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i70.GSR = "ENABLED";
    FD1S3AX d5_i71 (.D(d5_71__N_706[71]), .CK(osc_clk), .Q(d5[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i71.GSR = "ENABLED";
    FD1P3AX d6_i0_i1 (.D(d6_71__N_1459[1]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d6_i0_i2 (.D(d6_71__N_1459[2]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d6_i0_i3 (.D(d6_71__N_1459[3]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d6_i0_i4 (.D(d6_71__N_1459[4]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d6_i0_i5 (.D(d6_71__N_1459[5]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d6_i0_i6 (.D(d6_71__N_1459[6]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d6_i0_i7 (.D(d6_71__N_1459[7]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d6_i0_i8 (.D(d6_71__N_1459[8]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d6_i0_i9 (.D(d6_71__N_1459[9]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d6_i0_i10 (.D(d6_71__N_1459[10]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d6_i0_i11 (.D(d6_71__N_1459[11]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d6_i0_i12 (.D(d6_71__N_1459[12]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d6_i0_i13 (.D(d6_71__N_1459[13]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d6_i0_i14 (.D(d6_71__N_1459[14]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d6_i0_i15 (.D(d6_71__N_1459[15]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d6_i0_i16 (.D(d6_71__N_1459[16]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d6_i0_i17 (.D(d6_71__N_1459[17]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d6_i0_i18 (.D(d6_71__N_1459[18]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d6_i0_i19 (.D(d6_71__N_1459[19]), .SP(osc_clk_enable_147), .CK(osc_clk), 
            .Q(d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d6_i0_i20 (.D(d6_71__N_1459[20]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d6_i0_i21 (.D(d6_71__N_1459[21]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d6_i0_i22 (.D(d6_71__N_1459[22]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d6_i0_i23 (.D(d6_71__N_1459[23]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d6_i0_i24 (.D(d6_71__N_1459[24]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d6_i0_i25 (.D(d6_71__N_1459[25]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d6_i0_i26 (.D(d6_71__N_1459[26]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d6_i0_i27 (.D(d6_71__N_1459[27]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d6_i0_i28 (.D(d6_71__N_1459[28]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d6_i0_i29 (.D(d6_71__N_1459[29]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d6_i0_i30 (.D(d6_71__N_1459[30]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d6_i0_i31 (.D(d6_71__N_1459[31]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d6_i0_i32 (.D(d6_71__N_1459[32]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d6_i0_i33 (.D(d6_71__N_1459[33]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d6_i0_i34 (.D(d6_71__N_1459[34]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d6_i0_i35 (.D(d6_71__N_1459[35]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d6_i0_i36 (.D(d6_71__N_1459[36]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d6_i0_i37 (.D(d6_71__N_1459[37]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d6_i0_i38 (.D(d6_71__N_1459[38]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d6_i0_i39 (.D(d6_71__N_1459[39]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d6_i0_i40 (.D(d6_71__N_1459[40]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d6_i0_i41 (.D(d6_71__N_1459[41]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d6_i0_i42 (.D(d6_71__N_1459[42]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d6_i0_i43 (.D(d6_71__N_1459[43]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d6_i0_i44 (.D(d6_71__N_1459[44]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d6_i0_i45 (.D(d6_71__N_1459[45]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d6_i0_i46 (.D(d6_71__N_1459[46]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d6_i0_i47 (.D(d6_71__N_1459[47]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d6_i0_i48 (.D(d6_71__N_1459[48]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d6_i0_i49 (.D(d6_71__N_1459[49]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d6_i0_i50 (.D(d6_71__N_1459[50]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d6_i0_i51 (.D(d6_71__N_1459[51]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d6_i0_i52 (.D(d6_71__N_1459[52]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d6_i0_i53 (.D(d6_71__N_1459[53]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d6_i0_i54 (.D(d6_71__N_1459[54]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d6_i0_i55 (.D(d6_71__N_1459[55]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d6_i0_i56 (.D(d6_71__N_1459[56]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d6_i0_i57 (.D(d6_71__N_1459[57]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d6_i0_i58 (.D(d6_71__N_1459[58]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d6_i0_i59 (.D(d6_71__N_1459[59]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d6_i0_i60 (.D(d6_71__N_1459[60]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d6_i0_i61 (.D(d6_71__N_1459[61]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d6_i0_i62 (.D(d6_71__N_1459[62]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d6_i0_i63 (.D(d6_71__N_1459[63]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d6_i0_i64 (.D(d6_71__N_1459[64]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d6_i0_i65 (.D(d6_71__N_1459[65]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d6_i0_i66 (.D(d6_71__N_1459[66]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d6_i0_i67 (.D(d6_71__N_1459[67]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d6_i0_i68 (.D(d6_71__N_1459[68]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d6_i0_i69 (.D(d6_71__N_1459[69]), .SP(osc_clk_enable_197), .CK(osc_clk), 
            .Q(d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d6_i0_i70 (.D(d6_71__N_1459[70]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d6_i0_i71 (.D(d6_71__N_1459[71]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i1 (.D(d6[1]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i2 (.D(d6[2]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i3 (.D(d6[3]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i4 (.D(d6[4]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i5 (.D(d6[5]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i6 (.D(d6[6]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i7 (.D(d6[7]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i8 (.D(d6[8]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i9 (.D(d6[9]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i10 (.D(d6[10]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i11 (.D(d6[11]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i12 (.D(d6[12]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i13 (.D(d6[13]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i14 (.D(d6[14]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i15 (.D(d6[15]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i16 (.D(d6[16]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i17 (.D(d6[17]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i18 (.D(d6[18]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i19 (.D(d6[19]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i20 (.D(d6[20]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i21 (.D(d6[21]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i22 (.D(d6[22]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i23 (.D(d6[23]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i24 (.D(d6[24]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i25 (.D(d6[25]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i26 (.D(d6[26]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i27 (.D(d6[27]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i28 (.D(d6[28]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i29 (.D(d6[29]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i30 (.D(d6[30]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i31 (.D(d6[31]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i32 (.D(d6[32]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i33 (.D(d6[33]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i34 (.D(d6[34]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i35 (.D(d6[35]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i36 (.D(d6[36]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i37 (.D(d6[37]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i38 (.D(d6[38]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i39 (.D(d6[39]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i40 (.D(d6[40]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i41 (.D(d6[41]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i42 (.D(d6[42]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i43 (.D(d6[43]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i44 (.D(d6[44]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i45 (.D(d6[45]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i46 (.D(d6[46]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i47 (.D(d6[47]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i48 (.D(d6[48]), .SP(osc_clk_enable_247), .CK(osc_clk), 
            .Q(d_d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i49 (.D(d6[49]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d_d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i50 (.D(d6[50]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d_d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i51 (.D(d6[51]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d_d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i52 (.D(d6[52]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d_d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i53 (.D(d6[53]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d_d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i54 (.D(d6[54]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d_d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i55 (.D(d6[55]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d_d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i56 (.D(d6[56]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d_d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i57 (.D(d6[57]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d_d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i58 (.D(d6[58]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d_d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i59 (.D(d6[59]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d_d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i60 (.D(d6[60]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d_d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i61 (.D(d6[61]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d_d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i62 (.D(d6[62]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d_d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i63 (.D(d6[63]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d_d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i64 (.D(d6[64]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d_d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i65 (.D(d6[65]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d_d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i66 (.D(d6[66]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d_d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i67 (.D(d6[67]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d_d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i68 (.D(d6[68]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d_d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i69 (.D(d6[69]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d_d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i70 (.D(d6[70]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d_d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i71 (.D(d6[71]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d_d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d7_i0_i1 (.D(d7_71__N_1531[1]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d7_i0_i2 (.D(d7_71__N_1531[2]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d7_i0_i3 (.D(d7_71__N_1531[3]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d7_i0_i4 (.D(d7_71__N_1531[4]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d7_i0_i5 (.D(d7_71__N_1531[5]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d7_i0_i6 (.D(d7_71__N_1531[6]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d7_i0_i7 (.D(d7_71__N_1531[7]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d7_i0_i8 (.D(d7_71__N_1531[8]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d7_i0_i9 (.D(d7_71__N_1531[9]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d7_i0_i10 (.D(d7_71__N_1531[10]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d7_i0_i11 (.D(d7_71__N_1531[11]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d7_i0_i12 (.D(d7_71__N_1531[12]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d7_i0_i13 (.D(d7_71__N_1531[13]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d7_i0_i14 (.D(d7_71__N_1531[14]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d7_i0_i15 (.D(d7_71__N_1531[15]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d7_i0_i16 (.D(d7_71__N_1531[16]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d7_i0_i17 (.D(d7_71__N_1531[17]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d7_i0_i18 (.D(d7_71__N_1531[18]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d7_i0_i19 (.D(d7_71__N_1531[19]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d7_i0_i20 (.D(d7_71__N_1531[20]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d7_i0_i21 (.D(d7_71__N_1531[21]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d7_i0_i22 (.D(d7_71__N_1531[22]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d7_i0_i23 (.D(d7_71__N_1531[23]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d7_i0_i24 (.D(d7_71__N_1531[24]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d7_i0_i25 (.D(d7_71__N_1531[25]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d7_i0_i26 (.D(d7_71__N_1531[26]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d7_i0_i27 (.D(d7_71__N_1531[27]), .SP(osc_clk_enable_297), .CK(osc_clk), 
            .Q(d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d7_i0_i28 (.D(d7_71__N_1531[28]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d7_i0_i29 (.D(d7_71__N_1531[29]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d7_i0_i30 (.D(d7_71__N_1531[30]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d7_i0_i31 (.D(d7_71__N_1531[31]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d7_i0_i32 (.D(d7_71__N_1531[32]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d7_i0_i33 (.D(d7_71__N_1531[33]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d7_i0_i34 (.D(d7_71__N_1531[34]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d7_i0_i35 (.D(d7_71__N_1531[35]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d7_i0_i36 (.D(d7_71__N_1531[36]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d7_i0_i37 (.D(d7_71__N_1531[37]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d7_i0_i38 (.D(d7_71__N_1531[38]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d7_i0_i39 (.D(d7_71__N_1531[39]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d7_i0_i40 (.D(d7_71__N_1531[40]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d7_i0_i41 (.D(d7_71__N_1531[41]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d7_i0_i42 (.D(d7_71__N_1531[42]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d7_i0_i43 (.D(d7_71__N_1531[43]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d7_i0_i44 (.D(d7_71__N_1531[44]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d7_i0_i45 (.D(d7_71__N_1531[45]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d7_i0_i46 (.D(d7_71__N_1531[46]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d7_i0_i47 (.D(d7_71__N_1531[47]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d7_i0_i48 (.D(d7_71__N_1531[48]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d7_i0_i49 (.D(d7_71__N_1531[49]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d7_i0_i50 (.D(d7_71__N_1531[50]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d7_i0_i51 (.D(d7_71__N_1531[51]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d7_i0_i52 (.D(d7_71__N_1531[52]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d7_i0_i53 (.D(d7_71__N_1531[53]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d7_i0_i54 (.D(d7_71__N_1531[54]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d7_i0_i55 (.D(d7_71__N_1531[55]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d7_i0_i56 (.D(d7_71__N_1531[56]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d7_i0_i57 (.D(d7_71__N_1531[57]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d7_i0_i58 (.D(d7_71__N_1531[58]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d7_i0_i59 (.D(d7_71__N_1531[59]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d7_i0_i60 (.D(d7_71__N_1531[60]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d7_i0_i61 (.D(d7_71__N_1531[61]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d7_i0_i62 (.D(d7_71__N_1531[62]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d7_i0_i63 (.D(d7_71__N_1531[63]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d7_i0_i64 (.D(d7_71__N_1531[64]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d7_i0_i65 (.D(d7_71__N_1531[65]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d7_i0_i66 (.D(d7_71__N_1531[66]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d7_i0_i67 (.D(d7_71__N_1531[67]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d7_i0_i68 (.D(d7_71__N_1531[68]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d7_i0_i69 (.D(d7_71__N_1531[69]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d7_i0_i70 (.D(d7_71__N_1531[70]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d7_i0_i71 (.D(d7_71__N_1531[71]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i1 (.D(d7[1]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d_d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i2 (.D(d7[2]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d_d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i3 (.D(d7[3]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d_d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i4 (.D(d7[4]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d_d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i5 (.D(d7[5]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d_d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i6 (.D(d7[6]), .SP(osc_clk_enable_347), .CK(osc_clk), 
            .Q(d_d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i7 (.D(d7[7]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i8 (.D(d7[8]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i9 (.D(d7[9]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i10 (.D(d7[10]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i11 (.D(d7[11]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i12 (.D(d7[12]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i13 (.D(d7[13]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i14 (.D(d7[14]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i15 (.D(d7[15]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i16 (.D(d7[16]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i17 (.D(d7[17]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i18 (.D(d7[18]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i19 (.D(d7[19]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i20 (.D(d7[20]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i21 (.D(d7[21]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i22 (.D(d7[22]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i23 (.D(d7[23]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i24 (.D(d7[24]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i25 (.D(d7[25]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i26 (.D(d7[26]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i27 (.D(d7[27]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i28 (.D(d7[28]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i29 (.D(d7[29]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i30 (.D(d7[30]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i31 (.D(d7[31]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i32 (.D(d7[32]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i33 (.D(d7[33]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i34 (.D(d7[34]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i35 (.D(d7[35]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i36 (.D(d7[36]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i37 (.D(d7[37]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i38 (.D(d7[38]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i39 (.D(d7[39]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i40 (.D(d7[40]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i41 (.D(d7[41]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i42 (.D(d7[42]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i43 (.D(d7[43]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i44 (.D(d7[44]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i45 (.D(d7[45]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i46 (.D(d7[46]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i47 (.D(d7[47]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i48 (.D(d7[48]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i49 (.D(d7[49]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i50 (.D(d7[50]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i51 (.D(d7[51]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i52 (.D(d7[52]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i53 (.D(d7[53]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i54 (.D(d7[54]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i55 (.D(d7[55]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i56 (.D(d7[56]), .SP(osc_clk_enable_397), .CK(osc_clk), 
            .Q(d_d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i57 (.D(d7[57]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d_d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i58 (.D(d7[58]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d_d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i59 (.D(d7[59]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d_d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i60 (.D(d7[60]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d_d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i61 (.D(d7[61]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d_d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i62 (.D(d7[62]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d_d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i63 (.D(d7[63]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d_d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i64 (.D(d7[64]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d_d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i65 (.D(d7[65]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d_d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i66 (.D(d7[66]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d_d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i67 (.D(d7[67]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d_d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i68 (.D(d7[68]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d_d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i69 (.D(d7[69]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d_d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i70 (.D(d7[70]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d_d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i71 (.D(d7[71]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d_d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d8_i0_i1 (.D(d8_71__N_1603[1]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d8_i0_i2 (.D(d8_71__N_1603[2]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d8_i0_i3 (.D(d8_71__N_1603[3]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d8_i0_i4 (.D(d8_71__N_1603[4]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d8_i0_i5 (.D(d8_71__N_1603[5]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d8_i0_i6 (.D(d8_71__N_1603[6]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d8_i0_i7 (.D(d8_71__N_1603[7]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d8_i0_i8 (.D(d8_71__N_1603[8]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d8_i0_i9 (.D(d8_71__N_1603[9]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d8_i0_i10 (.D(d8_71__N_1603[10]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d8_i0_i11 (.D(d8_71__N_1603[11]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d8_i0_i12 (.D(d8_71__N_1603[12]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d8_i0_i13 (.D(d8_71__N_1603[13]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d8_i0_i14 (.D(d8_71__N_1603[14]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d8_i0_i15 (.D(d8_71__N_1603[15]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d8_i0_i16 (.D(d8_71__N_1603[16]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d8_i0_i17 (.D(d8_71__N_1603[17]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d8_i0_i18 (.D(d8_71__N_1603[18]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d8_i0_i19 (.D(d8_71__N_1603[19]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d8_i0_i20 (.D(d8_71__N_1603[20]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d8_i0_i21 (.D(d8_71__N_1603[21]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d8_i0_i22 (.D(d8_71__N_1603[22]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d8_i0_i23 (.D(d8_71__N_1603[23]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d8_i0_i24 (.D(d8_71__N_1603[24]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d8_i0_i25 (.D(d8_71__N_1603[25]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d8_i0_i26 (.D(d8_71__N_1603[26]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d8_i0_i27 (.D(d8_71__N_1603[27]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d8_i0_i28 (.D(d8_71__N_1603[28]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d8_i0_i29 (.D(d8_71__N_1603[29]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d8_i0_i30 (.D(d8_71__N_1603[30]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d8_i0_i31 (.D(d8_71__N_1603[31]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d8_i0_i32 (.D(d8_71__N_1603[32]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d8_i0_i33 (.D(d8_71__N_1603[33]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d8_i0_i34 (.D(d8_71__N_1603[34]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d8_i0_i35 (.D(d8_71__N_1603[35]), .SP(osc_clk_enable_447), .CK(osc_clk), 
            .Q(d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d8_i0_i36 (.D(d8_71__N_1603[36]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d8_i0_i37 (.D(d8_71__N_1603[37]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d8_i0_i38 (.D(d8_71__N_1603[38]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d8_i0_i39 (.D(d8_71__N_1603[39]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d8_i0_i40 (.D(d8_71__N_1603[40]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d8_i0_i41 (.D(d8_71__N_1603[41]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d8_i0_i42 (.D(d8_71__N_1603[42]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d8_i0_i43 (.D(d8_71__N_1603[43]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d8_i0_i44 (.D(d8_71__N_1603[44]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d8_i0_i45 (.D(d8_71__N_1603[45]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d8_i0_i46 (.D(d8_71__N_1603[46]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d8_i0_i47 (.D(d8_71__N_1603[47]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d8_i0_i48 (.D(d8_71__N_1603[48]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d8_i0_i49 (.D(d8_71__N_1603[49]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d8_i0_i50 (.D(d8_71__N_1603[50]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d8_i0_i51 (.D(d8_71__N_1603[51]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d8_i0_i52 (.D(d8_71__N_1603[52]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d8_i0_i53 (.D(d8_71__N_1603[53]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d8_i0_i54 (.D(d8_71__N_1603[54]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d8_i0_i55 (.D(d8_71__N_1603[55]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d8_i0_i56 (.D(d8_71__N_1603[56]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d8_i0_i57 (.D(d8_71__N_1603[57]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d8_i0_i58 (.D(d8_71__N_1603[58]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d8_i0_i59 (.D(d8_71__N_1603[59]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d8_i0_i60 (.D(d8_71__N_1603[60]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d8_i0_i61 (.D(d8_71__N_1603[61]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d8_i0_i62 (.D(d8_71__N_1603[62]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d8_i0_i63 (.D(d8_71__N_1603[63]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d8_i0_i64 (.D(d8_71__N_1603[64]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d8_i0_i65 (.D(d8_71__N_1603[65]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d8_i0_i66 (.D(d8_71__N_1603[66]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d8_i0_i67 (.D(d8_71__N_1603[67]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d8_i0_i68 (.D(d8_71__N_1603[68]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d8_i0_i69 (.D(d8_71__N_1603[69]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d8_i0_i70 (.D(d8_71__N_1603[70]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d8_i0_i71 (.D(d8_71__N_1603[71]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i1 (.D(d8[1]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d_d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i2 (.D(d8[2]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d_d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i3 (.D(d8[3]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d_d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i4 (.D(d8[4]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d_d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i5 (.D(d8[5]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d_d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i6 (.D(d8[6]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d_d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i7 (.D(d8[7]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d_d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i8 (.D(d8[8]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d_d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i9 (.D(d8[9]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d_d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i10 (.D(d8[10]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d_d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i11 (.D(d8[11]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d_d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i12 (.D(d8[12]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d_d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i13 (.D(d8[13]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d_d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i14 (.D(d8[14]), .SP(osc_clk_enable_497), .CK(osc_clk), 
            .Q(d_d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i15 (.D(d8[15]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i16 (.D(d8[16]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i17 (.D(d8[17]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i18 (.D(d8[18]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i19 (.D(d8[19]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i20 (.D(d8[20]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i21 (.D(d8[21]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i22 (.D(d8[22]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i23 (.D(d8[23]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i24 (.D(d8[24]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i25 (.D(d8[25]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i26 (.D(d8[26]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i27 (.D(d8[27]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i28 (.D(d8[28]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i29 (.D(d8[29]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i30 (.D(d8[30]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i31 (.D(d8[31]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i32 (.D(d8[32]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i33 (.D(d8[33]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i34 (.D(d8[34]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i35 (.D(d8[35]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i36 (.D(d8[36]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i37 (.D(d8[37]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i38 (.D(d8[38]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i39 (.D(d8[39]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i40 (.D(d8[40]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i41 (.D(d8[41]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i42 (.D(d8[42]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i43 (.D(d8[43]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i44 (.D(d8[44]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i45 (.D(d8[45]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i46 (.D(d8[46]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i47 (.D(d8[47]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i48 (.D(d8[48]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i49 (.D(d8[49]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i50 (.D(d8[50]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i51 (.D(d8[51]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i52 (.D(d8[52]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i53 (.D(d8[53]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i54 (.D(d8[54]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i55 (.D(d8[55]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i56 (.D(d8[56]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i57 (.D(d8[57]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i58 (.D(d8[58]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i59 (.D(d8[59]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i60 (.D(d8[60]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i61 (.D(d8[61]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i62 (.D(d8[62]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i63 (.D(d8[63]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i64 (.D(d8[64]), .SP(osc_clk_enable_547), .CK(osc_clk), 
            .Q(d_d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i65 (.D(d8[65]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d_d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i66 (.D(d8[66]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d_d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i67 (.D(d8[67]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d_d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i68 (.D(d8[68]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d_d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i69 (.D(d8[69]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d_d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i70 (.D(d8[70]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d_d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i71 (.D(d8[71]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d_d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d9_i0_i1 (.D(d9_71__N_1675[1]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d9_i0_i2 (.D(d9_71__N_1675[2]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d9_i0_i3 (.D(d9_71__N_1675[3]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d9_i0_i4 (.D(d9_71__N_1675[4]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d9_i0_i5 (.D(d9_71__N_1675[5]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d9_i0_i6 (.D(d9_71__N_1675[6]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d9_i0_i7 (.D(d9_71__N_1675[7]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d9_i0_i8 (.D(d9_71__N_1675[8]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d9_i0_i9 (.D(d9_71__N_1675[9]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d9_i0_i10 (.D(d9_71__N_1675[10]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d9_i0_i11 (.D(d9_71__N_1675[11]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d9_i0_i12 (.D(d9_71__N_1675[12]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d9_i0_i13 (.D(d9_71__N_1675[13]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d9_i0_i14 (.D(d9_71__N_1675[14]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d9_i0_i15 (.D(d9_71__N_1675[15]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d9_i0_i16 (.D(d9_71__N_1675[16]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d9_i0_i17 (.D(d9_71__N_1675[17]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d9_i0_i18 (.D(d9_71__N_1675[18]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d9_i0_i19 (.D(d9_71__N_1675[19]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d9_i0_i20 (.D(d9_71__N_1675[20]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d9_i0_i21 (.D(d9_71__N_1675[21]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d9_i0_i22 (.D(d9_71__N_1675[22]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d9_i0_i23 (.D(d9_71__N_1675[23]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d9_i0_i24 (.D(d9_71__N_1675[24]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d9_i0_i25 (.D(d9_71__N_1675[25]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d9_i0_i26 (.D(d9_71__N_1675[26]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d9_i0_i27 (.D(d9_71__N_1675[27]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d9_i0_i28 (.D(d9_71__N_1675[28]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d9_i0_i29 (.D(d9_71__N_1675[29]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d9_i0_i30 (.D(d9_71__N_1675[30]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d9_i0_i31 (.D(d9_71__N_1675[31]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d9_i0_i32 (.D(d9_71__N_1675[32]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d9_i0_i33 (.D(d9_71__N_1675[33]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d9_i0_i34 (.D(d9_71__N_1675[34]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d9_i0_i35 (.D(d9_71__N_1675[35]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d9_i0_i36 (.D(d9_71__N_1675[36]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d9_i0_i37 (.D(d9_71__N_1675[37]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d9_i0_i38 (.D(d9_71__N_1675[38]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d9_i0_i39 (.D(d9_71__N_1675[39]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d9_i0_i40 (.D(d9_71__N_1675[40]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d9_i0_i41 (.D(d9_71__N_1675[41]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d9_i0_i42 (.D(d9_71__N_1675[42]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d9_i0_i43 (.D(d9_71__N_1675[43]), .SP(osc_clk_enable_597), .CK(osc_clk), 
            .Q(d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d9_i0_i44 (.D(d9_71__N_1675[44]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d9_i0_i45 (.D(d9_71__N_1675[45]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d9_i0_i46 (.D(d9_71__N_1675[46]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d9_i0_i47 (.D(d9_71__N_1675[47]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d9_i0_i48 (.D(d9_71__N_1675[48]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d9_i0_i49 (.D(d9_71__N_1675[49]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d9_i0_i50 (.D(d9_71__N_1675[50]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d9_i0_i51 (.D(d9_71__N_1675[51]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d9_i0_i52 (.D(d9_71__N_1675[52]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d9_i0_i53 (.D(d9_71__N_1675[53]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d9_i0_i54 (.D(d9_71__N_1675[54]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d9_i0_i55 (.D(d9_71__N_1675[55]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d9_i0_i56 (.D(d9_71__N_1675[56]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d9_i0_i57 (.D(d9_71__N_1675[57]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d9_i0_i58 (.D(d9_71__N_1675[58]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d9_i0_i59 (.D(d9_71__N_1675[59]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d9_i0_i60 (.D(d9_71__N_1675[60]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d9_i0_i61 (.D(d9_71__N_1675[61]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d9_i0_i62 (.D(d9_71__N_1675[62]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d9_i0_i63 (.D(d9_71__N_1675[63]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d9_i0_i64 (.D(d9_71__N_1675[64]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d9_i0_i65 (.D(d9_71__N_1675[65]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d9_i0_i66 (.D(d9_71__N_1675[66]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d9_i0_i67 (.D(d9_71__N_1675[67]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d9_i0_i68 (.D(d9_71__N_1675[68]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d9_i0_i69 (.D(d9_71__N_1675[69]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d9_i0_i70 (.D(d9_71__N_1675[70]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d9_i0_i71 (.D(d9_71__N_1675[71]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i1 (.D(d9[1]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d_d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i2 (.D(d9[2]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d_d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i3 (.D(d9[3]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d_d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i4 (.D(d9[4]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d_d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i5 (.D(d9[5]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d_d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i6 (.D(d9[6]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d_d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i7 (.D(d9[7]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d_d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i8 (.D(d9[8]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d_d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i9 (.D(d9[9]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d_d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i10 (.D(d9[10]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d_d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i11 (.D(d9[11]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d_d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i12 (.D(d9[12]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d_d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i13 (.D(d9[13]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d_d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i14 (.D(d9[14]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d_d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i15 (.D(d9[15]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d_d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i16 (.D(d9[16]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d_d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i17 (.D(d9[17]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d_d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i18 (.D(d9[18]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d_d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i19 (.D(d9[19]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d_d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i20 (.D(d9[20]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d_d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i21 (.D(d9[21]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d_d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i22 (.D(d9[22]), .SP(osc_clk_enable_647), .CK(osc_clk), 
            .Q(d_d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i23 (.D(d9[23]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i24 (.D(d9[24]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i25 (.D(d9[25]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i26 (.D(d9[26]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i27 (.D(d9[27]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i28 (.D(d9[28]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i29 (.D(d9[29]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i30 (.D(d9[30]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i31 (.D(d9[31]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i32 (.D(d9[32]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i33 (.D(d9[33]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i34 (.D(d9[34]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i35 (.D(d9[35]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i36 (.D(d9[36]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i37 (.D(d9[37]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i38 (.D(d9[38]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i39 (.D(d9[39]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i40 (.D(d9[40]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i41 (.D(d9[41]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i42 (.D(d9[42]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i43 (.D(d9[43]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i44 (.D(d9[44]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i45 (.D(d9[45]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i46 (.D(d9[46]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i47 (.D(d9[47]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i48 (.D(d9[48]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i49 (.D(d9[49]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i50 (.D(d9[50]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i51 (.D(d9[51]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i52 (.D(d9[52]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i53 (.D(d9[53]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i54 (.D(d9[54]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i55 (.D(d9[55]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i56 (.D(d9[56]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i57 (.D(d9[57]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i58 (.D(d9[58]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i59 (.D(d9[59]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i60 (.D(d9[60]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i61 (.D(d9[61]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i62 (.D(d9[62]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i63 (.D(d9[63]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i64 (.D(d9[64]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i65 (.D(d9[65]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i66 (.D(d9[66]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i67 (.D(d9[67]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i68 (.D(d9[68]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i69 (.D(d9[69]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i70 (.D(d9[70]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i71 (.D(d9[71]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d_d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d10__i2 (.D(d10_71__N_1747[57]), .SP(osc_clk_enable_697), .CK(osc_clk), 
            .Q(d10[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i2.GSR = "ENABLED";
    FD1P3AX d10__i3 (.D(d10_71__N_1747[58]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i3.GSR = "ENABLED";
    FD1P3AX d10__i4 (.D(d10_71__N_1747[59]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i4.GSR = "ENABLED";
    FD1P3AX d10__i5 (.D(d10_71__N_1747[60]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i5.GSR = "ENABLED";
    FD1P3AX d10__i6 (.D(d10_71__N_1747[61]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i6.GSR = "ENABLED";
    FD1P3AX d10__i7 (.D(d10_71__N_1747[62]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i7.GSR = "ENABLED";
    FD1P3AX d10__i8 (.D(d10_71__N_1747[63]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i8.GSR = "ENABLED";
    FD1P3AX d10__i9 (.D(d10_71__N_1747[64]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i9.GSR = "ENABLED";
    FD1P3AX d10__i10 (.D(d10_71__N_1747[65]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i10.GSR = "ENABLED";
    FD1P3AX d10__i11 (.D(d10_71__N_1747[66]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i11.GSR = "ENABLED";
    FD1P3AX d10__i12 (.D(d10_71__N_1747[67]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i12.GSR = "ENABLED";
    FD1P3AX d10__i13 (.D(d10_71__N_1747[68]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i13.GSR = "ENABLED";
    FD1P3AX d10__i14 (.D(d10_71__N_1747[69]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i14.GSR = "ENABLED";
    FD1P3AX d10__i15 (.D(d10_71__N_1747[70]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i15.GSR = "ENABLED";
    FD1P3AX d10__i16 (.D(d10_71__N_1747[71]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i16.GSR = "ENABLED";
    FD1P3AX d_out_i0_i1 (.D(d_out_11__N_1819[1]), .SP(v_comb), .CK(osc_clk), 
            .Q(\CIC1_outSin[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i1.GSR = "ENABLED";
    FD1P3AX d_out_i0_i2 (.D(d_out_11__N_1819[2]), .SP(v_comb), .CK(osc_clk), 
            .Q(\CIC1_outSin[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i2.GSR = "ENABLED";
    FD1P3AX d_out_i0_i3 (.D(d_out_11__N_1819[3]), .SP(v_comb), .CK(osc_clk), 
            .Q(\CIC1_outSin[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i3.GSR = "ENABLED";
    FD1P3AX d_out_i0_i4 (.D(d_out_11__N_1819[4]), .SP(v_comb), .CK(osc_clk), 
            .Q(\CIC1_outSin[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i4.GSR = "ENABLED";
    FD1P3AX d_out_i0_i5 (.D(d_out_11__N_1819[5]), .SP(v_comb), .CK(osc_clk), 
            .Q(\CIC1_outSin[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i5.GSR = "ENABLED";
    FD1P3AX d_out_i0_i6 (.D(d_out_11__N_1819[6]), .SP(v_comb), .CK(osc_clk), 
            .Q(MYLED_c_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i6.GSR = "ENABLED";
    FD1P3AX d_out_i0_i7 (.D(d_out_11__N_1819[7]), .SP(v_comb), .CK(osc_clk), 
            .Q(MYLED_c_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i7.GSR = "ENABLED";
    FD1P3AX d_out_i0_i8 (.D(d_out_11__N_1819[8]), .SP(v_comb), .CK(osc_clk), 
            .Q(MYLED_c_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i8.GSR = "ENABLED";
    FD1P3AX d_out_i0_i9 (.D(d_out_11__N_1819[9]), .SP(v_comb), .CK(osc_clk), 
            .Q(MYLED_c_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i9.GSR = "ENABLED";
    FD1P3AX d_out_i0_i10 (.D(d_out_11__N_1819[10]), .SP(v_comb), .CK(osc_clk), 
            .Q(MYLED_c_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i10.GSR = "ENABLED";
    FD1P3AX d_out_i0_i11 (.D(d_out_11__N_1819[11]), .SP(v_comb), .CK(osc_clk), 
            .Q(MYLED_c_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i11.GSR = "ENABLED";
    FD1S3AX d1_i1 (.D(d1_71__N_418[1]), .CK(osc_clk), .Q(d1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i1.GSR = "ENABLED";
    FD1S3AX d1_i2 (.D(d1_71__N_418[2]), .CK(osc_clk), .Q(d1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i2.GSR = "ENABLED";
    FD1S3AX d1_i3 (.D(d1_71__N_418[3]), .CK(osc_clk), .Q(d1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i3.GSR = "ENABLED";
    FD1S3AX d1_i4 (.D(d1_71__N_418[4]), .CK(osc_clk), .Q(d1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i4.GSR = "ENABLED";
    FD1S3AX d1_i5 (.D(d1_71__N_418[5]), .CK(osc_clk), .Q(d1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i5.GSR = "ENABLED";
    FD1S3AX d1_i6 (.D(d1_71__N_418[6]), .CK(osc_clk), .Q(d1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i6.GSR = "ENABLED";
    FD1S3AX d1_i7 (.D(d1_71__N_418[7]), .CK(osc_clk), .Q(d1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i7.GSR = "ENABLED";
    FD1S3AX d1_i8 (.D(d1_71__N_418[8]), .CK(osc_clk), .Q(d1[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i8.GSR = "ENABLED";
    FD1S3AX d1_i9 (.D(d1_71__N_418[9]), .CK(osc_clk), .Q(d1[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i9.GSR = "ENABLED";
    FD1S3AX d1_i10 (.D(d1_71__N_418[10]), .CK(osc_clk), .Q(d1[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i10.GSR = "ENABLED";
    FD1S3AX d1_i11 (.D(d1_71__N_418[11]), .CK(osc_clk), .Q(d1[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i11.GSR = "ENABLED";
    FD1S3AX d1_i12 (.D(d1_71__N_418[12]), .CK(osc_clk), .Q(d1[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i12.GSR = "ENABLED";
    FD1S3AX d1_i13 (.D(d1_71__N_418[13]), .CK(osc_clk), .Q(d1[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i13.GSR = "ENABLED";
    FD1S3AX d1_i14 (.D(d1_71__N_418[14]), .CK(osc_clk), .Q(d1[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i14.GSR = "ENABLED";
    FD1S3AX d1_i15 (.D(d1_71__N_418[15]), .CK(osc_clk), .Q(d1[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i15.GSR = "ENABLED";
    FD1S3AX d1_i16 (.D(d1_71__N_418[16]), .CK(osc_clk), .Q(d1[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i16.GSR = "ENABLED";
    FD1S3AX d1_i17 (.D(d1_71__N_418[17]), .CK(osc_clk), .Q(d1[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i17.GSR = "ENABLED";
    FD1S3AX d1_i18 (.D(d1_71__N_418[18]), .CK(osc_clk), .Q(d1[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i18.GSR = "ENABLED";
    FD1S3AX d1_i19 (.D(d1_71__N_418[19]), .CK(osc_clk), .Q(d1[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i19.GSR = "ENABLED";
    FD1S3AX d1_i20 (.D(d1_71__N_418[20]), .CK(osc_clk), .Q(d1[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i20.GSR = "ENABLED";
    FD1S3AX d1_i21 (.D(d1_71__N_418[21]), .CK(osc_clk), .Q(d1[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i21.GSR = "ENABLED";
    FD1S3AX d1_i22 (.D(d1_71__N_418[22]), .CK(osc_clk), .Q(d1[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i22.GSR = "ENABLED";
    FD1S3AX d1_i23 (.D(d1_71__N_418[23]), .CK(osc_clk), .Q(d1[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i23.GSR = "ENABLED";
    FD1S3AX d1_i24 (.D(d1_71__N_418[24]), .CK(osc_clk), .Q(d1[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i24.GSR = "ENABLED";
    FD1S3AX d1_i25 (.D(d1_71__N_418[25]), .CK(osc_clk), .Q(d1[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i25.GSR = "ENABLED";
    FD1S3AX d1_i26 (.D(d1_71__N_418[26]), .CK(osc_clk), .Q(d1[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i26.GSR = "ENABLED";
    FD1S3AX d1_i27 (.D(d1_71__N_418[27]), .CK(osc_clk), .Q(d1[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i27.GSR = "ENABLED";
    FD1S3AX d1_i28 (.D(d1_71__N_418[28]), .CK(osc_clk), .Q(d1[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i28.GSR = "ENABLED";
    FD1S3AX d1_i29 (.D(d1_71__N_418[29]), .CK(osc_clk), .Q(d1[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i29.GSR = "ENABLED";
    FD1S3AX d1_i30 (.D(d1_71__N_418[30]), .CK(osc_clk), .Q(d1[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i30.GSR = "ENABLED";
    FD1S3AX d1_i31 (.D(d1_71__N_418[31]), .CK(osc_clk), .Q(d1[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i31.GSR = "ENABLED";
    FD1S3AX d1_i32 (.D(d1_71__N_418[32]), .CK(osc_clk), .Q(d1[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i32.GSR = "ENABLED";
    FD1S3AX d1_i33 (.D(d1_71__N_418[33]), .CK(osc_clk), .Q(d1[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i33.GSR = "ENABLED";
    FD1S3AX d1_i34 (.D(d1_71__N_418[34]), .CK(osc_clk), .Q(d1[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i34.GSR = "ENABLED";
    FD1S3AX d1_i35 (.D(d1_71__N_418[35]), .CK(osc_clk), .Q(d1[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i35.GSR = "ENABLED";
    FD1S3AX d1_i36 (.D(d1_71__N_418[36]), .CK(osc_clk), .Q(d1[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i36.GSR = "ENABLED";
    FD1S3AX d1_i37 (.D(d1_71__N_418[37]), .CK(osc_clk), .Q(d1[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i37.GSR = "ENABLED";
    FD1S3AX d1_i38 (.D(d1_71__N_418[38]), .CK(osc_clk), .Q(d1[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i38.GSR = "ENABLED";
    FD1S3AX d1_i39 (.D(d1_71__N_418[39]), .CK(osc_clk), .Q(d1[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i39.GSR = "ENABLED";
    FD1S3AX d1_i40 (.D(d1_71__N_418[40]), .CK(osc_clk), .Q(d1[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i40.GSR = "ENABLED";
    FD1S3AX d1_i41 (.D(d1_71__N_418[41]), .CK(osc_clk), .Q(d1[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i41.GSR = "ENABLED";
    FD1S3AX d1_i42 (.D(d1_71__N_418[42]), .CK(osc_clk), .Q(d1[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i42.GSR = "ENABLED";
    FD1S3AX d1_i43 (.D(d1_71__N_418[43]), .CK(osc_clk), .Q(d1[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i43.GSR = "ENABLED";
    FD1S3AX d1_i44 (.D(d1_71__N_418[44]), .CK(osc_clk), .Q(d1[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i44.GSR = "ENABLED";
    FD1S3AX d1_i45 (.D(d1_71__N_418[45]), .CK(osc_clk), .Q(d1[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i45.GSR = "ENABLED";
    FD1S3AX d1_i46 (.D(d1_71__N_418[46]), .CK(osc_clk), .Q(d1[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i46.GSR = "ENABLED";
    FD1S3AX d1_i47 (.D(d1_71__N_418[47]), .CK(osc_clk), .Q(d1[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i47.GSR = "ENABLED";
    FD1S3AX d1_i48 (.D(d1_71__N_418[48]), .CK(osc_clk), .Q(d1[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i48.GSR = "ENABLED";
    FD1S3AX d1_i49 (.D(d1_71__N_418[49]), .CK(osc_clk), .Q(d1[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i49.GSR = "ENABLED";
    FD1S3AX d1_i50 (.D(d1_71__N_418[50]), .CK(osc_clk), .Q(d1[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i50.GSR = "ENABLED";
    FD1S3AX d1_i51 (.D(d1_71__N_418[51]), .CK(osc_clk), .Q(d1[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i51.GSR = "ENABLED";
    FD1S3AX d1_i52 (.D(d1_71__N_418[52]), .CK(osc_clk), .Q(d1[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i52.GSR = "ENABLED";
    FD1S3AX d1_i53 (.D(d1_71__N_418[53]), .CK(osc_clk), .Q(d1[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i53.GSR = "ENABLED";
    FD1S3AX d1_i54 (.D(d1_71__N_418[54]), .CK(osc_clk), .Q(d1[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i54.GSR = "ENABLED";
    FD1S3AX d1_i55 (.D(d1_71__N_418[55]), .CK(osc_clk), .Q(d1[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i55.GSR = "ENABLED";
    FD1S3AX d1_i56 (.D(d1_71__N_418[56]), .CK(osc_clk), .Q(d1[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i56.GSR = "ENABLED";
    FD1S3AX d1_i57 (.D(d1_71__N_418[57]), .CK(osc_clk), .Q(d1[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i57.GSR = "ENABLED";
    FD1S3AX d1_i58 (.D(d1_71__N_418[58]), .CK(osc_clk), .Q(d1[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i58.GSR = "ENABLED";
    FD1S3AX d1_i59 (.D(d1_71__N_418[59]), .CK(osc_clk), .Q(d1[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i59.GSR = "ENABLED";
    FD1S3AX d1_i60 (.D(d1_71__N_418[60]), .CK(osc_clk), .Q(d1[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i60.GSR = "ENABLED";
    FD1S3AX d1_i61 (.D(d1_71__N_418[61]), .CK(osc_clk), .Q(d1[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i61.GSR = "ENABLED";
    FD1S3AX d1_i62 (.D(d1_71__N_418[62]), .CK(osc_clk), .Q(d1[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i62.GSR = "ENABLED";
    FD1S3AX d1_i63 (.D(d1_71__N_418[63]), .CK(osc_clk), .Q(d1[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i63.GSR = "ENABLED";
    FD1S3AX d1_i64 (.D(d1_71__N_418[64]), .CK(osc_clk), .Q(d1[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i64.GSR = "ENABLED";
    FD1S3AX d1_i65 (.D(d1_71__N_418[65]), .CK(osc_clk), .Q(d1[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i65.GSR = "ENABLED";
    FD1S3AX d1_i66 (.D(d1_71__N_418[66]), .CK(osc_clk), .Q(d1[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i66.GSR = "ENABLED";
    FD1S3AX d1_i67 (.D(d1_71__N_418[67]), .CK(osc_clk), .Q(d1[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i67.GSR = "ENABLED";
    FD1S3AX d1_i68 (.D(d1_71__N_418[68]), .CK(osc_clk), .Q(d1[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i68.GSR = "ENABLED";
    FD1S3AX d1_i69 (.D(d1_71__N_418[69]), .CK(osc_clk), .Q(d1[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i69.GSR = "ENABLED";
    FD1S3AX d1_i70 (.D(d1_71__N_418[70]), .CK(osc_clk), .Q(d1[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i70.GSR = "ENABLED";
    FD1S3AX d1_i71 (.D(d1_71__N_418[71]), .CK(osc_clk), .Q(d1[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i71.GSR = "ENABLED";
    CCU2D add_1049_6 (.A0(d1[40]), .B0(d2[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[41]), .B1(d2[41]), .C1(GND_net), .D1(GND_net), .CIN(n12233), 
          .COUT(n12234), .S0(n4429[4]), .S1(n4429[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1049_6.INIT0 = 16'h5666;
    defparam add_1049_6.INIT1 = 16'h5666;
    defparam add_1049_6.INJECT1_0 = "NO";
    defparam add_1049_6.INJECT1_1 = "NO";
    CCU2D add_1049_4 (.A0(d1[38]), .B0(d2[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[39]), .B1(d2[39]), .C1(GND_net), .D1(GND_net), .CIN(n12232), 
          .COUT(n12233), .S0(n4429[2]), .S1(n4429[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1049_4.INIT0 = 16'h5666;
    defparam add_1049_4.INIT1 = 16'h5666;
    defparam add_1049_4.INJECT1_0 = "NO";
    defparam add_1049_4.INJECT1_1 = "NO";
    CCU2D add_1049_2 (.A0(d1[36]), .B0(d2[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[37]), .B1(d2[37]), .C1(GND_net), .D1(GND_net), .COUT(n12232), 
          .S1(n4429[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1049_2.INIT0 = 16'h7000;
    defparam add_1049_2.INIT1 = 16'h5666;
    defparam add_1049_2.INJECT1_0 = "NO";
    defparam add_1049_2.INJECT1_1 = "NO";
    CCU2D add_1050_37 (.A0(d2[70]), .B0(n4428), .C0(n4429[34]), .D0(d1[70]), 
          .A1(d2[71]), .B1(n4428), .C1(n4429[35]), .D1(d1[71]), .CIN(n12229), 
          .S0(d2_71__N_490[70]), .S1(d2_71__N_490[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1050_37.INIT0 = 16'h74b8;
    defparam add_1050_37.INIT1 = 16'h74b8;
    defparam add_1050_37.INJECT1_0 = "NO";
    defparam add_1050_37.INJECT1_1 = "NO";
    CCU2D add_1050_35 (.A0(d2[68]), .B0(n4428), .C0(n4429[32]), .D0(d1[68]), 
          .A1(d2[69]), .B1(n4428), .C1(n4429[33]), .D1(d1[69]), .CIN(n12228), 
          .COUT(n12229), .S0(d2_71__N_490[68]), .S1(d2_71__N_490[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1050_35.INIT0 = 16'h74b8;
    defparam add_1050_35.INIT1 = 16'h74b8;
    defparam add_1050_35.INJECT1_0 = "NO";
    defparam add_1050_35.INJECT1_1 = "NO";
    CCU2D add_1050_33 (.A0(d2[66]), .B0(n4428), .C0(n4429[30]), .D0(d1[66]), 
          .A1(d2[67]), .B1(n4428), .C1(n4429[31]), .D1(d1[67]), .CIN(n12227), 
          .COUT(n12228), .S0(d2_71__N_490[66]), .S1(d2_71__N_490[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1050_33.INIT0 = 16'h74b8;
    defparam add_1050_33.INIT1 = 16'h74b8;
    defparam add_1050_33.INJECT1_0 = "NO";
    defparam add_1050_33.INJECT1_1 = "NO";
    CCU2D add_1050_31 (.A0(d2[64]), .B0(n4428), .C0(n4429[28]), .D0(d1[64]), 
          .A1(d2[65]), .B1(n4428), .C1(n4429[29]), .D1(d1[65]), .CIN(n12226), 
          .COUT(n12227), .S0(d2_71__N_490[64]), .S1(d2_71__N_490[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1050_31.INIT0 = 16'h74b8;
    defparam add_1050_31.INIT1 = 16'h74b8;
    defparam add_1050_31.INJECT1_0 = "NO";
    defparam add_1050_31.INJECT1_1 = "NO";
    CCU2D add_1050_29 (.A0(d2[62]), .B0(n4428), .C0(n4429[26]), .D0(d1[62]), 
          .A1(d2[63]), .B1(n4428), .C1(n4429[27]), .D1(d1[63]), .CIN(n12225), 
          .COUT(n12226), .S0(d2_71__N_490[62]), .S1(d2_71__N_490[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1050_29.INIT0 = 16'h74b8;
    defparam add_1050_29.INIT1 = 16'h74b8;
    defparam add_1050_29.INJECT1_0 = "NO";
    defparam add_1050_29.INJECT1_1 = "NO";
    CCU2D add_1050_27 (.A0(d2[60]), .B0(n4428), .C0(n4429[24]), .D0(d1[60]), 
          .A1(d2[61]), .B1(n4428), .C1(n4429[25]), .D1(d1[61]), .CIN(n12224), 
          .COUT(n12225), .S0(d2_71__N_490[60]), .S1(d2_71__N_490[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1050_27.INIT0 = 16'h74b8;
    defparam add_1050_27.INIT1 = 16'h74b8;
    defparam add_1050_27.INJECT1_0 = "NO";
    defparam add_1050_27.INJECT1_1 = "NO";
    CCU2D add_1050_25 (.A0(d2[58]), .B0(n4428), .C0(n4429[22]), .D0(d1[58]), 
          .A1(d2[59]), .B1(n4428), .C1(n4429[23]), .D1(d1[59]), .CIN(n12223), 
          .COUT(n12224), .S0(d2_71__N_490[58]), .S1(d2_71__N_490[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1050_25.INIT0 = 16'h74b8;
    defparam add_1050_25.INIT1 = 16'h74b8;
    defparam add_1050_25.INJECT1_0 = "NO";
    defparam add_1050_25.INJECT1_1 = "NO";
    CCU2D add_1050_23 (.A0(d2[56]), .B0(n4428), .C0(n4429[20]), .D0(d1[56]), 
          .A1(d2[57]), .B1(n4428), .C1(n4429[21]), .D1(d1[57]), .CIN(n12222), 
          .COUT(n12223), .S0(d2_71__N_490[56]), .S1(d2_71__N_490[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1050_23.INIT0 = 16'h74b8;
    defparam add_1050_23.INIT1 = 16'h74b8;
    defparam add_1050_23.INJECT1_0 = "NO";
    defparam add_1050_23.INJECT1_1 = "NO";
    CCU2D add_1050_21 (.A0(d2[54]), .B0(n4428), .C0(n4429[18]), .D0(d1[54]), 
          .A1(d2[55]), .B1(n4428), .C1(n4429[19]), .D1(d1[55]), .CIN(n12221), 
          .COUT(n12222), .S0(d2_71__N_490[54]), .S1(d2_71__N_490[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1050_21.INIT0 = 16'h74b8;
    defparam add_1050_21.INIT1 = 16'h74b8;
    defparam add_1050_21.INJECT1_0 = "NO";
    defparam add_1050_21.INJECT1_1 = "NO";
    FD1S3IX count__i2 (.D(n375[2]), .CK(osc_clk), .CD(n8376), .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n375[3]), .CK(osc_clk), .CD(n8376), .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n375[4]), .CK(osc_clk), .CD(n8376), .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n375[5]), .CK(osc_clk), .CD(n8376), .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n375[6]), .CK(osc_clk), .CD(n8376), .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n375[7]), .CK(osc_clk), .CD(n8376), .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n375[8]), .CK(osc_clk), .CD(n8376), .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n375[9]), .CK(osc_clk), .CD(n8376), .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n375[10]), .CK(osc_clk), .CD(n8376), .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_15__N_1442[11]), .CK(osc_clk), .CD(d_clk_tmp_N_1831), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(n375[12]), .CK(osc_clk), .CD(n8376), .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(n375[13]), .CK(osc_clk), .CD(n8376), .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(n375[14]), .CK(osc_clk), .CD(n8376), .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(n375[15]), .CK(osc_clk), .CD(n8376), .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i15.GSR = "ENABLED";
    CCU2D add_1050_19 (.A0(d2[52]), .B0(n4428), .C0(n4429[16]), .D0(d1[52]), 
          .A1(d2[53]), .B1(n4428), .C1(n4429[17]), .D1(d1[53]), .CIN(n12220), 
          .COUT(n12221), .S0(d2_71__N_490[52]), .S1(d2_71__N_490[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1050_19.INIT0 = 16'h74b8;
    defparam add_1050_19.INIT1 = 16'h74b8;
    defparam add_1050_19.INJECT1_0 = "NO";
    defparam add_1050_19.INJECT1_1 = "NO";
    LUT4 i2849_2_lut (.A(n375[0]), .B(n31), .Z(count_15__N_1442[0])) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(86[13] 89[16])
    defparam i2849_2_lut.init = 16'hbbbb;
    LUT4 shift_right_31_i131_3_lut_4_lut_adj_42 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n61_adj_2521), .D(d10[59]), .Z(n131)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i131_3_lut_4_lut_adj_42.init = 16'hf960;
    CCU2D add_1050_17 (.A0(d2[50]), .B0(n4428), .C0(n4429[14]), .D0(d1[50]), 
          .A1(d2[51]), .B1(n4428), .C1(n4429[15]), .D1(d1[51]), .CIN(n12219), 
          .COUT(n12220), .S0(d2_71__N_490[50]), .S1(d2_71__N_490[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1050_17.INIT0 = 16'h74b8;
    defparam add_1050_17.INIT1 = 16'h74b8;
    defparam add_1050_17.INJECT1_0 = "NO";
    defparam add_1050_17.INJECT1_1 = "NO";
    CCU2D add_1050_15 (.A0(d2[48]), .B0(n4428), .C0(n4429[12]), .D0(d1[48]), 
          .A1(d2[49]), .B1(n4428), .C1(n4429[13]), .D1(d1[49]), .CIN(n12218), 
          .COUT(n12219), .S0(d2_71__N_490[48]), .S1(d2_71__N_490[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1050_15.INIT0 = 16'h74b8;
    defparam add_1050_15.INIT1 = 16'h74b8;
    defparam add_1050_15.INJECT1_0 = "NO";
    defparam add_1050_15.INJECT1_1 = "NO";
    CCU2D add_1050_13 (.A0(d2[46]), .B0(n4428), .C0(n4429[10]), .D0(d1[46]), 
          .A1(d2[47]), .B1(n4428), .C1(n4429[11]), .D1(d1[47]), .CIN(n12217), 
          .COUT(n12218), .S0(d2_71__N_490[46]), .S1(d2_71__N_490[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1050_13.INIT0 = 16'h74b8;
    defparam add_1050_13.INIT1 = 16'h74b8;
    defparam add_1050_13.INJECT1_0 = "NO";
    defparam add_1050_13.INJECT1_1 = "NO";
    CCU2D add_1050_11 (.A0(d2[44]), .B0(n4428), .C0(n4429[8]), .D0(d1[44]), 
          .A1(d2[45]), .B1(n4428), .C1(n4429[9]), .D1(d1[45]), .CIN(n12216), 
          .COUT(n12217), .S0(d2_71__N_490[44]), .S1(d2_71__N_490[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1050_11.INIT0 = 16'h74b8;
    defparam add_1050_11.INIT1 = 16'h74b8;
    defparam add_1050_11.INJECT1_0 = "NO";
    defparam add_1050_11.INJECT1_1 = "NO";
    CCU2D add_1050_9 (.A0(d2[42]), .B0(n4428), .C0(n4429[6]), .D0(d1[42]), 
          .A1(d2[43]), .B1(n4428), .C1(n4429[7]), .D1(d1[43]), .CIN(n12215), 
          .COUT(n12216), .S0(d2_71__N_490[42]), .S1(d2_71__N_490[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1050_9.INIT0 = 16'h74b8;
    defparam add_1050_9.INIT1 = 16'h74b8;
    defparam add_1050_9.INJECT1_0 = "NO";
    defparam add_1050_9.INJECT1_1 = "NO";
    CCU2D add_1050_7 (.A0(d2[40]), .B0(n4428), .C0(n4429[4]), .D0(d1[40]), 
          .A1(d2[41]), .B1(n4428), .C1(n4429[5]), .D1(d1[41]), .CIN(n12214), 
          .COUT(n12215), .S0(d2_71__N_490[40]), .S1(d2_71__N_490[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1050_7.INIT0 = 16'h74b8;
    defparam add_1050_7.INIT1 = 16'h74b8;
    defparam add_1050_7.INJECT1_0 = "NO";
    defparam add_1050_7.INJECT1_1 = "NO";
    CCU2D add_1050_5 (.A0(d2[38]), .B0(n4428), .C0(n4429[2]), .D0(d1[38]), 
          .A1(d2[39]), .B1(n4428), .C1(n4429[3]), .D1(d1[39]), .CIN(n12213), 
          .COUT(n12214), .S0(d2_71__N_490[38]), .S1(d2_71__N_490[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1050_5.INIT0 = 16'h74b8;
    defparam add_1050_5.INIT1 = 16'h74b8;
    defparam add_1050_5.INJECT1_0 = "NO";
    defparam add_1050_5.INJECT1_1 = "NO";
    CCU2D add_1050_3 (.A0(d2[36]), .B0(n4428), .C0(n4429[0]), .D0(d1[36]), 
          .A1(d2[37]), .B1(n4428), .C1(n4429[1]), .D1(d1[37]), .CIN(n12212), 
          .COUT(n12213), .S0(d2_71__N_490[36]), .S1(d2_71__N_490[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1050_3.INIT0 = 16'h74b8;
    defparam add_1050_3.INIT1 = 16'h74b8;
    defparam add_1050_3.INJECT1_0 = "NO";
    defparam add_1050_3.INJECT1_1 = "NO";
    CCU2D add_1050_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n4428), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n12212));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1050_1.INIT0 = 16'hF000;
    defparam add_1050_1.INIT1 = 16'h0555;
    defparam add_1050_1.INJECT1_0 = "NO";
    defparam add_1050_1.INJECT1_1 = "NO";
    CCU2D add_1095_3 (.A0(d_d8[36]), .B0(n5796), .C0(n5797[0]), .D0(d8[36]), 
          .A1(d_d8[37]), .B1(n5796), .C1(n5797[1]), .D1(d8[37]), .CIN(n11844), 
          .COUT(n11845), .S0(d9_71__N_1675[36]), .S1(d9_71__N_1675[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1095_3.INIT0 = 16'hb874;
    defparam add_1095_3.INIT1 = 16'hb874;
    defparam add_1095_3.INJECT1_0 = "NO";
    defparam add_1095_3.INJECT1_1 = "NO";
    CCU2D add_1099_27 (.A0(d9[61]), .B0(d_d9[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[62]), .B1(d_d9[62]), .C1(GND_net), .D1(GND_net), .CIN(n11835), 
          .COUT(n11836), .S0(n5949[25]), .S1(n5949[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1099_27.INIT0 = 16'h5999;
    defparam add_1099_27.INIT1 = 16'h5999;
    defparam add_1099_27.INJECT1_0 = "NO";
    defparam add_1099_27.INJECT1_1 = "NO";
    CCU2D add_1099_25 (.A0(d9[59]), .B0(d_d9[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[60]), .B1(d_d9[60]), .C1(GND_net), .D1(GND_net), .CIN(n11834), 
          .COUT(n11835), .S0(n5949[23]), .S1(n5949[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1099_25.INIT0 = 16'h5999;
    defparam add_1099_25.INIT1 = 16'h5999;
    defparam add_1099_25.INJECT1_0 = "NO";
    defparam add_1099_25.INJECT1_1 = "NO";
    CCU2D add_1099_23 (.A0(d9[57]), .B0(d_d9[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[58]), .B1(d_d9[58]), .C1(GND_net), .D1(GND_net), .CIN(n11833), 
          .COUT(n11834), .S0(n5949[21]), .S1(n5949[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1099_23.INIT0 = 16'h5999;
    defparam add_1099_23.INIT1 = 16'h5999;
    defparam add_1099_23.INJECT1_0 = "NO";
    defparam add_1099_23.INJECT1_1 = "NO";
    CCU2D add_1054_36 (.A0(d2[70]), .B0(d3[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[71]), .B1(d3[71]), .C1(GND_net), .D1(GND_net), .CIN(n12207), 
          .S0(n4581[34]), .S1(n4581[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1054_36.INIT0 = 16'h5666;
    defparam add_1054_36.INIT1 = 16'h5666;
    defparam add_1054_36.INJECT1_0 = "NO";
    defparam add_1054_36.INJECT1_1 = "NO";
    CCU2D add_1054_34 (.A0(d2[68]), .B0(d3[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[69]), .B1(d3[69]), .C1(GND_net), .D1(GND_net), .CIN(n12206), 
          .COUT(n12207), .S0(n4581[32]), .S1(n4581[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1054_34.INIT0 = 16'h5666;
    defparam add_1054_34.INIT1 = 16'h5666;
    defparam add_1054_34.INJECT1_0 = "NO";
    defparam add_1054_34.INJECT1_1 = "NO";
    CCU2D add_1129_37 (.A0(d7[71]), .B0(d_d7[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11427), 
          .S0(n6861[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1129_37.INIT0 = 16'h5999;
    defparam add_1129_37.INIT1 = 16'h0000;
    defparam add_1129_37.INJECT1_0 = "NO";
    defparam add_1129_37.INJECT1_1 = "NO";
    CCU2D add_1129_35 (.A0(d7[69]), .B0(d_d7[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[70]), .B1(d_d7[70]), .C1(GND_net), .D1(GND_net), .CIN(n11426), 
          .COUT(n11427), .S0(n6861[33]), .S1(n6861[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1129_35.INIT0 = 16'h5999;
    defparam add_1129_35.INIT1 = 16'h5999;
    defparam add_1129_35.INJECT1_0 = "NO";
    defparam add_1129_35.INJECT1_1 = "NO";
    CCU2D add_1129_33 (.A0(d7[67]), .B0(d_d7[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[68]), .B1(d_d7[68]), .C1(GND_net), .D1(GND_net), .CIN(n11425), 
          .COUT(n11426), .S0(n6861[31]), .S1(n6861[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1129_33.INIT0 = 16'h5999;
    defparam add_1129_33.INIT1 = 16'h5999;
    defparam add_1129_33.INJECT1_0 = "NO";
    defparam add_1129_33.INJECT1_1 = "NO";
    CCU2D add_1129_31 (.A0(d7[65]), .B0(d_d7[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[66]), .B1(d_d7[66]), .C1(GND_net), .D1(GND_net), .CIN(n11424), 
          .COUT(n11425), .S0(n6861[29]), .S1(n6861[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1129_31.INIT0 = 16'h5999;
    defparam add_1129_31.INIT1 = 16'h5999;
    defparam add_1129_31.INJECT1_0 = "NO";
    defparam add_1129_31.INJECT1_1 = "NO";
    CCU2D add_1129_29 (.A0(d7[63]), .B0(d_d7[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[64]), .B1(d_d7[64]), .C1(GND_net), .D1(GND_net), .CIN(n11423), 
          .COUT(n11424), .S0(n6861[27]), .S1(n6861[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1129_29.INIT0 = 16'h5999;
    defparam add_1129_29.INIT1 = 16'h5999;
    defparam add_1129_29.INJECT1_0 = "NO";
    defparam add_1129_29.INJECT1_1 = "NO";
    CCU2D add_1129_27 (.A0(d7[61]), .B0(d_d7[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[62]), .B1(d_d7[62]), .C1(GND_net), .D1(GND_net), .CIN(n11422), 
          .COUT(n11423), .S0(n6861[25]), .S1(n6861[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1129_27.INIT0 = 16'h5999;
    defparam add_1129_27.INIT1 = 16'h5999;
    defparam add_1129_27.INJECT1_0 = "NO";
    defparam add_1129_27.INJECT1_1 = "NO";
    CCU2D add_1129_25 (.A0(d7[59]), .B0(d_d7[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[60]), .B1(d_d7[60]), .C1(GND_net), .D1(GND_net), .CIN(n11421), 
          .COUT(n11422), .S0(n6861[23]), .S1(n6861[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1129_25.INIT0 = 16'h5999;
    defparam add_1129_25.INIT1 = 16'h5999;
    defparam add_1129_25.INJECT1_0 = "NO";
    defparam add_1129_25.INJECT1_1 = "NO";
    CCU2D add_1129_23 (.A0(d7[57]), .B0(d_d7[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[58]), .B1(d_d7[58]), .C1(GND_net), .D1(GND_net), .CIN(n11420), 
          .COUT(n11421), .S0(n6861[21]), .S1(n6861[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1129_23.INIT0 = 16'h5999;
    defparam add_1129_23.INIT1 = 16'h5999;
    defparam add_1129_23.INJECT1_0 = "NO";
    defparam add_1129_23.INJECT1_1 = "NO";
    CCU2D add_1129_21 (.A0(d7[55]), .B0(d_d7[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[56]), .B1(d_d7[56]), .C1(GND_net), .D1(GND_net), .CIN(n11419), 
          .COUT(n11420), .S0(n6861[19]), .S1(n6861[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1129_21.INIT0 = 16'h5999;
    defparam add_1129_21.INIT1 = 16'h5999;
    defparam add_1129_21.INJECT1_0 = "NO";
    defparam add_1129_21.INJECT1_1 = "NO";
    CCU2D add_1129_19 (.A0(d7[53]), .B0(d_d7[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[54]), .B1(d_d7[54]), .C1(GND_net), .D1(GND_net), .CIN(n11418), 
          .COUT(n11419), .S0(n6861[17]), .S1(n6861[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1129_19.INIT0 = 16'h5999;
    defparam add_1129_19.INIT1 = 16'h5999;
    defparam add_1129_19.INJECT1_0 = "NO";
    defparam add_1129_19.INJECT1_1 = "NO";
    CCU2D add_1129_17 (.A0(d7[51]), .B0(d_d7[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[52]), .B1(d_d7[52]), .C1(GND_net), .D1(GND_net), .CIN(n11417), 
          .COUT(n11418), .S0(n6861[15]), .S1(n6861[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1129_17.INIT0 = 16'h5999;
    defparam add_1129_17.INIT1 = 16'h5999;
    defparam add_1129_17.INJECT1_0 = "NO";
    defparam add_1129_17.INJECT1_1 = "NO";
    CCU2D add_1129_15 (.A0(d7[49]), .B0(d_d7[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[50]), .B1(d_d7[50]), .C1(GND_net), .D1(GND_net), .CIN(n11416), 
          .COUT(n11417), .S0(n6861[13]), .S1(n6861[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1129_15.INIT0 = 16'h5999;
    defparam add_1129_15.INIT1 = 16'h5999;
    defparam add_1129_15.INJECT1_0 = "NO";
    defparam add_1129_15.INJECT1_1 = "NO";
    CCU2D add_1129_13 (.A0(d7[47]), .B0(d_d7[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[48]), .B1(d_d7[48]), .C1(GND_net), .D1(GND_net), .CIN(n11415), 
          .COUT(n11416), .S0(n6861[11]), .S1(n6861[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1129_13.INIT0 = 16'h5999;
    defparam add_1129_13.INIT1 = 16'h5999;
    defparam add_1129_13.INJECT1_0 = "NO";
    defparam add_1129_13.INJECT1_1 = "NO";
    CCU2D add_1129_11 (.A0(d7[45]), .B0(d_d7[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[46]), .B1(d_d7[46]), .C1(GND_net), .D1(GND_net), .CIN(n11414), 
          .COUT(n11415), .S0(n6861[9]), .S1(n6861[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1129_11.INIT0 = 16'h5999;
    defparam add_1129_11.INIT1 = 16'h5999;
    defparam add_1129_11.INJECT1_0 = "NO";
    defparam add_1129_11.INJECT1_1 = "NO";
    CCU2D add_1129_9 (.A0(d7[43]), .B0(d_d7[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[44]), .B1(d_d7[44]), .C1(GND_net), .D1(GND_net), .CIN(n11413), 
          .COUT(n11414), .S0(n6861[7]), .S1(n6861[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1129_9.INIT0 = 16'h5999;
    defparam add_1129_9.INIT1 = 16'h5999;
    defparam add_1129_9.INJECT1_0 = "NO";
    defparam add_1129_9.INJECT1_1 = "NO";
    CCU2D add_1129_7 (.A0(d7[41]), .B0(d_d7[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[42]), .B1(d_d7[42]), .C1(GND_net), .D1(GND_net), .CIN(n11412), 
          .COUT(n11413), .S0(n6861[5]), .S1(n6861[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1129_7.INIT0 = 16'h5999;
    defparam add_1129_7.INIT1 = 16'h5999;
    defparam add_1129_7.INJECT1_0 = "NO";
    defparam add_1129_7.INJECT1_1 = "NO";
    CCU2D add_1129_5 (.A0(d7[39]), .B0(d_d7[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[40]), .B1(d_d7[40]), .C1(GND_net), .D1(GND_net), .CIN(n11411), 
          .COUT(n11412), .S0(n6861[3]), .S1(n6861[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1129_5.INIT0 = 16'h5999;
    defparam add_1129_5.INIT1 = 16'h5999;
    defparam add_1129_5.INJECT1_0 = "NO";
    defparam add_1129_5.INJECT1_1 = "NO";
    CCU2D add_1129_3 (.A0(d7[37]), .B0(d_d7[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[38]), .B1(d_d7[38]), .C1(GND_net), .D1(GND_net), .CIN(n11410), 
          .COUT(n11411), .S0(n6861[1]), .S1(n6861[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1129_3.INIT0 = 16'h5999;
    defparam add_1129_3.INIT1 = 16'h5999;
    defparam add_1129_3.INJECT1_0 = "NO";
    defparam add_1129_3.INJECT1_1 = "NO";
    CCU2D add_1129_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d7[36]), .B1(d_d7[36]), .C1(GND_net), .D1(GND_net), .COUT(n11410), 
          .S1(n6861[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1129_1.INIT0 = 16'hF000;
    defparam add_1129_1.INIT1 = 16'h5999;
    defparam add_1129_1.INJECT1_0 = "NO";
    defparam add_1129_1.INJECT1_1 = "NO";
    CCU2D add_1130_37 (.A0(d_d7[70]), .B0(n6860), .C0(n6861[34]), .D0(d7[70]), 
          .A1(d_d7[71]), .B1(n6860), .C1(n6861[35]), .D1(d7[71]), .CIN(n11408), 
          .S0(d8_71__N_1603[70]), .S1(d8_71__N_1603[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1130_37.INIT0 = 16'hb874;
    defparam add_1130_37.INIT1 = 16'hb874;
    defparam add_1130_37.INJECT1_0 = "NO";
    defparam add_1130_37.INJECT1_1 = "NO";
    CCU2D add_1130_35 (.A0(d_d7[68]), .B0(n6860), .C0(n6861[32]), .D0(d7[68]), 
          .A1(d_d7[69]), .B1(n6860), .C1(n6861[33]), .D1(d7[69]), .CIN(n11407), 
          .COUT(n11408), .S0(d8_71__N_1603[68]), .S1(d8_71__N_1603[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1130_35.INIT0 = 16'hb874;
    defparam add_1130_35.INIT1 = 16'hb874;
    defparam add_1130_35.INJECT1_0 = "NO";
    defparam add_1130_35.INJECT1_1 = "NO";
    CCU2D add_1130_33 (.A0(d_d7[66]), .B0(n6860), .C0(n6861[30]), .D0(d7[66]), 
          .A1(d_d7[67]), .B1(n6860), .C1(n6861[31]), .D1(d7[67]), .CIN(n11406), 
          .COUT(n11407), .S0(d8_71__N_1603[66]), .S1(d8_71__N_1603[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1130_33.INIT0 = 16'hb874;
    defparam add_1130_33.INIT1 = 16'hb874;
    defparam add_1130_33.INJECT1_0 = "NO";
    defparam add_1130_33.INJECT1_1 = "NO";
    CCU2D add_1130_31 (.A0(d_d7[64]), .B0(n6860), .C0(n6861[28]), .D0(d7[64]), 
          .A1(d_d7[65]), .B1(n6860), .C1(n6861[29]), .D1(d7[65]), .CIN(n11405), 
          .COUT(n11406), .S0(d8_71__N_1603[64]), .S1(d8_71__N_1603[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1130_31.INIT0 = 16'hb874;
    defparam add_1130_31.INIT1 = 16'hb874;
    defparam add_1130_31.INJECT1_0 = "NO";
    defparam add_1130_31.INJECT1_1 = "NO";
    CCU2D add_1130_29 (.A0(d_d7[62]), .B0(n6860), .C0(n6861[26]), .D0(d7[62]), 
          .A1(d_d7[63]), .B1(n6860), .C1(n6861[27]), .D1(d7[63]), .CIN(n11404), 
          .COUT(n11405), .S0(d8_71__N_1603[62]), .S1(d8_71__N_1603[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1130_29.INIT0 = 16'hb874;
    defparam add_1130_29.INIT1 = 16'hb874;
    defparam add_1130_29.INJECT1_0 = "NO";
    defparam add_1130_29.INJECT1_1 = "NO";
    CCU2D add_1130_27 (.A0(d_d7[60]), .B0(n6860), .C0(n6861[24]), .D0(d7[60]), 
          .A1(d_d7[61]), .B1(n6860), .C1(n6861[25]), .D1(d7[61]), .CIN(n11403), 
          .COUT(n11404), .S0(d8_71__N_1603[60]), .S1(d8_71__N_1603[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1130_27.INIT0 = 16'hb874;
    defparam add_1130_27.INIT1 = 16'hb874;
    defparam add_1130_27.INJECT1_0 = "NO";
    defparam add_1130_27.INJECT1_1 = "NO";
    CCU2D add_1130_25 (.A0(d_d7[58]), .B0(n6860), .C0(n6861[22]), .D0(d7[58]), 
          .A1(d_d7[59]), .B1(n6860), .C1(n6861[23]), .D1(d7[59]), .CIN(n11402), 
          .COUT(n11403), .S0(d8_71__N_1603[58]), .S1(d8_71__N_1603[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1130_25.INIT0 = 16'hb874;
    defparam add_1130_25.INIT1 = 16'hb874;
    defparam add_1130_25.INJECT1_0 = "NO";
    defparam add_1130_25.INJECT1_1 = "NO";
    CCU2D add_1130_23 (.A0(d_d7[56]), .B0(n6860), .C0(n6861[20]), .D0(d7[56]), 
          .A1(d_d7[57]), .B1(n6860), .C1(n6861[21]), .D1(d7[57]), .CIN(n11401), 
          .COUT(n11402), .S0(d8_71__N_1603[56]), .S1(d8_71__N_1603[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1130_23.INIT0 = 16'hb874;
    defparam add_1130_23.INIT1 = 16'hb874;
    defparam add_1130_23.INJECT1_0 = "NO";
    defparam add_1130_23.INJECT1_1 = "NO";
    CCU2D add_1130_21 (.A0(d_d7[54]), .B0(n6860), .C0(n6861[18]), .D0(d7[54]), 
          .A1(d_d7[55]), .B1(n6860), .C1(n6861[19]), .D1(d7[55]), .CIN(n11400), 
          .COUT(n11401), .S0(d8_71__N_1603[54]), .S1(d8_71__N_1603[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1130_21.INIT0 = 16'hb874;
    defparam add_1130_21.INIT1 = 16'hb874;
    defparam add_1130_21.INJECT1_0 = "NO";
    defparam add_1130_21.INJECT1_1 = "NO";
    CCU2D add_1130_19 (.A0(d_d7[52]), .B0(n6860), .C0(n6861[16]), .D0(d7[52]), 
          .A1(d_d7[53]), .B1(n6860), .C1(n6861[17]), .D1(d7[53]), .CIN(n11399), 
          .COUT(n11400), .S0(d8_71__N_1603[52]), .S1(d8_71__N_1603[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1130_19.INIT0 = 16'hb874;
    defparam add_1130_19.INIT1 = 16'hb874;
    defparam add_1130_19.INJECT1_0 = "NO";
    defparam add_1130_19.INJECT1_1 = "NO";
    CCU2D add_1130_17 (.A0(d_d7[50]), .B0(n6860), .C0(n6861[14]), .D0(d7[50]), 
          .A1(d_d7[51]), .B1(n6860), .C1(n6861[15]), .D1(d7[51]), .CIN(n11398), 
          .COUT(n11399), .S0(d8_71__N_1603[50]), .S1(d8_71__N_1603[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1130_17.INIT0 = 16'hb874;
    defparam add_1130_17.INIT1 = 16'hb874;
    defparam add_1130_17.INJECT1_0 = "NO";
    defparam add_1130_17.INJECT1_1 = "NO";
    CCU2D add_1130_15 (.A0(d_d7[48]), .B0(n6860), .C0(n6861[12]), .D0(d7[48]), 
          .A1(d_d7[49]), .B1(n6860), .C1(n6861[13]), .D1(d7[49]), .CIN(n11397), 
          .COUT(n11398), .S0(d8_71__N_1603[48]), .S1(d8_71__N_1603[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1130_15.INIT0 = 16'hb874;
    defparam add_1130_15.INIT1 = 16'hb874;
    defparam add_1130_15.INJECT1_0 = "NO";
    defparam add_1130_15.INJECT1_1 = "NO";
    CCU2D add_1130_13 (.A0(d_d7[46]), .B0(n6860), .C0(n6861[10]), .D0(d7[46]), 
          .A1(d_d7[47]), .B1(n6860), .C1(n6861[11]), .D1(d7[47]), .CIN(n11396), 
          .COUT(n11397), .S0(d8_71__N_1603[46]), .S1(d8_71__N_1603[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1130_13.INIT0 = 16'hb874;
    defparam add_1130_13.INIT1 = 16'hb874;
    defparam add_1130_13.INJECT1_0 = "NO";
    defparam add_1130_13.INJECT1_1 = "NO";
    CCU2D add_1130_11 (.A0(d_d7[44]), .B0(n6860), .C0(n6861[8]), .D0(d7[44]), 
          .A1(d_d7[45]), .B1(n6860), .C1(n6861[9]), .D1(d7[45]), .CIN(n11395), 
          .COUT(n11396), .S0(d8_71__N_1603[44]), .S1(d8_71__N_1603[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1130_11.INIT0 = 16'hb874;
    defparam add_1130_11.INIT1 = 16'hb874;
    defparam add_1130_11.INJECT1_0 = "NO";
    defparam add_1130_11.INJECT1_1 = "NO";
    CCU2D add_1130_9 (.A0(d_d7[42]), .B0(n6860), .C0(n6861[6]), .D0(d7[42]), 
          .A1(d_d7[43]), .B1(n6860), .C1(n6861[7]), .D1(d7[43]), .CIN(n11394), 
          .COUT(n11395), .S0(d8_71__N_1603[42]), .S1(d8_71__N_1603[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1130_9.INIT0 = 16'hb874;
    defparam add_1130_9.INIT1 = 16'hb874;
    defparam add_1130_9.INJECT1_0 = "NO";
    defparam add_1130_9.INJECT1_1 = "NO";
    CCU2D add_1130_7 (.A0(d_d7[40]), .B0(n6860), .C0(n6861[4]), .D0(d7[40]), 
          .A1(d_d7[41]), .B1(n6860), .C1(n6861[5]), .D1(d7[41]), .CIN(n11393), 
          .COUT(n11394), .S0(d8_71__N_1603[40]), .S1(d8_71__N_1603[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1130_7.INIT0 = 16'hb874;
    defparam add_1130_7.INIT1 = 16'hb874;
    defparam add_1130_7.INJECT1_0 = "NO";
    defparam add_1130_7.INJECT1_1 = "NO";
    CCU2D add_1130_5 (.A0(d_d7[38]), .B0(n6860), .C0(n6861[2]), .D0(d7[38]), 
          .A1(d_d7[39]), .B1(n6860), .C1(n6861[3]), .D1(d7[39]), .CIN(n11392), 
          .COUT(n11393), .S0(d8_71__N_1603[38]), .S1(d8_71__N_1603[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1130_5.INIT0 = 16'hb874;
    defparam add_1130_5.INIT1 = 16'hb874;
    defparam add_1130_5.INJECT1_0 = "NO";
    defparam add_1130_5.INJECT1_1 = "NO";
    CCU2D add_1130_3 (.A0(d_d7[36]), .B0(n6860), .C0(n6861[0]), .D0(d7[36]), 
          .A1(d_d7[37]), .B1(n6860), .C1(n6861[1]), .D1(d7[37]), .CIN(n11391), 
          .COUT(n11392), .S0(d8_71__N_1603[36]), .S1(d8_71__N_1603[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1130_3.INIT0 = 16'hb874;
    defparam add_1130_3.INIT1 = 16'hb874;
    defparam add_1130_3.INJECT1_0 = "NO";
    defparam add_1130_3.INJECT1_1 = "NO";
    CCU2D add_1130_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n6860), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11391));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1130_1.INIT0 = 16'hF000;
    defparam add_1130_1.INIT1 = 16'h0555;
    defparam add_1130_1.INJECT1_0 = "NO";
    defparam add_1130_1.INJECT1_1 = "NO";
    CCU2D add_1134_37 (.A0(d6[71]), .B0(d_d6[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11387), 
          .S0(n7013[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1134_37.INIT0 = 16'h5999;
    defparam add_1134_37.INIT1 = 16'h0000;
    defparam add_1134_37.INJECT1_0 = "NO";
    defparam add_1134_37.INJECT1_1 = "NO";
    CCU2D add_1134_35 (.A0(d6[69]), .B0(d_d6[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[70]), .B1(d_d6[70]), .C1(GND_net), .D1(GND_net), .CIN(n11386), 
          .COUT(n11387), .S0(n7013[33]), .S1(n7013[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1134_35.INIT0 = 16'h5999;
    defparam add_1134_35.INIT1 = 16'h5999;
    defparam add_1134_35.INJECT1_0 = "NO";
    defparam add_1134_35.INJECT1_1 = "NO";
    CCU2D add_1134_33 (.A0(d6[67]), .B0(d_d6[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[68]), .B1(d_d6[68]), .C1(GND_net), .D1(GND_net), .CIN(n11385), 
          .COUT(n11386), .S0(n7013[31]), .S1(n7013[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1134_33.INIT0 = 16'h5999;
    defparam add_1134_33.INIT1 = 16'h5999;
    defparam add_1134_33.INJECT1_0 = "NO";
    defparam add_1134_33.INJECT1_1 = "NO";
    CCU2D add_1134_31 (.A0(d6[65]), .B0(d_d6[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[66]), .B1(d_d6[66]), .C1(GND_net), .D1(GND_net), .CIN(n11384), 
          .COUT(n11385), .S0(n7013[29]), .S1(n7013[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1134_31.INIT0 = 16'h5999;
    defparam add_1134_31.INIT1 = 16'h5999;
    defparam add_1134_31.INJECT1_0 = "NO";
    defparam add_1134_31.INJECT1_1 = "NO";
    CCU2D add_1134_29 (.A0(d6[63]), .B0(d_d6[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[64]), .B1(d_d6[64]), .C1(GND_net), .D1(GND_net), .CIN(n11383), 
          .COUT(n11384), .S0(n7013[27]), .S1(n7013[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1134_29.INIT0 = 16'h5999;
    defparam add_1134_29.INIT1 = 16'h5999;
    defparam add_1134_29.INJECT1_0 = "NO";
    defparam add_1134_29.INJECT1_1 = "NO";
    CCU2D add_1134_27 (.A0(d6[61]), .B0(d_d6[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[62]), .B1(d_d6[62]), .C1(GND_net), .D1(GND_net), .CIN(n11382), 
          .COUT(n11383), .S0(n7013[25]), .S1(n7013[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1134_27.INIT0 = 16'h5999;
    defparam add_1134_27.INIT1 = 16'h5999;
    defparam add_1134_27.INJECT1_0 = "NO";
    defparam add_1134_27.INJECT1_1 = "NO";
    CCU2D add_1134_25 (.A0(d6[59]), .B0(d_d6[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[60]), .B1(d_d6[60]), .C1(GND_net), .D1(GND_net), .CIN(n11381), 
          .COUT(n11382), .S0(n7013[23]), .S1(n7013[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1134_25.INIT0 = 16'h5999;
    defparam add_1134_25.INIT1 = 16'h5999;
    defparam add_1134_25.INJECT1_0 = "NO";
    defparam add_1134_25.INJECT1_1 = "NO";
    CCU2D add_1134_23 (.A0(d6[57]), .B0(d_d6[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[58]), .B1(d_d6[58]), .C1(GND_net), .D1(GND_net), .CIN(n11380), 
          .COUT(n11381), .S0(n7013[21]), .S1(n7013[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1134_23.INIT0 = 16'h5999;
    defparam add_1134_23.INIT1 = 16'h5999;
    defparam add_1134_23.INJECT1_0 = "NO";
    defparam add_1134_23.INJECT1_1 = "NO";
    CCU2D add_1134_21 (.A0(d6[55]), .B0(d_d6[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[56]), .B1(d_d6[56]), .C1(GND_net), .D1(GND_net), .CIN(n11379), 
          .COUT(n11380), .S0(n7013[19]), .S1(n7013[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1134_21.INIT0 = 16'h5999;
    defparam add_1134_21.INIT1 = 16'h5999;
    defparam add_1134_21.INJECT1_0 = "NO";
    defparam add_1134_21.INJECT1_1 = "NO";
    CCU2D add_1134_19 (.A0(d6[53]), .B0(d_d6[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[54]), .B1(d_d6[54]), .C1(GND_net), .D1(GND_net), .CIN(n11378), 
          .COUT(n11379), .S0(n7013[17]), .S1(n7013[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1134_19.INIT0 = 16'h5999;
    defparam add_1134_19.INIT1 = 16'h5999;
    defparam add_1134_19.INJECT1_0 = "NO";
    defparam add_1134_19.INJECT1_1 = "NO";
    CCU2D add_1134_17 (.A0(d6[51]), .B0(d_d6[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[52]), .B1(d_d6[52]), .C1(GND_net), .D1(GND_net), .CIN(n11377), 
          .COUT(n11378), .S0(n7013[15]), .S1(n7013[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1134_17.INIT0 = 16'h5999;
    defparam add_1134_17.INIT1 = 16'h5999;
    defparam add_1134_17.INJECT1_0 = "NO";
    defparam add_1134_17.INJECT1_1 = "NO";
    CCU2D add_1134_15 (.A0(d6[49]), .B0(d_d6[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[50]), .B1(d_d6[50]), .C1(GND_net), .D1(GND_net), .CIN(n11376), 
          .COUT(n11377), .S0(n7013[13]), .S1(n7013[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1134_15.INIT0 = 16'h5999;
    defparam add_1134_15.INIT1 = 16'h5999;
    defparam add_1134_15.INJECT1_0 = "NO";
    defparam add_1134_15.INJECT1_1 = "NO";
    CCU2D add_1134_13 (.A0(d6[47]), .B0(d_d6[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[48]), .B1(d_d6[48]), .C1(GND_net), .D1(GND_net), .CIN(n11375), 
          .COUT(n11376), .S0(n7013[11]), .S1(n7013[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1134_13.INIT0 = 16'h5999;
    defparam add_1134_13.INIT1 = 16'h5999;
    defparam add_1134_13.INJECT1_0 = "NO";
    defparam add_1134_13.INJECT1_1 = "NO";
    CCU2D add_1134_11 (.A0(d6[45]), .B0(d_d6[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[46]), .B1(d_d6[46]), .C1(GND_net), .D1(GND_net), .CIN(n11374), 
          .COUT(n11375), .S0(n7013[9]), .S1(n7013[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1134_11.INIT0 = 16'h5999;
    defparam add_1134_11.INIT1 = 16'h5999;
    defparam add_1134_11.INJECT1_0 = "NO";
    defparam add_1134_11.INJECT1_1 = "NO";
    CCU2D add_1134_9 (.A0(d6[43]), .B0(d_d6[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[44]), .B1(d_d6[44]), .C1(GND_net), .D1(GND_net), .CIN(n11373), 
          .COUT(n11374), .S0(n7013[7]), .S1(n7013[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1134_9.INIT0 = 16'h5999;
    defparam add_1134_9.INIT1 = 16'h5999;
    defparam add_1134_9.INJECT1_0 = "NO";
    defparam add_1134_9.INJECT1_1 = "NO";
    CCU2D add_1134_7 (.A0(d6[41]), .B0(d_d6[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[42]), .B1(d_d6[42]), .C1(GND_net), .D1(GND_net), .CIN(n11372), 
          .COUT(n11373), .S0(n7013[5]), .S1(n7013[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1134_7.INIT0 = 16'h5999;
    defparam add_1134_7.INIT1 = 16'h5999;
    defparam add_1134_7.INJECT1_0 = "NO";
    defparam add_1134_7.INJECT1_1 = "NO";
    CCU2D add_1134_5 (.A0(d6[39]), .B0(d_d6[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[40]), .B1(d_d6[40]), .C1(GND_net), .D1(GND_net), .CIN(n11371), 
          .COUT(n11372), .S0(n7013[3]), .S1(n7013[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1134_5.INIT0 = 16'h5999;
    defparam add_1134_5.INIT1 = 16'h5999;
    defparam add_1134_5.INJECT1_0 = "NO";
    defparam add_1134_5.INJECT1_1 = "NO";
    CCU2D add_1134_3 (.A0(d6[37]), .B0(d_d6[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[38]), .B1(d_d6[38]), .C1(GND_net), .D1(GND_net), .CIN(n11370), 
          .COUT(n11371), .S0(n7013[1]), .S1(n7013[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1134_3.INIT0 = 16'h5999;
    defparam add_1134_3.INIT1 = 16'h5999;
    defparam add_1134_3.INJECT1_0 = "NO";
    defparam add_1134_3.INJECT1_1 = "NO";
    CCU2D add_1134_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d6[36]), .B1(d_d6[36]), .C1(GND_net), .D1(GND_net), .COUT(n11370), 
          .S1(n7013[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1134_1.INIT0 = 16'hF000;
    defparam add_1134_1.INIT1 = 16'h5999;
    defparam add_1134_1.INJECT1_0 = "NO";
    defparam add_1134_1.INJECT1_1 = "NO";
    CCU2D add_1135_37 (.A0(d_d6[70]), .B0(n7012), .C0(n7013[34]), .D0(d6[70]), 
          .A1(d_d6[71]), .B1(n7012), .C1(n7013[35]), .D1(d6[71]), .CIN(n11368), 
          .S0(d7_71__N_1531[70]), .S1(d7_71__N_1531[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1135_37.INIT0 = 16'hb874;
    defparam add_1135_37.INIT1 = 16'hb874;
    defparam add_1135_37.INJECT1_0 = "NO";
    defparam add_1135_37.INJECT1_1 = "NO";
    CCU2D add_1135_35 (.A0(d_d6[68]), .B0(n7012), .C0(n7013[32]), .D0(d6[68]), 
          .A1(d_d6[69]), .B1(n7012), .C1(n7013[33]), .D1(d6[69]), .CIN(n11367), 
          .COUT(n11368), .S0(d7_71__N_1531[68]), .S1(d7_71__N_1531[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1135_35.INIT0 = 16'hb874;
    defparam add_1135_35.INIT1 = 16'hb874;
    defparam add_1135_35.INJECT1_0 = "NO";
    defparam add_1135_35.INJECT1_1 = "NO";
    CCU2D add_1135_33 (.A0(d_d6[66]), .B0(n7012), .C0(n7013[30]), .D0(d6[66]), 
          .A1(d_d6[67]), .B1(n7012), .C1(n7013[31]), .D1(d6[67]), .CIN(n11366), 
          .COUT(n11367), .S0(d7_71__N_1531[66]), .S1(d7_71__N_1531[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1135_33.INIT0 = 16'hb874;
    defparam add_1135_33.INIT1 = 16'hb874;
    defparam add_1135_33.INJECT1_0 = "NO";
    defparam add_1135_33.INJECT1_1 = "NO";
    CCU2D add_1135_31 (.A0(d_d6[64]), .B0(n7012), .C0(n7013[28]), .D0(d6[64]), 
          .A1(d_d6[65]), .B1(n7012), .C1(n7013[29]), .D1(d6[65]), .CIN(n11365), 
          .COUT(n11366), .S0(d7_71__N_1531[64]), .S1(d7_71__N_1531[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1135_31.INIT0 = 16'hb874;
    defparam add_1135_31.INIT1 = 16'hb874;
    defparam add_1135_31.INJECT1_0 = "NO";
    defparam add_1135_31.INJECT1_1 = "NO";
    CCU2D add_1135_29 (.A0(d_d6[62]), .B0(n7012), .C0(n7013[26]), .D0(d6[62]), 
          .A1(d_d6[63]), .B1(n7012), .C1(n7013[27]), .D1(d6[63]), .CIN(n11364), 
          .COUT(n11365), .S0(d7_71__N_1531[62]), .S1(d7_71__N_1531[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1135_29.INIT0 = 16'hb874;
    defparam add_1135_29.INIT1 = 16'hb874;
    defparam add_1135_29.INJECT1_0 = "NO";
    defparam add_1135_29.INJECT1_1 = "NO";
    CCU2D add_1135_27 (.A0(d_d6[60]), .B0(n7012), .C0(n7013[24]), .D0(d6[60]), 
          .A1(d_d6[61]), .B1(n7012), .C1(n7013[25]), .D1(d6[61]), .CIN(n11363), 
          .COUT(n11364), .S0(d7_71__N_1531[60]), .S1(d7_71__N_1531[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1135_27.INIT0 = 16'hb874;
    defparam add_1135_27.INIT1 = 16'hb874;
    defparam add_1135_27.INJECT1_0 = "NO";
    defparam add_1135_27.INJECT1_1 = "NO";
    CCU2D add_1135_25 (.A0(d_d6[58]), .B0(n7012), .C0(n7013[22]), .D0(d6[58]), 
          .A1(d_d6[59]), .B1(n7012), .C1(n7013[23]), .D1(d6[59]), .CIN(n11362), 
          .COUT(n11363), .S0(d7_71__N_1531[58]), .S1(d7_71__N_1531[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1135_25.INIT0 = 16'hb874;
    defparam add_1135_25.INIT1 = 16'hb874;
    defparam add_1135_25.INJECT1_0 = "NO";
    defparam add_1135_25.INJECT1_1 = "NO";
    CCU2D add_1135_23 (.A0(d_d6[56]), .B0(n7012), .C0(n7013[20]), .D0(d6[56]), 
          .A1(d_d6[57]), .B1(n7012), .C1(n7013[21]), .D1(d6[57]), .CIN(n11361), 
          .COUT(n11362), .S0(d7_71__N_1531[56]), .S1(d7_71__N_1531[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1135_23.INIT0 = 16'hb874;
    defparam add_1135_23.INIT1 = 16'hb874;
    defparam add_1135_23.INJECT1_0 = "NO";
    defparam add_1135_23.INJECT1_1 = "NO";
    CCU2D add_1135_21 (.A0(d_d6[54]), .B0(n7012), .C0(n7013[18]), .D0(d6[54]), 
          .A1(d_d6[55]), .B1(n7012), .C1(n7013[19]), .D1(d6[55]), .CIN(n11360), 
          .COUT(n11361), .S0(d7_71__N_1531[54]), .S1(d7_71__N_1531[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1135_21.INIT0 = 16'hb874;
    defparam add_1135_21.INIT1 = 16'hb874;
    defparam add_1135_21.INJECT1_0 = "NO";
    defparam add_1135_21.INJECT1_1 = "NO";
    CCU2D add_1135_19 (.A0(d_d6[52]), .B0(n7012), .C0(n7013[16]), .D0(d6[52]), 
          .A1(d_d6[53]), .B1(n7012), .C1(n7013[17]), .D1(d6[53]), .CIN(n11359), 
          .COUT(n11360), .S0(d7_71__N_1531[52]), .S1(d7_71__N_1531[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1135_19.INIT0 = 16'hb874;
    defparam add_1135_19.INIT1 = 16'hb874;
    defparam add_1135_19.INJECT1_0 = "NO";
    defparam add_1135_19.INJECT1_1 = "NO";
    CCU2D add_1135_17 (.A0(d_d6[50]), .B0(n7012), .C0(n7013[14]), .D0(d6[50]), 
          .A1(d_d6[51]), .B1(n7012), .C1(n7013[15]), .D1(d6[51]), .CIN(n11358), 
          .COUT(n11359), .S0(d7_71__N_1531[50]), .S1(d7_71__N_1531[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1135_17.INIT0 = 16'hb874;
    defparam add_1135_17.INIT1 = 16'hb874;
    defparam add_1135_17.INJECT1_0 = "NO";
    defparam add_1135_17.INJECT1_1 = "NO";
    CCU2D add_1135_15 (.A0(d_d6[48]), .B0(n7012), .C0(n7013[12]), .D0(d6[48]), 
          .A1(d_d6[49]), .B1(n7012), .C1(n7013[13]), .D1(d6[49]), .CIN(n11357), 
          .COUT(n11358), .S0(d7_71__N_1531[48]), .S1(d7_71__N_1531[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1135_15.INIT0 = 16'hb874;
    defparam add_1135_15.INIT1 = 16'hb874;
    defparam add_1135_15.INJECT1_0 = "NO";
    defparam add_1135_15.INJECT1_1 = "NO";
    CCU2D add_1135_13 (.A0(d_d6[46]), .B0(n7012), .C0(n7013[10]), .D0(d6[46]), 
          .A1(d_d6[47]), .B1(n7012), .C1(n7013[11]), .D1(d6[47]), .CIN(n11356), 
          .COUT(n11357), .S0(d7_71__N_1531[46]), .S1(d7_71__N_1531[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1135_13.INIT0 = 16'hb874;
    defparam add_1135_13.INIT1 = 16'hb874;
    defparam add_1135_13.INJECT1_0 = "NO";
    defparam add_1135_13.INJECT1_1 = "NO";
    CCU2D add_1135_11 (.A0(d_d6[44]), .B0(n7012), .C0(n7013[8]), .D0(d6[44]), 
          .A1(d_d6[45]), .B1(n7012), .C1(n7013[9]), .D1(d6[45]), .CIN(n11355), 
          .COUT(n11356), .S0(d7_71__N_1531[44]), .S1(d7_71__N_1531[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1135_11.INIT0 = 16'hb874;
    defparam add_1135_11.INIT1 = 16'hb874;
    defparam add_1135_11.INJECT1_0 = "NO";
    defparam add_1135_11.INJECT1_1 = "NO";
    CCU2D add_1135_9 (.A0(d_d6[42]), .B0(n7012), .C0(n7013[6]), .D0(d6[42]), 
          .A1(d_d6[43]), .B1(n7012), .C1(n7013[7]), .D1(d6[43]), .CIN(n11354), 
          .COUT(n11355), .S0(d7_71__N_1531[42]), .S1(d7_71__N_1531[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1135_9.INIT0 = 16'hb874;
    defparam add_1135_9.INIT1 = 16'hb874;
    defparam add_1135_9.INJECT1_0 = "NO";
    defparam add_1135_9.INJECT1_1 = "NO";
    CCU2D add_1135_7 (.A0(d_d6[40]), .B0(n7012), .C0(n7013[4]), .D0(d6[40]), 
          .A1(d_d6[41]), .B1(n7012), .C1(n7013[5]), .D1(d6[41]), .CIN(n11353), 
          .COUT(n11354), .S0(d7_71__N_1531[40]), .S1(d7_71__N_1531[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1135_7.INIT0 = 16'hb874;
    defparam add_1135_7.INIT1 = 16'hb874;
    defparam add_1135_7.INJECT1_0 = "NO";
    defparam add_1135_7.INJECT1_1 = "NO";
    CCU2D add_1135_5 (.A0(d_d6[38]), .B0(n7012), .C0(n7013[2]), .D0(d6[38]), 
          .A1(d_d6[39]), .B1(n7012), .C1(n7013[3]), .D1(d6[39]), .CIN(n11352), 
          .COUT(n11353), .S0(d7_71__N_1531[38]), .S1(d7_71__N_1531[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1135_5.INIT0 = 16'hb874;
    defparam add_1135_5.INIT1 = 16'hb874;
    defparam add_1135_5.INJECT1_0 = "NO";
    defparam add_1135_5.INJECT1_1 = "NO";
    CCU2D add_1135_3 (.A0(d_d6[36]), .B0(n7012), .C0(n7013[0]), .D0(d6[36]), 
          .A1(d_d6[37]), .B1(n7012), .C1(n7013[1]), .D1(d6[37]), .CIN(n11351), 
          .COUT(n11352), .S0(d7_71__N_1531[36]), .S1(d7_71__N_1531[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1135_3.INIT0 = 16'hb874;
    defparam add_1135_3.INIT1 = 16'hb874;
    defparam add_1135_3.INJECT1_0 = "NO";
    defparam add_1135_3.INJECT1_1 = "NO";
    CCU2D add_1135_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n7012), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11351));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1135_1.INIT0 = 16'hF000;
    defparam add_1135_1.INIT1 = 16'h0555;
    defparam add_1135_1.INJECT1_0 = "NO";
    defparam add_1135_1.INJECT1_1 = "NO";
    CCU2D add_1038_37 (.A0(d_tmp[35]), .B0(d_d_tmp[35]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11262), .S0(d6_71__N_1459[35]), .S1(n4124));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1038_37.INIT0 = 16'h5999;
    defparam add_1038_37.INIT1 = 16'h0000;
    defparam add_1038_37.INJECT1_0 = "NO";
    defparam add_1038_37.INJECT1_1 = "NO";
    CCU2D add_1038_35 (.A0(d_tmp[33]), .B0(d_d_tmp[33]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[34]), .B1(d_d_tmp[34]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11261), .COUT(n11262), .S0(d6_71__N_1459[33]), 
          .S1(d6_71__N_1459[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1038_35.INIT0 = 16'h5999;
    defparam add_1038_35.INIT1 = 16'h5999;
    defparam add_1038_35.INJECT1_0 = "NO";
    defparam add_1038_35.INJECT1_1 = "NO";
    CCU2D add_1038_33 (.A0(d_tmp[31]), .B0(d_d_tmp[31]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[32]), .B1(d_d_tmp[32]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11260), .COUT(n11261), .S0(d6_71__N_1459[31]), 
          .S1(d6_71__N_1459[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1038_33.INIT0 = 16'h5999;
    defparam add_1038_33.INIT1 = 16'h5999;
    defparam add_1038_33.INJECT1_0 = "NO";
    defparam add_1038_33.INJECT1_1 = "NO";
    CCU2D add_1038_31 (.A0(d_tmp[29]), .B0(d_d_tmp[29]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[30]), .B1(d_d_tmp[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11259), .COUT(n11260), .S0(d6_71__N_1459[29]), 
          .S1(d6_71__N_1459[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1038_31.INIT0 = 16'h5999;
    defparam add_1038_31.INIT1 = 16'h5999;
    defparam add_1038_31.INJECT1_0 = "NO";
    defparam add_1038_31.INJECT1_1 = "NO";
    CCU2D add_1038_29 (.A0(d_tmp[27]), .B0(d_d_tmp[27]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[28]), .B1(d_d_tmp[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11258), .COUT(n11259), .S0(d6_71__N_1459[27]), 
          .S1(d6_71__N_1459[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1038_29.INIT0 = 16'h5999;
    defparam add_1038_29.INIT1 = 16'h5999;
    defparam add_1038_29.INJECT1_0 = "NO";
    defparam add_1038_29.INJECT1_1 = "NO";
    CCU2D add_1038_27 (.A0(d_tmp[25]), .B0(d_d_tmp[25]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[26]), .B1(d_d_tmp[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11257), .COUT(n11258), .S0(d6_71__N_1459[25]), 
          .S1(d6_71__N_1459[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1038_27.INIT0 = 16'h5999;
    defparam add_1038_27.INIT1 = 16'h5999;
    defparam add_1038_27.INJECT1_0 = "NO";
    defparam add_1038_27.INJECT1_1 = "NO";
    CCU2D add_1038_25 (.A0(d_tmp[23]), .B0(d_d_tmp[23]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[24]), .B1(d_d_tmp[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11256), .COUT(n11257), .S0(d6_71__N_1459[23]), 
          .S1(d6_71__N_1459[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1038_25.INIT0 = 16'h5999;
    defparam add_1038_25.INIT1 = 16'h5999;
    defparam add_1038_25.INJECT1_0 = "NO";
    defparam add_1038_25.INJECT1_1 = "NO";
    CCU2D add_1038_23 (.A0(d_tmp[21]), .B0(d_d_tmp[21]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[22]), .B1(d_d_tmp[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11255), .COUT(n11256), .S0(d6_71__N_1459[21]), 
          .S1(d6_71__N_1459[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1038_23.INIT0 = 16'h5999;
    defparam add_1038_23.INIT1 = 16'h5999;
    defparam add_1038_23.INJECT1_0 = "NO";
    defparam add_1038_23.INJECT1_1 = "NO";
    CCU2D add_1038_21 (.A0(d_tmp[19]), .B0(d_d_tmp[19]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[20]), .B1(d_d_tmp[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11254), .COUT(n11255), .S0(d6_71__N_1459[19]), 
          .S1(d6_71__N_1459[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1038_21.INIT0 = 16'h5999;
    defparam add_1038_21.INIT1 = 16'h5999;
    defparam add_1038_21.INJECT1_0 = "NO";
    defparam add_1038_21.INJECT1_1 = "NO";
    CCU2D add_1038_19 (.A0(d_tmp[17]), .B0(d_d_tmp[17]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[18]), .B1(d_d_tmp[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11253), .COUT(n11254), .S0(d6_71__N_1459[17]), 
          .S1(d6_71__N_1459[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1038_19.INIT0 = 16'h5999;
    defparam add_1038_19.INIT1 = 16'h5999;
    defparam add_1038_19.INJECT1_0 = "NO";
    defparam add_1038_19.INJECT1_1 = "NO";
    CCU2D add_1038_17 (.A0(d_tmp[15]), .B0(d_d_tmp[15]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[16]), .B1(d_d_tmp[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11252), .COUT(n11253), .S0(d6_71__N_1459[15]), 
          .S1(d6_71__N_1459[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1038_17.INIT0 = 16'h5999;
    defparam add_1038_17.INIT1 = 16'h5999;
    defparam add_1038_17.INJECT1_0 = "NO";
    defparam add_1038_17.INJECT1_1 = "NO";
    CCU2D add_1038_15 (.A0(d_tmp[13]), .B0(d_d_tmp[13]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[14]), .B1(d_d_tmp[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11251), .COUT(n11252), .S0(d6_71__N_1459[13]), 
          .S1(d6_71__N_1459[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1038_15.INIT0 = 16'h5999;
    defparam add_1038_15.INIT1 = 16'h5999;
    defparam add_1038_15.INJECT1_0 = "NO";
    defparam add_1038_15.INJECT1_1 = "NO";
    CCU2D add_1038_13 (.A0(d_tmp[11]), .B0(d_d_tmp[11]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[12]), .B1(d_d_tmp[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11250), .COUT(n11251), .S0(d6_71__N_1459[11]), 
          .S1(d6_71__N_1459[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1038_13.INIT0 = 16'h5999;
    defparam add_1038_13.INIT1 = 16'h5999;
    defparam add_1038_13.INJECT1_0 = "NO";
    defparam add_1038_13.INJECT1_1 = "NO";
    CCU2D add_1038_11 (.A0(d_tmp[9]), .B0(d_d_tmp[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[10]), .B1(d_d_tmp[10]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11249), .COUT(n11250), .S0(d6_71__N_1459[9]), .S1(d6_71__N_1459[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1038_11.INIT0 = 16'h5999;
    defparam add_1038_11.INIT1 = 16'h5999;
    defparam add_1038_11.INJECT1_0 = "NO";
    defparam add_1038_11.INJECT1_1 = "NO";
    CCU2D add_1038_9 (.A0(d_tmp[7]), .B0(d_d_tmp[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[8]), .B1(d_d_tmp[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11248), .COUT(n11249), .S0(d6_71__N_1459[7]), .S1(d6_71__N_1459[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1038_9.INIT0 = 16'h5999;
    defparam add_1038_9.INIT1 = 16'h5999;
    defparam add_1038_9.INJECT1_0 = "NO";
    defparam add_1038_9.INJECT1_1 = "NO";
    CCU2D add_1038_7 (.A0(d_tmp[5]), .B0(d_d_tmp[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[6]), .B1(d_d_tmp[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11247), .COUT(n11248), .S0(d6_71__N_1459[5]), .S1(d6_71__N_1459[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1038_7.INIT0 = 16'h5999;
    defparam add_1038_7.INIT1 = 16'h5999;
    defparam add_1038_7.INJECT1_0 = "NO";
    defparam add_1038_7.INJECT1_1 = "NO";
    CCU2D add_1038_5 (.A0(d_tmp[3]), .B0(d_d_tmp[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[4]), .B1(d_d_tmp[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11246), .COUT(n11247), .S0(d6_71__N_1459[3]), .S1(d6_71__N_1459[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1038_5.INIT0 = 16'h5999;
    defparam add_1038_5.INIT1 = 16'h5999;
    defparam add_1038_5.INJECT1_0 = "NO";
    defparam add_1038_5.INJECT1_1 = "NO";
    CCU2D add_1038_3 (.A0(d_tmp[1]), .B0(d_d_tmp[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[2]), .B1(d_d_tmp[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11245), .COUT(n11246), .S0(d6_71__N_1459[1]), .S1(d6_71__N_1459[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1038_3.INIT0 = 16'h5999;
    defparam add_1038_3.INIT1 = 16'h5999;
    defparam add_1038_3.INJECT1_0 = "NO";
    defparam add_1038_3.INJECT1_1 = "NO";
    CCU2D add_1038_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[0]), .B1(d_d_tmp[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n11245), .S1(d6_71__N_1459[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1038_1.INIT0 = 16'h0000;
    defparam add_1038_1.INIT1 = 16'h5999;
    defparam add_1038_1.INJECT1_0 = "NO";
    defparam add_1038_1.INJECT1_1 = "NO";
    CCU2D add_1093_37 (.A0(d8[35]), .B0(d_d8[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11223), 
          .S0(d9_71__N_1675[35]), .S1(n5796));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1093_37.INIT0 = 16'h5999;
    defparam add_1093_37.INIT1 = 16'h0000;
    defparam add_1093_37.INJECT1_0 = "NO";
    defparam add_1093_37.INJECT1_1 = "NO";
    CCU2D add_1093_35 (.A0(d8[33]), .B0(d_d8[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[34]), .B1(d_d8[34]), .C1(GND_net), .D1(GND_net), .CIN(n11222), 
          .COUT(n11223), .S0(d9_71__N_1675[33]), .S1(d9_71__N_1675[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1093_35.INIT0 = 16'h5999;
    defparam add_1093_35.INIT1 = 16'h5999;
    defparam add_1093_35.INJECT1_0 = "NO";
    defparam add_1093_35.INJECT1_1 = "NO";
    CCU2D add_1093_33 (.A0(d8[31]), .B0(d_d8[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[32]), .B1(d_d8[32]), .C1(GND_net), .D1(GND_net), .CIN(n11221), 
          .COUT(n11222), .S0(d9_71__N_1675[31]), .S1(d9_71__N_1675[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1093_33.INIT0 = 16'h5999;
    defparam add_1093_33.INIT1 = 16'h5999;
    defparam add_1093_33.INJECT1_0 = "NO";
    defparam add_1093_33.INJECT1_1 = "NO";
    CCU2D add_1093_31 (.A0(d8[29]), .B0(d_d8[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[30]), .B1(d_d8[30]), .C1(GND_net), .D1(GND_net), .CIN(n11220), 
          .COUT(n11221), .S0(d9_71__N_1675[29]), .S1(d9_71__N_1675[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1093_31.INIT0 = 16'h5999;
    defparam add_1093_31.INIT1 = 16'h5999;
    defparam add_1093_31.INJECT1_0 = "NO";
    defparam add_1093_31.INJECT1_1 = "NO";
    CCU2D add_1093_29 (.A0(d8[27]), .B0(d_d8[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[28]), .B1(d_d8[28]), .C1(GND_net), .D1(GND_net), .CIN(n11219), 
          .COUT(n11220), .S0(d9_71__N_1675[27]), .S1(d9_71__N_1675[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1093_29.INIT0 = 16'h5999;
    defparam add_1093_29.INIT1 = 16'h5999;
    defparam add_1093_29.INJECT1_0 = "NO";
    defparam add_1093_29.INJECT1_1 = "NO";
    CCU2D add_1093_27 (.A0(d8[25]), .B0(d_d8[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[26]), .B1(d_d8[26]), .C1(GND_net), .D1(GND_net), .CIN(n11218), 
          .COUT(n11219), .S0(d9_71__N_1675[25]), .S1(d9_71__N_1675[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1093_27.INIT0 = 16'h5999;
    defparam add_1093_27.INIT1 = 16'h5999;
    defparam add_1093_27.INJECT1_0 = "NO";
    defparam add_1093_27.INJECT1_1 = "NO";
    CCU2D add_1093_25 (.A0(d8[23]), .B0(d_d8[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[24]), .B1(d_d8[24]), .C1(GND_net), .D1(GND_net), .CIN(n11217), 
          .COUT(n11218), .S0(d9_71__N_1675[23]), .S1(d9_71__N_1675[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1093_25.INIT0 = 16'h5999;
    defparam add_1093_25.INIT1 = 16'h5999;
    defparam add_1093_25.INJECT1_0 = "NO";
    defparam add_1093_25.INJECT1_1 = "NO";
    CCU2D add_1093_23 (.A0(d8[21]), .B0(d_d8[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[22]), .B1(d_d8[22]), .C1(GND_net), .D1(GND_net), .CIN(n11216), 
          .COUT(n11217), .S0(d9_71__N_1675[21]), .S1(d9_71__N_1675[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1093_23.INIT0 = 16'h5999;
    defparam add_1093_23.INIT1 = 16'h5999;
    defparam add_1093_23.INJECT1_0 = "NO";
    defparam add_1093_23.INJECT1_1 = "NO";
    CCU2D add_1093_21 (.A0(d8[19]), .B0(d_d8[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[20]), .B1(d_d8[20]), .C1(GND_net), .D1(GND_net), .CIN(n11215), 
          .COUT(n11216), .S0(d9_71__N_1675[19]), .S1(d9_71__N_1675[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1093_21.INIT0 = 16'h5999;
    defparam add_1093_21.INIT1 = 16'h5999;
    defparam add_1093_21.INJECT1_0 = "NO";
    defparam add_1093_21.INJECT1_1 = "NO";
    CCU2D add_1093_19 (.A0(d8[17]), .B0(d_d8[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[18]), .B1(d_d8[18]), .C1(GND_net), .D1(GND_net), .CIN(n11214), 
          .COUT(n11215), .S0(d9_71__N_1675[17]), .S1(d9_71__N_1675[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1093_19.INIT0 = 16'h5999;
    defparam add_1093_19.INIT1 = 16'h5999;
    defparam add_1093_19.INJECT1_0 = "NO";
    defparam add_1093_19.INJECT1_1 = "NO";
    CCU2D add_1093_17 (.A0(d8[15]), .B0(d_d8[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[16]), .B1(d_d8[16]), .C1(GND_net), .D1(GND_net), .CIN(n11213), 
          .COUT(n11214), .S0(d9_71__N_1675[15]), .S1(d9_71__N_1675[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1093_17.INIT0 = 16'h5999;
    defparam add_1093_17.INIT1 = 16'h5999;
    defparam add_1093_17.INJECT1_0 = "NO";
    defparam add_1093_17.INJECT1_1 = "NO";
    CCU2D add_1093_15 (.A0(d8[13]), .B0(d_d8[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[14]), .B1(d_d8[14]), .C1(GND_net), .D1(GND_net), .CIN(n11212), 
          .COUT(n11213), .S0(d9_71__N_1675[13]), .S1(d9_71__N_1675[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1093_15.INIT0 = 16'h5999;
    defparam add_1093_15.INIT1 = 16'h5999;
    defparam add_1093_15.INJECT1_0 = "NO";
    defparam add_1093_15.INJECT1_1 = "NO";
    CCU2D add_1093_13 (.A0(d8[11]), .B0(d_d8[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[12]), .B1(d_d8[12]), .C1(GND_net), .D1(GND_net), .CIN(n11211), 
          .COUT(n11212), .S0(d9_71__N_1675[11]), .S1(d9_71__N_1675[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1093_13.INIT0 = 16'h5999;
    defparam add_1093_13.INIT1 = 16'h5999;
    defparam add_1093_13.INJECT1_0 = "NO";
    defparam add_1093_13.INJECT1_1 = "NO";
    CCU2D add_1093_11 (.A0(d8[9]), .B0(d_d8[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[10]), .B1(d_d8[10]), .C1(GND_net), .D1(GND_net), .CIN(n11210), 
          .COUT(n11211), .S0(d9_71__N_1675[9]), .S1(d9_71__N_1675[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1093_11.INIT0 = 16'h5999;
    defparam add_1093_11.INIT1 = 16'h5999;
    defparam add_1093_11.INJECT1_0 = "NO";
    defparam add_1093_11.INJECT1_1 = "NO";
    CCU2D add_1093_9 (.A0(d8[7]), .B0(d_d8[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[8]), .B1(d_d8[8]), .C1(GND_net), .D1(GND_net), .CIN(n11209), 
          .COUT(n11210), .S0(d9_71__N_1675[7]), .S1(d9_71__N_1675[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1093_9.INIT0 = 16'h5999;
    defparam add_1093_9.INIT1 = 16'h5999;
    defparam add_1093_9.INJECT1_0 = "NO";
    defparam add_1093_9.INJECT1_1 = "NO";
    CCU2D add_1093_7 (.A0(d8[5]), .B0(d_d8[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[6]), .B1(d_d8[6]), .C1(GND_net), .D1(GND_net), .CIN(n11208), 
          .COUT(n11209), .S0(d9_71__N_1675[5]), .S1(d9_71__N_1675[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1093_7.INIT0 = 16'h5999;
    defparam add_1093_7.INIT1 = 16'h5999;
    defparam add_1093_7.INJECT1_0 = "NO";
    defparam add_1093_7.INJECT1_1 = "NO";
    CCU2D add_1093_5 (.A0(d8[3]), .B0(d_d8[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[4]), .B1(d_d8[4]), .C1(GND_net), .D1(GND_net), .CIN(n11207), 
          .COUT(n11208), .S0(d9_71__N_1675[3]), .S1(d9_71__N_1675[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1093_5.INIT0 = 16'h5999;
    defparam add_1093_5.INIT1 = 16'h5999;
    defparam add_1093_5.INJECT1_0 = "NO";
    defparam add_1093_5.INJECT1_1 = "NO";
    CCU2D add_1093_3 (.A0(d8[1]), .B0(d_d8[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[2]), .B1(d_d8[2]), .C1(GND_net), .D1(GND_net), .CIN(n11206), 
          .COUT(n11207), .S0(d9_71__N_1675[1]), .S1(d9_71__N_1675[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1093_3.INIT0 = 16'h5999;
    defparam add_1093_3.INIT1 = 16'h5999;
    defparam add_1093_3.INJECT1_0 = "NO";
    defparam add_1093_3.INJECT1_1 = "NO";
    CCU2D add_1093_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d8[0]), .B1(d_d8[0]), .C1(GND_net), .D1(GND_net), .COUT(n11206), 
          .S1(d9_71__N_1675[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1093_1.INIT0 = 16'h0000;
    defparam add_1093_1.INIT1 = 16'h5999;
    defparam add_1093_1.INJECT1_0 = "NO";
    defparam add_1093_1.INJECT1_1 = "NO";
    CCU2D add_10_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11099), 
          .S0(n375[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_17.INIT0 = 16'h5aaa;
    defparam add_10_17.INIT1 = 16'h0000;
    defparam add_10_17.INJECT1_0 = "NO";
    defparam add_10_17.INJECT1_1 = "NO";
    CCU2D add_10_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11098), .COUT(n11099), .S0(n375[13]), .S1(n375[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_15.INIT0 = 16'h5aaa;
    defparam add_10_15.INIT1 = 16'h5aaa;
    defparam add_10_15.INJECT1_0 = "NO";
    defparam add_10_15.INJECT1_1 = "NO";
    CCU2D add_10_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11097), .COUT(n11098), .S0(n375[11]), .S1(n375[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_13.INIT0 = 16'h5aaa;
    defparam add_10_13.INIT1 = 16'h5aaa;
    defparam add_10_13.INJECT1_0 = "NO";
    defparam add_10_13.INJECT1_1 = "NO";
    CCU2D add_10_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11096), .COUT(n11097), .S0(n375[9]), .S1(n375[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_11.INIT0 = 16'h5aaa;
    defparam add_10_11.INIT1 = 16'h5aaa;
    defparam add_10_11.INJECT1_0 = "NO";
    defparam add_10_11.INJECT1_1 = "NO";
    CCU2D add_10_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11095), 
          .COUT(n11096), .S0(n375[7]), .S1(n375[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_9.INIT0 = 16'h5aaa;
    defparam add_10_9.INIT1 = 16'h5aaa;
    defparam add_10_9.INJECT1_0 = "NO";
    defparam add_10_9.INJECT1_1 = "NO";
    CCU2D add_10_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11094), 
          .COUT(n11095), .S0(n375[5]), .S1(n375[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_7.INIT0 = 16'h5aaa;
    defparam add_10_7.INIT1 = 16'h5aaa;
    defparam add_10_7.INJECT1_0 = "NO";
    defparam add_10_7.INJECT1_1 = "NO";
    CCU2D add_10_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11093), 
          .COUT(n11094), .S0(n375[3]), .S1(n375[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_5.INIT0 = 16'h5aaa;
    defparam add_10_5.INIT1 = 16'h5aaa;
    defparam add_10_5.INJECT1_0 = "NO";
    defparam add_10_5.INJECT1_1 = "NO";
    CCU2D add_10_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11092), 
          .COUT(n11093), .S0(n375[1]), .S1(n375[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_3.INIT0 = 16'h5aaa;
    defparam add_10_3.INIT1 = 16'h5aaa;
    defparam add_10_3.INJECT1_0 = "NO";
    defparam add_10_3.INJECT1_1 = "NO";
    CCU2D add_10_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11092), 
          .S1(n375[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_1.INIT0 = 16'hF000;
    defparam add_10_1.INIT1 = 16'h5555;
    defparam add_10_1.INJECT1_0 = "NO";
    defparam add_10_1.INJECT1_1 = "NO";
    CCU2D add_1063_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11072), 
          .S0(n4884));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1063_cout.INIT0 = 16'h0000;
    defparam add_1063_cout.INIT1 = 16'h0000;
    defparam add_1063_cout.INJECT1_0 = "NO";
    defparam add_1063_cout.INJECT1_1 = "NO";
    CCU2D add_1063_36 (.A0(d4[34]), .B0(d5[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[35]), .B1(d5[35]), .C1(GND_net), .D1(GND_net), .CIN(n11071), 
          .COUT(n11072), .S0(d5_71__N_706[34]), .S1(d5_71__N_706[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1063_36.INIT0 = 16'h5666;
    defparam add_1063_36.INIT1 = 16'h5666;
    defparam add_1063_36.INJECT1_0 = "NO";
    defparam add_1063_36.INJECT1_1 = "NO";
    CCU2D add_1063_34 (.A0(d4[32]), .B0(d5[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[33]), .B1(d5[33]), .C1(GND_net), .D1(GND_net), .CIN(n11070), 
          .COUT(n11071), .S0(d5_71__N_706[32]), .S1(d5_71__N_706[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1063_34.INIT0 = 16'h5666;
    defparam add_1063_34.INIT1 = 16'h5666;
    defparam add_1063_34.INJECT1_0 = "NO";
    defparam add_1063_34.INJECT1_1 = "NO";
    CCU2D add_1063_32 (.A0(d4[30]), .B0(d5[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[31]), .B1(d5[31]), .C1(GND_net), .D1(GND_net), .CIN(n11069), 
          .COUT(n11070), .S0(d5_71__N_706[30]), .S1(d5_71__N_706[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1063_32.INIT0 = 16'h5666;
    defparam add_1063_32.INIT1 = 16'h5666;
    defparam add_1063_32.INJECT1_0 = "NO";
    defparam add_1063_32.INJECT1_1 = "NO";
    CCU2D add_1063_30 (.A0(d4[28]), .B0(d5[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[29]), .B1(d5[29]), .C1(GND_net), .D1(GND_net), .CIN(n11068), 
          .COUT(n11069), .S0(d5_71__N_706[28]), .S1(d5_71__N_706[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1063_30.INIT0 = 16'h5666;
    defparam add_1063_30.INIT1 = 16'h5666;
    defparam add_1063_30.INJECT1_0 = "NO";
    defparam add_1063_30.INJECT1_1 = "NO";
    CCU2D add_1063_28 (.A0(d4[26]), .B0(d5[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[27]), .B1(d5[27]), .C1(GND_net), .D1(GND_net), .CIN(n11067), 
          .COUT(n11068), .S0(d5_71__N_706[26]), .S1(d5_71__N_706[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1063_28.INIT0 = 16'h5666;
    defparam add_1063_28.INIT1 = 16'h5666;
    defparam add_1063_28.INJECT1_0 = "NO";
    defparam add_1063_28.INJECT1_1 = "NO";
    CCU2D add_1063_26 (.A0(d4[24]), .B0(d5[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[25]), .B1(d5[25]), .C1(GND_net), .D1(GND_net), .CIN(n11066), 
          .COUT(n11067), .S0(d5_71__N_706[24]), .S1(d5_71__N_706[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1063_26.INIT0 = 16'h5666;
    defparam add_1063_26.INIT1 = 16'h5666;
    defparam add_1063_26.INJECT1_0 = "NO";
    defparam add_1063_26.INJECT1_1 = "NO";
    CCU2D add_1063_24 (.A0(d4[22]), .B0(d5[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[23]), .B1(d5[23]), .C1(GND_net), .D1(GND_net), .CIN(n11065), 
          .COUT(n11066), .S0(d5_71__N_706[22]), .S1(d5_71__N_706[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1063_24.INIT0 = 16'h5666;
    defparam add_1063_24.INIT1 = 16'h5666;
    defparam add_1063_24.INJECT1_0 = "NO";
    defparam add_1063_24.INJECT1_1 = "NO";
    CCU2D add_1063_22 (.A0(d4[20]), .B0(d5[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[21]), .B1(d5[21]), .C1(GND_net), .D1(GND_net), .CIN(n11064), 
          .COUT(n11065), .S0(d5_71__N_706[20]), .S1(d5_71__N_706[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1063_22.INIT0 = 16'h5666;
    defparam add_1063_22.INIT1 = 16'h5666;
    defparam add_1063_22.INJECT1_0 = "NO";
    defparam add_1063_22.INJECT1_1 = "NO";
    CCU2D add_1063_20 (.A0(d4[18]), .B0(d5[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[19]), .B1(d5[19]), .C1(GND_net), .D1(GND_net), .CIN(n11063), 
          .COUT(n11064), .S0(d5_71__N_706[18]), .S1(d5_71__N_706[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1063_20.INIT0 = 16'h5666;
    defparam add_1063_20.INIT1 = 16'h5666;
    defparam add_1063_20.INJECT1_0 = "NO";
    defparam add_1063_20.INJECT1_1 = "NO";
    CCU2D add_1063_18 (.A0(d4[16]), .B0(d5[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[17]), .B1(d5[17]), .C1(GND_net), .D1(GND_net), .CIN(n11062), 
          .COUT(n11063), .S0(d5_71__N_706[16]), .S1(d5_71__N_706[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1063_18.INIT0 = 16'h5666;
    defparam add_1063_18.INIT1 = 16'h5666;
    defparam add_1063_18.INJECT1_0 = "NO";
    defparam add_1063_18.INJECT1_1 = "NO";
    CCU2D add_1063_16 (.A0(d4[14]), .B0(d5[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[15]), .B1(d5[15]), .C1(GND_net), .D1(GND_net), .CIN(n11061), 
          .COUT(n11062), .S0(d5_71__N_706[14]), .S1(d5_71__N_706[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1063_16.INIT0 = 16'h5666;
    defparam add_1063_16.INIT1 = 16'h5666;
    defparam add_1063_16.INJECT1_0 = "NO";
    defparam add_1063_16.INJECT1_1 = "NO";
    CCU2D add_1063_14 (.A0(d4[12]), .B0(d5[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[13]), .B1(d5[13]), .C1(GND_net), .D1(GND_net), .CIN(n11060), 
          .COUT(n11061), .S0(d5_71__N_706[12]), .S1(d5_71__N_706[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1063_14.INIT0 = 16'h5666;
    defparam add_1063_14.INIT1 = 16'h5666;
    defparam add_1063_14.INJECT1_0 = "NO";
    defparam add_1063_14.INJECT1_1 = "NO";
    CCU2D add_1063_12 (.A0(d4[10]), .B0(d5[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[11]), .B1(d5[11]), .C1(GND_net), .D1(GND_net), .CIN(n11059), 
          .COUT(n11060), .S0(d5_71__N_706[10]), .S1(d5_71__N_706[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1063_12.INIT0 = 16'h5666;
    defparam add_1063_12.INIT1 = 16'h5666;
    defparam add_1063_12.INJECT1_0 = "NO";
    defparam add_1063_12.INJECT1_1 = "NO";
    CCU2D add_1063_10 (.A0(d4[8]), .B0(d5[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[9]), .B1(d5[9]), .C1(GND_net), .D1(GND_net), .CIN(n11058), 
          .COUT(n11059), .S0(d5_71__N_706[8]), .S1(d5_71__N_706[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1063_10.INIT0 = 16'h5666;
    defparam add_1063_10.INIT1 = 16'h5666;
    defparam add_1063_10.INJECT1_0 = "NO";
    defparam add_1063_10.INJECT1_1 = "NO";
    CCU2D add_1063_8 (.A0(d4[6]), .B0(d5[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[7]), .B1(d5[7]), .C1(GND_net), .D1(GND_net), .CIN(n11057), 
          .COUT(n11058), .S0(d5_71__N_706[6]), .S1(d5_71__N_706[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1063_8.INIT0 = 16'h5666;
    defparam add_1063_8.INIT1 = 16'h5666;
    defparam add_1063_8.INJECT1_0 = "NO";
    defparam add_1063_8.INJECT1_1 = "NO";
    CCU2D add_1063_6 (.A0(d4[4]), .B0(d5[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[5]), .B1(d5[5]), .C1(GND_net), .D1(GND_net), .CIN(n11056), 
          .COUT(n11057), .S0(d5_71__N_706[4]), .S1(d5_71__N_706[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1063_6.INIT0 = 16'h5666;
    defparam add_1063_6.INIT1 = 16'h5666;
    defparam add_1063_6.INJECT1_0 = "NO";
    defparam add_1063_6.INJECT1_1 = "NO";
    CCU2D add_1063_4 (.A0(d4[2]), .B0(d5[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[3]), .B1(d5[3]), .C1(GND_net), .D1(GND_net), .CIN(n11055), 
          .COUT(n11056), .S0(d5_71__N_706[2]), .S1(d5_71__N_706[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1063_4.INIT0 = 16'h5666;
    defparam add_1063_4.INIT1 = 16'h5666;
    defparam add_1063_4.INJECT1_0 = "NO";
    defparam add_1063_4.INJECT1_1 = "NO";
    CCU2D add_1063_2 (.A0(d4[0]), .B0(d5[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[1]), .B1(d5[1]), .C1(GND_net), .D1(GND_net), .COUT(n11055), 
          .S1(d5_71__N_706[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1063_2.INIT0 = 16'h7000;
    defparam add_1063_2.INIT1 = 16'h5666;
    defparam add_1063_2.INJECT1_0 = "NO";
    defparam add_1063_2.INJECT1_1 = "NO";
    CCU2D add_1058_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11053), 
          .S0(n4732));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1058_cout.INIT0 = 16'h0000;
    defparam add_1058_cout.INIT1 = 16'h0000;
    defparam add_1058_cout.INJECT1_0 = "NO";
    defparam add_1058_cout.INJECT1_1 = "NO";
    CCU2D add_1058_36 (.A0(d3[34]), .B0(d4[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[35]), .B1(d4[35]), .C1(GND_net), .D1(GND_net), .CIN(n11052), 
          .COUT(n11053), .S0(d4_71__N_634[34]), .S1(d4_71__N_634[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1058_36.INIT0 = 16'h5666;
    defparam add_1058_36.INIT1 = 16'h5666;
    defparam add_1058_36.INJECT1_0 = "NO";
    defparam add_1058_36.INJECT1_1 = "NO";
    CCU2D add_1058_34 (.A0(d3[32]), .B0(d4[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[33]), .B1(d4[33]), .C1(GND_net), .D1(GND_net), .CIN(n11051), 
          .COUT(n11052), .S0(d4_71__N_634[32]), .S1(d4_71__N_634[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1058_34.INIT0 = 16'h5666;
    defparam add_1058_34.INIT1 = 16'h5666;
    defparam add_1058_34.INJECT1_0 = "NO";
    defparam add_1058_34.INJECT1_1 = "NO";
    CCU2D add_1058_32 (.A0(d3[30]), .B0(d4[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[31]), .B1(d4[31]), .C1(GND_net), .D1(GND_net), .CIN(n11050), 
          .COUT(n11051), .S0(d4_71__N_634[30]), .S1(d4_71__N_634[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1058_32.INIT0 = 16'h5666;
    defparam add_1058_32.INIT1 = 16'h5666;
    defparam add_1058_32.INJECT1_0 = "NO";
    defparam add_1058_32.INJECT1_1 = "NO";
    CCU2D add_1058_30 (.A0(d3[28]), .B0(d4[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[29]), .B1(d4[29]), .C1(GND_net), .D1(GND_net), .CIN(n11049), 
          .COUT(n11050), .S0(d4_71__N_634[28]), .S1(d4_71__N_634[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1058_30.INIT0 = 16'h5666;
    defparam add_1058_30.INIT1 = 16'h5666;
    defparam add_1058_30.INJECT1_0 = "NO";
    defparam add_1058_30.INJECT1_1 = "NO";
    CCU2D add_1058_28 (.A0(d3[26]), .B0(d4[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[27]), .B1(d4[27]), .C1(GND_net), .D1(GND_net), .CIN(n11048), 
          .COUT(n11049), .S0(d4_71__N_634[26]), .S1(d4_71__N_634[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1058_28.INIT0 = 16'h5666;
    defparam add_1058_28.INIT1 = 16'h5666;
    defparam add_1058_28.INJECT1_0 = "NO";
    defparam add_1058_28.INJECT1_1 = "NO";
    CCU2D add_1058_26 (.A0(d3[24]), .B0(d4[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[25]), .B1(d4[25]), .C1(GND_net), .D1(GND_net), .CIN(n11047), 
          .COUT(n11048), .S0(d4_71__N_634[24]), .S1(d4_71__N_634[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1058_26.INIT0 = 16'h5666;
    defparam add_1058_26.INIT1 = 16'h5666;
    defparam add_1058_26.INJECT1_0 = "NO";
    defparam add_1058_26.INJECT1_1 = "NO";
    CCU2D add_1058_24 (.A0(d3[22]), .B0(d4[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[23]), .B1(d4[23]), .C1(GND_net), .D1(GND_net), .CIN(n11046), 
          .COUT(n11047), .S0(d4_71__N_634[22]), .S1(d4_71__N_634[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1058_24.INIT0 = 16'h5666;
    defparam add_1058_24.INIT1 = 16'h5666;
    defparam add_1058_24.INJECT1_0 = "NO";
    defparam add_1058_24.INJECT1_1 = "NO";
    CCU2D add_1058_22 (.A0(d3[20]), .B0(d4[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[21]), .B1(d4[21]), .C1(GND_net), .D1(GND_net), .CIN(n11045), 
          .COUT(n11046), .S0(d4_71__N_634[20]), .S1(d4_71__N_634[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1058_22.INIT0 = 16'h5666;
    defparam add_1058_22.INIT1 = 16'h5666;
    defparam add_1058_22.INJECT1_0 = "NO";
    defparam add_1058_22.INJECT1_1 = "NO";
    CCU2D add_1058_20 (.A0(d3[18]), .B0(d4[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[19]), .B1(d4[19]), .C1(GND_net), .D1(GND_net), .CIN(n11044), 
          .COUT(n11045), .S0(d4_71__N_634[18]), .S1(d4_71__N_634[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1058_20.INIT0 = 16'h5666;
    defparam add_1058_20.INIT1 = 16'h5666;
    defparam add_1058_20.INJECT1_0 = "NO";
    defparam add_1058_20.INJECT1_1 = "NO";
    CCU2D add_1058_18 (.A0(d3[16]), .B0(d4[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[17]), .B1(d4[17]), .C1(GND_net), .D1(GND_net), .CIN(n11043), 
          .COUT(n11044), .S0(d4_71__N_634[16]), .S1(d4_71__N_634[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1058_18.INIT0 = 16'h5666;
    defparam add_1058_18.INIT1 = 16'h5666;
    defparam add_1058_18.INJECT1_0 = "NO";
    defparam add_1058_18.INJECT1_1 = "NO";
    CCU2D add_1058_16 (.A0(d3[14]), .B0(d4[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[15]), .B1(d4[15]), .C1(GND_net), .D1(GND_net), .CIN(n11042), 
          .COUT(n11043), .S0(d4_71__N_634[14]), .S1(d4_71__N_634[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1058_16.INIT0 = 16'h5666;
    defparam add_1058_16.INIT1 = 16'h5666;
    defparam add_1058_16.INJECT1_0 = "NO";
    defparam add_1058_16.INJECT1_1 = "NO";
    CCU2D add_1058_14 (.A0(d3[12]), .B0(d4[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[13]), .B1(d4[13]), .C1(GND_net), .D1(GND_net), .CIN(n11041), 
          .COUT(n11042), .S0(d4_71__N_634[12]), .S1(d4_71__N_634[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1058_14.INIT0 = 16'h5666;
    defparam add_1058_14.INIT1 = 16'h5666;
    defparam add_1058_14.INJECT1_0 = "NO";
    defparam add_1058_14.INJECT1_1 = "NO";
    CCU2D add_1058_12 (.A0(d3[10]), .B0(d4[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[11]), .B1(d4[11]), .C1(GND_net), .D1(GND_net), .CIN(n11040), 
          .COUT(n11041), .S0(d4_71__N_634[10]), .S1(d4_71__N_634[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1058_12.INIT0 = 16'h5666;
    defparam add_1058_12.INIT1 = 16'h5666;
    defparam add_1058_12.INJECT1_0 = "NO";
    defparam add_1058_12.INJECT1_1 = "NO";
    CCU2D add_1058_10 (.A0(d3[8]), .B0(d4[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[9]), .B1(d4[9]), .C1(GND_net), .D1(GND_net), .CIN(n11039), 
          .COUT(n11040), .S0(d4_71__N_634[8]), .S1(d4_71__N_634[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1058_10.INIT0 = 16'h5666;
    defparam add_1058_10.INIT1 = 16'h5666;
    defparam add_1058_10.INJECT1_0 = "NO";
    defparam add_1058_10.INJECT1_1 = "NO";
    CCU2D add_1058_8 (.A0(d3[6]), .B0(d4[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[7]), .B1(d4[7]), .C1(GND_net), .D1(GND_net), .CIN(n11038), 
          .COUT(n11039), .S0(d4_71__N_634[6]), .S1(d4_71__N_634[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1058_8.INIT0 = 16'h5666;
    defparam add_1058_8.INIT1 = 16'h5666;
    defparam add_1058_8.INJECT1_0 = "NO";
    defparam add_1058_8.INJECT1_1 = "NO";
    CCU2D add_1058_6 (.A0(d3[4]), .B0(d4[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[5]), .B1(d4[5]), .C1(GND_net), .D1(GND_net), .CIN(n11037), 
          .COUT(n11038), .S0(d4_71__N_634[4]), .S1(d4_71__N_634[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1058_6.INIT0 = 16'h5666;
    defparam add_1058_6.INIT1 = 16'h5666;
    defparam add_1058_6.INJECT1_0 = "NO";
    defparam add_1058_6.INJECT1_1 = "NO";
    CCU2D add_1058_4 (.A0(d3[2]), .B0(d4[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[3]), .B1(d4[3]), .C1(GND_net), .D1(GND_net), .CIN(n11036), 
          .COUT(n11037), .S0(d4_71__N_634[2]), .S1(d4_71__N_634[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1058_4.INIT0 = 16'h5666;
    defparam add_1058_4.INIT1 = 16'h5666;
    defparam add_1058_4.INJECT1_0 = "NO";
    defparam add_1058_4.INJECT1_1 = "NO";
    CCU2D add_1058_2 (.A0(d3[0]), .B0(d4[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[1]), .B1(d4[1]), .C1(GND_net), .D1(GND_net), .COUT(n11036), 
          .S1(d4_71__N_634[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1058_2.INIT0 = 16'h7000;
    defparam add_1058_2.INIT1 = 16'h5666;
    defparam add_1058_2.INJECT1_0 = "NO";
    defparam add_1058_2.INJECT1_1 = "NO";
    CCU2D add_1053_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11034), 
          .S0(n4580));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1053_cout.INIT0 = 16'h0000;
    defparam add_1053_cout.INIT1 = 16'h0000;
    defparam add_1053_cout.INJECT1_0 = "NO";
    defparam add_1053_cout.INJECT1_1 = "NO";
    CCU2D add_1053_36 (.A0(d2[34]), .B0(d3[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[35]), .B1(d3[35]), .C1(GND_net), .D1(GND_net), .CIN(n11033), 
          .COUT(n11034), .S0(d3_71__N_562[34]), .S1(d3_71__N_562[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1053_36.INIT0 = 16'h5666;
    defparam add_1053_36.INIT1 = 16'h5666;
    defparam add_1053_36.INJECT1_0 = "NO";
    defparam add_1053_36.INJECT1_1 = "NO";
    CCU2D add_1053_34 (.A0(d2[32]), .B0(d3[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[33]), .B1(d3[33]), .C1(GND_net), .D1(GND_net), .CIN(n11032), 
          .COUT(n11033), .S0(d3_71__N_562[32]), .S1(d3_71__N_562[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1053_34.INIT0 = 16'h5666;
    defparam add_1053_34.INIT1 = 16'h5666;
    defparam add_1053_34.INJECT1_0 = "NO";
    defparam add_1053_34.INJECT1_1 = "NO";
    CCU2D add_1053_32 (.A0(d2[30]), .B0(d3[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[31]), .B1(d3[31]), .C1(GND_net), .D1(GND_net), .CIN(n11031), 
          .COUT(n11032), .S0(d3_71__N_562[30]), .S1(d3_71__N_562[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1053_32.INIT0 = 16'h5666;
    defparam add_1053_32.INIT1 = 16'h5666;
    defparam add_1053_32.INJECT1_0 = "NO";
    defparam add_1053_32.INJECT1_1 = "NO";
    CCU2D add_1053_30 (.A0(d2[28]), .B0(d3[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[29]), .B1(d3[29]), .C1(GND_net), .D1(GND_net), .CIN(n11030), 
          .COUT(n11031), .S0(d3_71__N_562[28]), .S1(d3_71__N_562[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1053_30.INIT0 = 16'h5666;
    defparam add_1053_30.INIT1 = 16'h5666;
    defparam add_1053_30.INJECT1_0 = "NO";
    defparam add_1053_30.INJECT1_1 = "NO";
    CCU2D add_1053_28 (.A0(d2[26]), .B0(d3[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[27]), .B1(d3[27]), .C1(GND_net), .D1(GND_net), .CIN(n11029), 
          .COUT(n11030), .S0(d3_71__N_562[26]), .S1(d3_71__N_562[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1053_28.INIT0 = 16'h5666;
    defparam add_1053_28.INIT1 = 16'h5666;
    defparam add_1053_28.INJECT1_0 = "NO";
    defparam add_1053_28.INJECT1_1 = "NO";
    CCU2D add_1053_26 (.A0(d2[24]), .B0(d3[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[25]), .B1(d3[25]), .C1(GND_net), .D1(GND_net), .CIN(n11028), 
          .COUT(n11029), .S0(d3_71__N_562[24]), .S1(d3_71__N_562[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1053_26.INIT0 = 16'h5666;
    defparam add_1053_26.INIT1 = 16'h5666;
    defparam add_1053_26.INJECT1_0 = "NO";
    defparam add_1053_26.INJECT1_1 = "NO";
    CCU2D add_1053_24 (.A0(d2[22]), .B0(d3[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[23]), .B1(d3[23]), .C1(GND_net), .D1(GND_net), .CIN(n11027), 
          .COUT(n11028), .S0(d3_71__N_562[22]), .S1(d3_71__N_562[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1053_24.INIT0 = 16'h5666;
    defparam add_1053_24.INIT1 = 16'h5666;
    defparam add_1053_24.INJECT1_0 = "NO";
    defparam add_1053_24.INJECT1_1 = "NO";
    CCU2D add_1053_22 (.A0(d2[20]), .B0(d3[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[21]), .B1(d3[21]), .C1(GND_net), .D1(GND_net), .CIN(n11026), 
          .COUT(n11027), .S0(d3_71__N_562[20]), .S1(d3_71__N_562[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1053_22.INIT0 = 16'h5666;
    defparam add_1053_22.INIT1 = 16'h5666;
    defparam add_1053_22.INJECT1_0 = "NO";
    defparam add_1053_22.INJECT1_1 = "NO";
    CCU2D add_1053_20 (.A0(d2[18]), .B0(d3[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[19]), .B1(d3[19]), .C1(GND_net), .D1(GND_net), .CIN(n11025), 
          .COUT(n11026), .S0(d3_71__N_562[18]), .S1(d3_71__N_562[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1053_20.INIT0 = 16'h5666;
    defparam add_1053_20.INIT1 = 16'h5666;
    defparam add_1053_20.INJECT1_0 = "NO";
    defparam add_1053_20.INJECT1_1 = "NO";
    CCU2D add_1053_18 (.A0(d2[16]), .B0(d3[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[17]), .B1(d3[17]), .C1(GND_net), .D1(GND_net), .CIN(n11024), 
          .COUT(n11025), .S0(d3_71__N_562[16]), .S1(d3_71__N_562[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1053_18.INIT0 = 16'h5666;
    defparam add_1053_18.INIT1 = 16'h5666;
    defparam add_1053_18.INJECT1_0 = "NO";
    defparam add_1053_18.INJECT1_1 = "NO";
    CCU2D add_1053_16 (.A0(d2[14]), .B0(d3[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[15]), .B1(d3[15]), .C1(GND_net), .D1(GND_net), .CIN(n11023), 
          .COUT(n11024), .S0(d3_71__N_562[14]), .S1(d3_71__N_562[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1053_16.INIT0 = 16'h5666;
    defparam add_1053_16.INIT1 = 16'h5666;
    defparam add_1053_16.INJECT1_0 = "NO";
    defparam add_1053_16.INJECT1_1 = "NO";
    CCU2D add_1053_14 (.A0(d2[12]), .B0(d3[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[13]), .B1(d3[13]), .C1(GND_net), .D1(GND_net), .CIN(n11022), 
          .COUT(n11023), .S0(d3_71__N_562[12]), .S1(d3_71__N_562[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1053_14.INIT0 = 16'h5666;
    defparam add_1053_14.INIT1 = 16'h5666;
    defparam add_1053_14.INJECT1_0 = "NO";
    defparam add_1053_14.INJECT1_1 = "NO";
    CCU2D add_1053_12 (.A0(d2[10]), .B0(d3[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[11]), .B1(d3[11]), .C1(GND_net), .D1(GND_net), .CIN(n11021), 
          .COUT(n11022), .S0(d3_71__N_562[10]), .S1(d3_71__N_562[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1053_12.INIT0 = 16'h5666;
    defparam add_1053_12.INIT1 = 16'h5666;
    defparam add_1053_12.INJECT1_0 = "NO";
    defparam add_1053_12.INJECT1_1 = "NO";
    CCU2D add_1053_10 (.A0(d2[8]), .B0(d3[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[9]), .B1(d3[9]), .C1(GND_net), .D1(GND_net), .CIN(n11020), 
          .COUT(n11021), .S0(d3_71__N_562[8]), .S1(d3_71__N_562[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1053_10.INIT0 = 16'h5666;
    defparam add_1053_10.INIT1 = 16'h5666;
    defparam add_1053_10.INJECT1_0 = "NO";
    defparam add_1053_10.INJECT1_1 = "NO";
    CCU2D add_1053_8 (.A0(d2[6]), .B0(d3[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[7]), .B1(d3[7]), .C1(GND_net), .D1(GND_net), .CIN(n11019), 
          .COUT(n11020), .S0(d3_71__N_562[6]), .S1(d3_71__N_562[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1053_8.INIT0 = 16'h5666;
    defparam add_1053_8.INIT1 = 16'h5666;
    defparam add_1053_8.INJECT1_0 = "NO";
    defparam add_1053_8.INJECT1_1 = "NO";
    CCU2D add_1053_6 (.A0(d2[4]), .B0(d3[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[5]), .B1(d3[5]), .C1(GND_net), .D1(GND_net), .CIN(n11018), 
          .COUT(n11019), .S0(d3_71__N_562[4]), .S1(d3_71__N_562[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1053_6.INIT0 = 16'h5666;
    defparam add_1053_6.INIT1 = 16'h5666;
    defparam add_1053_6.INJECT1_0 = "NO";
    defparam add_1053_6.INJECT1_1 = "NO";
    CCU2D add_1053_4 (.A0(d2[2]), .B0(d3[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[3]), .B1(d3[3]), .C1(GND_net), .D1(GND_net), .CIN(n11017), 
          .COUT(n11018), .S0(d3_71__N_562[2]), .S1(d3_71__N_562[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1053_4.INIT0 = 16'h5666;
    defparam add_1053_4.INIT1 = 16'h5666;
    defparam add_1053_4.INJECT1_0 = "NO";
    defparam add_1053_4.INJECT1_1 = "NO";
    CCU2D add_1053_2 (.A0(d2[0]), .B0(d3[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[1]), .B1(d3[1]), .C1(GND_net), .D1(GND_net), .COUT(n11017), 
          .S1(d3_71__N_562[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1053_2.INIT0 = 16'h7000;
    defparam add_1053_2.INIT1 = 16'h5666;
    defparam add_1053_2.INJECT1_0 = "NO";
    defparam add_1053_2.INJECT1_1 = "NO";
    CCU2D add_1048_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11015), 
          .S0(n4428));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1048_cout.INIT0 = 16'h0000;
    defparam add_1048_cout.INIT1 = 16'h0000;
    defparam add_1048_cout.INJECT1_0 = "NO";
    defparam add_1048_cout.INJECT1_1 = "NO";
    CCU2D add_1048_36 (.A0(d1[34]), .B0(d2[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[35]), .B1(d2[35]), .C1(GND_net), .D1(GND_net), .CIN(n11014), 
          .COUT(n11015), .S0(d2_71__N_490[34]), .S1(d2_71__N_490[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1048_36.INIT0 = 16'h5666;
    defparam add_1048_36.INIT1 = 16'h5666;
    defparam add_1048_36.INJECT1_0 = "NO";
    defparam add_1048_36.INJECT1_1 = "NO";
    CCU2D add_1048_34 (.A0(d1[32]), .B0(d2[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[33]), .B1(d2[33]), .C1(GND_net), .D1(GND_net), .CIN(n11013), 
          .COUT(n11014), .S0(d2_71__N_490[32]), .S1(d2_71__N_490[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1048_34.INIT0 = 16'h5666;
    defparam add_1048_34.INIT1 = 16'h5666;
    defparam add_1048_34.INJECT1_0 = "NO";
    defparam add_1048_34.INJECT1_1 = "NO";
    CCU2D add_1048_32 (.A0(d1[30]), .B0(d2[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[31]), .B1(d2[31]), .C1(GND_net), .D1(GND_net), .CIN(n11012), 
          .COUT(n11013), .S0(d2_71__N_490[30]), .S1(d2_71__N_490[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1048_32.INIT0 = 16'h5666;
    defparam add_1048_32.INIT1 = 16'h5666;
    defparam add_1048_32.INJECT1_0 = "NO";
    defparam add_1048_32.INJECT1_1 = "NO";
    CCU2D add_1048_30 (.A0(d1[28]), .B0(d2[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[29]), .B1(d2[29]), .C1(GND_net), .D1(GND_net), .CIN(n11011), 
          .COUT(n11012), .S0(d2_71__N_490[28]), .S1(d2_71__N_490[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1048_30.INIT0 = 16'h5666;
    defparam add_1048_30.INIT1 = 16'h5666;
    defparam add_1048_30.INJECT1_0 = "NO";
    defparam add_1048_30.INJECT1_1 = "NO";
    CCU2D add_1048_28 (.A0(d1[26]), .B0(d2[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[27]), .B1(d2[27]), .C1(GND_net), .D1(GND_net), .CIN(n11010), 
          .COUT(n11011), .S0(d2_71__N_490[26]), .S1(d2_71__N_490[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1048_28.INIT0 = 16'h5666;
    defparam add_1048_28.INIT1 = 16'h5666;
    defparam add_1048_28.INJECT1_0 = "NO";
    defparam add_1048_28.INJECT1_1 = "NO";
    CCU2D add_1048_26 (.A0(d1[24]), .B0(d2[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[25]), .B1(d2[25]), .C1(GND_net), .D1(GND_net), .CIN(n11009), 
          .COUT(n11010), .S0(d2_71__N_490[24]), .S1(d2_71__N_490[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1048_26.INIT0 = 16'h5666;
    defparam add_1048_26.INIT1 = 16'h5666;
    defparam add_1048_26.INJECT1_0 = "NO";
    defparam add_1048_26.INJECT1_1 = "NO";
    CCU2D add_1048_24 (.A0(d1[22]), .B0(d2[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[23]), .B1(d2[23]), .C1(GND_net), .D1(GND_net), .CIN(n11008), 
          .COUT(n11009), .S0(d2_71__N_490[22]), .S1(d2_71__N_490[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1048_24.INIT0 = 16'h5666;
    defparam add_1048_24.INIT1 = 16'h5666;
    defparam add_1048_24.INJECT1_0 = "NO";
    defparam add_1048_24.INJECT1_1 = "NO";
    CCU2D add_1048_22 (.A0(d1[20]), .B0(d2[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[21]), .B1(d2[21]), .C1(GND_net), .D1(GND_net), .CIN(n11007), 
          .COUT(n11008), .S0(d2_71__N_490[20]), .S1(d2_71__N_490[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1048_22.INIT0 = 16'h5666;
    defparam add_1048_22.INIT1 = 16'h5666;
    defparam add_1048_22.INJECT1_0 = "NO";
    defparam add_1048_22.INJECT1_1 = "NO";
    CCU2D add_1048_20 (.A0(d1[18]), .B0(d2[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[19]), .B1(d2[19]), .C1(GND_net), .D1(GND_net), .CIN(n11006), 
          .COUT(n11007), .S0(d2_71__N_490[18]), .S1(d2_71__N_490[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1048_20.INIT0 = 16'h5666;
    defparam add_1048_20.INIT1 = 16'h5666;
    defparam add_1048_20.INJECT1_0 = "NO";
    defparam add_1048_20.INJECT1_1 = "NO";
    CCU2D add_1048_18 (.A0(d1[16]), .B0(d2[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[17]), .B1(d2[17]), .C1(GND_net), .D1(GND_net), .CIN(n11005), 
          .COUT(n11006), .S0(d2_71__N_490[16]), .S1(d2_71__N_490[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1048_18.INIT0 = 16'h5666;
    defparam add_1048_18.INIT1 = 16'h5666;
    defparam add_1048_18.INJECT1_0 = "NO";
    defparam add_1048_18.INJECT1_1 = "NO";
    CCU2D add_1048_16 (.A0(d1[14]), .B0(d2[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[15]), .B1(d2[15]), .C1(GND_net), .D1(GND_net), .CIN(n11004), 
          .COUT(n11005), .S0(d2_71__N_490[14]), .S1(d2_71__N_490[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1048_16.INIT0 = 16'h5666;
    defparam add_1048_16.INIT1 = 16'h5666;
    defparam add_1048_16.INJECT1_0 = "NO";
    defparam add_1048_16.INJECT1_1 = "NO";
    CCU2D add_1048_14 (.A0(d1[12]), .B0(d2[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[13]), .B1(d2[13]), .C1(GND_net), .D1(GND_net), .CIN(n11003), 
          .COUT(n11004), .S0(d2_71__N_490[12]), .S1(d2_71__N_490[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1048_14.INIT0 = 16'h5666;
    defparam add_1048_14.INIT1 = 16'h5666;
    defparam add_1048_14.INJECT1_0 = "NO";
    defparam add_1048_14.INJECT1_1 = "NO";
    CCU2D add_1048_12 (.A0(d1[10]), .B0(d2[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[11]), .B1(d2[11]), .C1(GND_net), .D1(GND_net), .CIN(n11002), 
          .COUT(n11003), .S0(d2_71__N_490[10]), .S1(d2_71__N_490[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1048_12.INIT0 = 16'h5666;
    defparam add_1048_12.INIT1 = 16'h5666;
    defparam add_1048_12.INJECT1_0 = "NO";
    defparam add_1048_12.INJECT1_1 = "NO";
    CCU2D add_1048_10 (.A0(d1[8]), .B0(d2[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[9]), .B1(d2[9]), .C1(GND_net), .D1(GND_net), .CIN(n11001), 
          .COUT(n11002), .S0(d2_71__N_490[8]), .S1(d2_71__N_490[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1048_10.INIT0 = 16'h5666;
    defparam add_1048_10.INIT1 = 16'h5666;
    defparam add_1048_10.INJECT1_0 = "NO";
    defparam add_1048_10.INJECT1_1 = "NO";
    CCU2D add_1048_8 (.A0(d1[6]), .B0(d2[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[7]), .B1(d2[7]), .C1(GND_net), .D1(GND_net), .CIN(n11000), 
          .COUT(n11001), .S0(d2_71__N_490[6]), .S1(d2_71__N_490[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1048_8.INIT0 = 16'h5666;
    defparam add_1048_8.INIT1 = 16'h5666;
    defparam add_1048_8.INJECT1_0 = "NO";
    defparam add_1048_8.INJECT1_1 = "NO";
    CCU2D add_1048_6 (.A0(d1[4]), .B0(d2[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[5]), .B1(d2[5]), .C1(GND_net), .D1(GND_net), .CIN(n10999), 
          .COUT(n11000), .S0(d2_71__N_490[4]), .S1(d2_71__N_490[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1048_6.INIT0 = 16'h5666;
    defparam add_1048_6.INIT1 = 16'h5666;
    defparam add_1048_6.INJECT1_0 = "NO";
    defparam add_1048_6.INJECT1_1 = "NO";
    CCU2D add_1048_4 (.A0(d1[2]), .B0(d2[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[3]), .B1(d2[3]), .C1(GND_net), .D1(GND_net), .CIN(n10998), 
          .COUT(n10999), .S0(d2_71__N_490[2]), .S1(d2_71__N_490[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1048_4.INIT0 = 16'h5666;
    defparam add_1048_4.INIT1 = 16'h5666;
    defparam add_1048_4.INJECT1_0 = "NO";
    defparam add_1048_4.INJECT1_1 = "NO";
    CCU2D add_1048_2 (.A0(d1[0]), .B0(d2[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[1]), .B1(d2[1]), .C1(GND_net), .D1(GND_net), .COUT(n10998), 
          .S1(d2_71__N_490[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1048_2.INIT0 = 16'h7000;
    defparam add_1048_2.INIT1 = 16'h5666;
    defparam add_1048_2.INJECT1_0 = "NO";
    defparam add_1048_2.INJECT1_1 = "NO";
    CCU2D add_1043_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10953), 
          .S0(n4276));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1043_cout.INIT0 = 16'h0000;
    defparam add_1043_cout.INIT1 = 16'h0000;
    defparam add_1043_cout.INJECT1_0 = "NO";
    defparam add_1043_cout.INJECT1_1 = "NO";
    CCU2D add_1043_36 (.A0(MixerOutSin[11]), .B0(d1[34]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[35]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10952), .COUT(n10953), .S0(d1_71__N_418[34]), 
          .S1(d1_71__N_418[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1043_36.INIT0 = 16'h5666;
    defparam add_1043_36.INIT1 = 16'h5666;
    defparam add_1043_36.INJECT1_0 = "NO";
    defparam add_1043_36.INJECT1_1 = "NO";
    CCU2D add_1043_34 (.A0(MixerOutSin[11]), .B0(d1[32]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[33]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10951), .COUT(n10952), .S0(d1_71__N_418[32]), 
          .S1(d1_71__N_418[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1043_34.INIT0 = 16'h5666;
    defparam add_1043_34.INIT1 = 16'h5666;
    defparam add_1043_34.INJECT1_0 = "NO";
    defparam add_1043_34.INJECT1_1 = "NO";
    CCU2D add_1043_32 (.A0(MixerOutSin[11]), .B0(d1[30]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10950), .COUT(n10951), .S0(d1_71__N_418[30]), 
          .S1(d1_71__N_418[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1043_32.INIT0 = 16'h5666;
    defparam add_1043_32.INIT1 = 16'h5666;
    defparam add_1043_32.INJECT1_0 = "NO";
    defparam add_1043_32.INJECT1_1 = "NO";
    CCU2D add_1043_30 (.A0(MixerOutSin[11]), .B0(d1[28]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10949), .COUT(n10950), .S0(d1_71__N_418[28]), 
          .S1(d1_71__N_418[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1043_30.INIT0 = 16'h5666;
    defparam add_1043_30.INIT1 = 16'h5666;
    defparam add_1043_30.INJECT1_0 = "NO";
    defparam add_1043_30.INJECT1_1 = "NO";
    CCU2D add_1043_28 (.A0(MixerOutSin[11]), .B0(d1[26]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10948), .COUT(n10949), .S0(d1_71__N_418[26]), 
          .S1(d1_71__N_418[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1043_28.INIT0 = 16'h5666;
    defparam add_1043_28.INIT1 = 16'h5666;
    defparam add_1043_28.INJECT1_0 = "NO";
    defparam add_1043_28.INJECT1_1 = "NO";
    CCU2D add_1043_26 (.A0(MixerOutSin[11]), .B0(d1[24]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10947), .COUT(n10948), .S0(d1_71__N_418[24]), 
          .S1(d1_71__N_418[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1043_26.INIT0 = 16'h5666;
    defparam add_1043_26.INIT1 = 16'h5666;
    defparam add_1043_26.INJECT1_0 = "NO";
    defparam add_1043_26.INJECT1_1 = "NO";
    CCU2D add_1043_24 (.A0(MixerOutSin[11]), .B0(d1[22]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10946), .COUT(n10947), .S0(d1_71__N_418[22]), 
          .S1(d1_71__N_418[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1043_24.INIT0 = 16'h5666;
    defparam add_1043_24.INIT1 = 16'h5666;
    defparam add_1043_24.INJECT1_0 = "NO";
    defparam add_1043_24.INJECT1_1 = "NO";
    CCU2D add_1043_22 (.A0(MixerOutSin[11]), .B0(d1[20]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10945), .COUT(n10946), .S0(d1_71__N_418[20]), 
          .S1(d1_71__N_418[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1043_22.INIT0 = 16'h5666;
    defparam add_1043_22.INIT1 = 16'h5666;
    defparam add_1043_22.INJECT1_0 = "NO";
    defparam add_1043_22.INJECT1_1 = "NO";
    CCU2D add_1043_20 (.A0(MixerOutSin[11]), .B0(d1[18]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10944), .COUT(n10945), .S0(d1_71__N_418[18]), 
          .S1(d1_71__N_418[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1043_20.INIT0 = 16'h5666;
    defparam add_1043_20.INIT1 = 16'h5666;
    defparam add_1043_20.INJECT1_0 = "NO";
    defparam add_1043_20.INJECT1_1 = "NO";
    CCU2D add_1043_18 (.A0(MixerOutSin[11]), .B0(d1[16]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10943), .COUT(n10944), .S0(d1_71__N_418[16]), 
          .S1(d1_71__N_418[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1043_18.INIT0 = 16'h5666;
    defparam add_1043_18.INIT1 = 16'h5666;
    defparam add_1043_18.INJECT1_0 = "NO";
    defparam add_1043_18.INJECT1_1 = "NO";
    CCU2D add_1043_16 (.A0(MixerOutSin[11]), .B0(d1[14]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10942), .COUT(n10943), .S0(d1_71__N_418[14]), 
          .S1(d1_71__N_418[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1043_16.INIT0 = 16'h5666;
    defparam add_1043_16.INIT1 = 16'h5666;
    defparam add_1043_16.INJECT1_0 = "NO";
    defparam add_1043_16.INJECT1_1 = "NO";
    CCU2D add_1043_14 (.A0(MixerOutSin[11]), .B0(d1[12]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10941), .COUT(n10942), .S0(d1_71__N_418[12]), 
          .S1(d1_71__N_418[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1043_14.INIT0 = 16'h5666;
    defparam add_1043_14.INIT1 = 16'h5666;
    defparam add_1043_14.INJECT1_0 = "NO";
    defparam add_1043_14.INJECT1_1 = "NO";
    CCU2D add_1043_12 (.A0(MixerOutSin[10]), .B0(d1[10]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10940), .COUT(n10941), .S0(d1_71__N_418[10]), 
          .S1(d1_71__N_418[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1043_12.INIT0 = 16'h5666;
    defparam add_1043_12.INIT1 = 16'h5666;
    defparam add_1043_12.INJECT1_0 = "NO";
    defparam add_1043_12.INJECT1_1 = "NO";
    CCU2D add_1043_10 (.A0(MixerOutSin[8]), .B0(d1[8]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[9]), .B1(d1[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10939), .COUT(n10940), .S0(d1_71__N_418[8]), 
          .S1(d1_71__N_418[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1043_10.INIT0 = 16'h5666;
    defparam add_1043_10.INIT1 = 16'h5666;
    defparam add_1043_10.INJECT1_0 = "NO";
    defparam add_1043_10.INJECT1_1 = "NO";
    CCU2D add_1043_8 (.A0(MixerOutSin[6]), .B0(d1[6]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutSin[7]), .B1(d1[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10938), .COUT(n10939), .S0(d1_71__N_418[6]), .S1(d1_71__N_418[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1043_8.INIT0 = 16'h5666;
    defparam add_1043_8.INIT1 = 16'h5666;
    defparam add_1043_8.INJECT1_0 = "NO";
    defparam add_1043_8.INJECT1_1 = "NO";
    CCU2D add_1043_6 (.A0(MixerOutSin[4]), .B0(d1[4]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutSin[5]), .B1(d1[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10937), .COUT(n10938), .S0(d1_71__N_418[4]), .S1(d1_71__N_418[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1043_6.INIT0 = 16'h5666;
    defparam add_1043_6.INIT1 = 16'h5666;
    defparam add_1043_6.INJECT1_0 = "NO";
    defparam add_1043_6.INJECT1_1 = "NO";
    CCU2D add_1043_4 (.A0(MixerOutSin[2]), .B0(d1[2]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutSin[3]), .B1(d1[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10936), .COUT(n10937), .S0(d1_71__N_418[2]), .S1(d1_71__N_418[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1043_4.INIT0 = 16'h5666;
    defparam add_1043_4.INIT1 = 16'h5666;
    defparam add_1043_4.INJECT1_0 = "NO";
    defparam add_1043_4.INJECT1_1 = "NO";
    CCU2D add_1043_2 (.A0(MixerOutSin[0]), .B0(d1[0]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutSin[1]), .B1(d1[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n10936), .S1(d1_71__N_418[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1043_2.INIT0 = 16'h7000;
    defparam add_1043_2.INIT1 = 16'h5666;
    defparam add_1043_2.INJECT1_0 = "NO";
    defparam add_1043_2.INJECT1_1 = "NO";
    CCU2D add_1133_37 (.A0(d6[35]), .B0(d_d6[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n12424), 
          .S0(d7_71__N_1531[35]), .S1(n7012));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1133_37.INIT0 = 16'h5999;
    defparam add_1133_37.INIT1 = 16'h0000;
    defparam add_1133_37.INJECT1_0 = "NO";
    defparam add_1133_37.INJECT1_1 = "NO";
    CCU2D add_1133_35 (.A0(d6[33]), .B0(d_d6[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[34]), .B1(d_d6[34]), .C1(GND_net), .D1(GND_net), .CIN(n12423), 
          .COUT(n12424), .S0(d7_71__N_1531[33]), .S1(d7_71__N_1531[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1133_35.INIT0 = 16'h5999;
    defparam add_1133_35.INIT1 = 16'h5999;
    defparam add_1133_35.INJECT1_0 = "NO";
    defparam add_1133_35.INJECT1_1 = "NO";
    CCU2D add_1133_33 (.A0(d6[31]), .B0(d_d6[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[32]), .B1(d_d6[32]), .C1(GND_net), .D1(GND_net), .CIN(n12422), 
          .COUT(n12423), .S0(d7_71__N_1531[31]), .S1(d7_71__N_1531[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1133_33.INIT0 = 16'h5999;
    defparam add_1133_33.INIT1 = 16'h5999;
    defparam add_1133_33.INJECT1_0 = "NO";
    defparam add_1133_33.INJECT1_1 = "NO";
    CCU2D add_1128_37 (.A0(d7[35]), .B0(d_d7[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11777), 
          .S0(d8_71__N_1603[35]), .S1(n6860));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1128_37.INIT0 = 16'h5999;
    defparam add_1128_37.INIT1 = 16'h0000;
    defparam add_1128_37.INJECT1_0 = "NO";
    defparam add_1128_37.INJECT1_1 = "NO";
    CCU2D add_1128_35 (.A0(d7[33]), .B0(d_d7[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[34]), .B1(d_d7[34]), .C1(GND_net), .D1(GND_net), .CIN(n11776), 
          .COUT(n11777), .S0(d8_71__N_1603[33]), .S1(d8_71__N_1603[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1128_35.INIT0 = 16'h5999;
    defparam add_1128_35.INIT1 = 16'h5999;
    defparam add_1128_35.INJECT1_0 = "NO";
    defparam add_1128_35.INJECT1_1 = "NO";
    CCU2D add_1128_33 (.A0(d7[31]), .B0(d_d7[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[32]), .B1(d_d7[32]), .C1(GND_net), .D1(GND_net), .CIN(n11775), 
          .COUT(n11776), .S0(d8_71__N_1603[31]), .S1(d8_71__N_1603[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1128_33.INIT0 = 16'h5999;
    defparam add_1128_33.INIT1 = 16'h5999;
    defparam add_1128_33.INJECT1_0 = "NO";
    defparam add_1128_33.INJECT1_1 = "NO";
    CCU2D add_1128_31 (.A0(d7[29]), .B0(d_d7[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[30]), .B1(d_d7[30]), .C1(GND_net), .D1(GND_net), .CIN(n11774), 
          .COUT(n11775), .S0(d8_71__N_1603[29]), .S1(d8_71__N_1603[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1128_31.INIT0 = 16'h5999;
    defparam add_1128_31.INIT1 = 16'h5999;
    defparam add_1128_31.INJECT1_0 = "NO";
    defparam add_1128_31.INJECT1_1 = "NO";
    CCU2D add_1128_29 (.A0(d7[27]), .B0(d_d7[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[28]), .B1(d_d7[28]), .C1(GND_net), .D1(GND_net), .CIN(n11773), 
          .COUT(n11774), .S0(d8_71__N_1603[27]), .S1(d8_71__N_1603[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1128_29.INIT0 = 16'h5999;
    defparam add_1128_29.INIT1 = 16'h5999;
    defparam add_1128_29.INJECT1_0 = "NO";
    defparam add_1128_29.INJECT1_1 = "NO";
    CCU2D add_1128_27 (.A0(d7[25]), .B0(d_d7[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[26]), .B1(d_d7[26]), .C1(GND_net), .D1(GND_net), .CIN(n11772), 
          .COUT(n11773), .S0(d8_71__N_1603[25]), .S1(d8_71__N_1603[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1128_27.INIT0 = 16'h5999;
    defparam add_1128_27.INIT1 = 16'h5999;
    defparam add_1128_27.INJECT1_0 = "NO";
    defparam add_1128_27.INJECT1_1 = "NO";
    CCU2D add_1128_25 (.A0(d7[23]), .B0(d_d7[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[24]), .B1(d_d7[24]), .C1(GND_net), .D1(GND_net), .CIN(n11771), 
          .COUT(n11772), .S0(d8_71__N_1603[23]), .S1(d8_71__N_1603[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1128_25.INIT0 = 16'h5999;
    defparam add_1128_25.INIT1 = 16'h5999;
    defparam add_1128_25.INJECT1_0 = "NO";
    defparam add_1128_25.INJECT1_1 = "NO";
    CCU2D add_1128_23 (.A0(d7[21]), .B0(d_d7[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[22]), .B1(d_d7[22]), .C1(GND_net), .D1(GND_net), .CIN(n11770), 
          .COUT(n11771), .S0(d8_71__N_1603[21]), .S1(d8_71__N_1603[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1128_23.INIT0 = 16'h5999;
    defparam add_1128_23.INIT1 = 16'h5999;
    defparam add_1128_23.INJECT1_0 = "NO";
    defparam add_1128_23.INJECT1_1 = "NO";
    CCU2D add_1128_21 (.A0(d7[19]), .B0(d_d7[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[20]), .B1(d_d7[20]), .C1(GND_net), .D1(GND_net), .CIN(n11769), 
          .COUT(n11770), .S0(d8_71__N_1603[19]), .S1(d8_71__N_1603[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1128_21.INIT0 = 16'h5999;
    defparam add_1128_21.INIT1 = 16'h5999;
    defparam add_1128_21.INJECT1_0 = "NO";
    defparam add_1128_21.INJECT1_1 = "NO";
    CCU2D add_1128_19 (.A0(d7[17]), .B0(d_d7[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[18]), .B1(d_d7[18]), .C1(GND_net), .D1(GND_net), .CIN(n11768), 
          .COUT(n11769), .S0(d8_71__N_1603[17]), .S1(d8_71__N_1603[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1128_19.INIT0 = 16'h5999;
    defparam add_1128_19.INIT1 = 16'h5999;
    defparam add_1128_19.INJECT1_0 = "NO";
    defparam add_1128_19.INJECT1_1 = "NO";
    CCU2D add_1128_17 (.A0(d7[15]), .B0(d_d7[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[16]), .B1(d_d7[16]), .C1(GND_net), .D1(GND_net), .CIN(n11767), 
          .COUT(n11768), .S0(d8_71__N_1603[15]), .S1(d8_71__N_1603[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1128_17.INIT0 = 16'h5999;
    defparam add_1128_17.INIT1 = 16'h5999;
    defparam add_1128_17.INJECT1_0 = "NO";
    defparam add_1128_17.INJECT1_1 = "NO";
    CCU2D add_1128_15 (.A0(d7[13]), .B0(d_d7[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[14]), .B1(d_d7[14]), .C1(GND_net), .D1(GND_net), .CIN(n11766), 
          .COUT(n11767), .S0(d8_71__N_1603[13]), .S1(d8_71__N_1603[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1128_15.INIT0 = 16'h5999;
    defparam add_1128_15.INIT1 = 16'h5999;
    defparam add_1128_15.INJECT1_0 = "NO";
    defparam add_1128_15.INJECT1_1 = "NO";
    CCU2D add_1128_13 (.A0(d7[11]), .B0(d_d7[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[12]), .B1(d_d7[12]), .C1(GND_net), .D1(GND_net), .CIN(n11765), 
          .COUT(n11766), .S0(d8_71__N_1603[11]), .S1(d8_71__N_1603[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1128_13.INIT0 = 16'h5999;
    defparam add_1128_13.INIT1 = 16'h5999;
    defparam add_1128_13.INJECT1_0 = "NO";
    defparam add_1128_13.INJECT1_1 = "NO";
    CCU2D add_1128_11 (.A0(d7[9]), .B0(d_d7[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[10]), .B1(d_d7[10]), .C1(GND_net), .D1(GND_net), .CIN(n11764), 
          .COUT(n11765), .S0(d8_71__N_1603[9]), .S1(d8_71__N_1603[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1128_11.INIT0 = 16'h5999;
    defparam add_1128_11.INIT1 = 16'h5999;
    defparam add_1128_11.INJECT1_0 = "NO";
    defparam add_1128_11.INJECT1_1 = "NO";
    CCU2D add_1128_9 (.A0(d7[7]), .B0(d_d7[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[8]), .B1(d_d7[8]), .C1(GND_net), .D1(GND_net), .CIN(n11763), 
          .COUT(n11764), .S0(d8_71__N_1603[7]), .S1(d8_71__N_1603[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1128_9.INIT0 = 16'h5999;
    defparam add_1128_9.INIT1 = 16'h5999;
    defparam add_1128_9.INJECT1_0 = "NO";
    defparam add_1128_9.INJECT1_1 = "NO";
    CCU2D add_1128_7 (.A0(d7[5]), .B0(d_d7[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[6]), .B1(d_d7[6]), .C1(GND_net), .D1(GND_net), .CIN(n11762), 
          .COUT(n11763), .S0(d8_71__N_1603[5]), .S1(d8_71__N_1603[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1128_7.INIT0 = 16'h5999;
    defparam add_1128_7.INIT1 = 16'h5999;
    defparam add_1128_7.INJECT1_0 = "NO";
    defparam add_1128_7.INJECT1_1 = "NO";
    CCU2D add_1128_5 (.A0(d7[3]), .B0(d_d7[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[4]), .B1(d_d7[4]), .C1(GND_net), .D1(GND_net), .CIN(n11761), 
          .COUT(n11762), .S0(d8_71__N_1603[3]), .S1(d8_71__N_1603[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1128_5.INIT0 = 16'h5999;
    defparam add_1128_5.INIT1 = 16'h5999;
    defparam add_1128_5.INJECT1_0 = "NO";
    defparam add_1128_5.INJECT1_1 = "NO";
    CCU2D add_1128_3 (.A0(d7[1]), .B0(d_d7[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[2]), .B1(d_d7[2]), .C1(GND_net), .D1(GND_net), .CIN(n11760), 
          .COUT(n11761), .S0(d8_71__N_1603[1]), .S1(d8_71__N_1603[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1128_3.INIT0 = 16'h5999;
    defparam add_1128_3.INIT1 = 16'h5999;
    defparam add_1128_3.INJECT1_0 = "NO";
    defparam add_1128_3.INJECT1_1 = "NO";
    CCU2D add_1128_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d7[0]), .B1(d_d7[0]), .C1(GND_net), .D1(GND_net), .COUT(n11760), 
          .S1(d8_71__N_1603[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1128_1.INIT0 = 16'h0000;
    defparam add_1128_1.INIT1 = 16'h5999;
    defparam add_1128_1.INJECT1_0 = "NO";
    defparam add_1128_1.INJECT1_1 = "NO";
    CCU2D add_1098_37 (.A0(d9[35]), .B0(d_d9[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11641), 
          .S1(n5948));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1098_37.INIT0 = 16'h5999;
    defparam add_1098_37.INIT1 = 16'h0000;
    defparam add_1098_37.INJECT1_0 = "NO";
    defparam add_1098_37.INJECT1_1 = "NO";
    CCU2D add_1098_35 (.A0(d9[33]), .B0(d_d9[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[34]), .B1(d_d9[34]), .C1(GND_net), .D1(GND_net), .CIN(n11640), 
          .COUT(n11641));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1098_35.INIT0 = 16'h5999;
    defparam add_1098_35.INIT1 = 16'h5999;
    defparam add_1098_35.INJECT1_0 = "NO";
    defparam add_1098_35.INJECT1_1 = "NO";
    CCU2D add_1098_33 (.A0(d9[31]), .B0(d_d9[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[32]), .B1(d_d9[32]), .C1(GND_net), .D1(GND_net), .CIN(n11639), 
          .COUT(n11640));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1098_33.INIT0 = 16'h5999;
    defparam add_1098_33.INIT1 = 16'h5999;
    defparam add_1098_33.INJECT1_0 = "NO";
    defparam add_1098_33.INJECT1_1 = "NO";
    CCU2D add_1098_31 (.A0(d9[29]), .B0(d_d9[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[30]), .B1(d_d9[30]), .C1(GND_net), .D1(GND_net), .CIN(n11638), 
          .COUT(n11639));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1098_31.INIT0 = 16'h5999;
    defparam add_1098_31.INIT1 = 16'h5999;
    defparam add_1098_31.INJECT1_0 = "NO";
    defparam add_1098_31.INJECT1_1 = "NO";
    CCU2D add_1098_29 (.A0(d9[27]), .B0(d_d9[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[28]), .B1(d_d9[28]), .C1(GND_net), .D1(GND_net), .CIN(n11637), 
          .COUT(n11638));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1098_29.INIT0 = 16'h5999;
    defparam add_1098_29.INIT1 = 16'h5999;
    defparam add_1098_29.INJECT1_0 = "NO";
    defparam add_1098_29.INJECT1_1 = "NO";
    CCU2D add_1098_27 (.A0(d9[25]), .B0(d_d9[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[26]), .B1(d_d9[26]), .C1(GND_net), .D1(GND_net), .CIN(n11636), 
          .COUT(n11637));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1098_27.INIT0 = 16'h5999;
    defparam add_1098_27.INIT1 = 16'h5999;
    defparam add_1098_27.INJECT1_0 = "NO";
    defparam add_1098_27.INJECT1_1 = "NO";
    CCU2D add_1098_25 (.A0(d9[23]), .B0(d_d9[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[24]), .B1(d_d9[24]), .C1(GND_net), .D1(GND_net), .CIN(n11635), 
          .COUT(n11636));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1098_25.INIT0 = 16'h5999;
    defparam add_1098_25.INIT1 = 16'h5999;
    defparam add_1098_25.INJECT1_0 = "NO";
    defparam add_1098_25.INJECT1_1 = "NO";
    CCU2D add_1098_23 (.A0(d9[21]), .B0(d_d9[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[22]), .B1(d_d9[22]), .C1(GND_net), .D1(GND_net), .CIN(n11634), 
          .COUT(n11635));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1098_23.INIT0 = 16'h5999;
    defparam add_1098_23.INIT1 = 16'h5999;
    defparam add_1098_23.INJECT1_0 = "NO";
    defparam add_1098_23.INJECT1_1 = "NO";
    CCU2D add_1098_21 (.A0(d9[19]), .B0(d_d9[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[20]), .B1(d_d9[20]), .C1(GND_net), .D1(GND_net), .CIN(n11633), 
          .COUT(n11634));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1098_21.INIT0 = 16'h5999;
    defparam add_1098_21.INIT1 = 16'h5999;
    defparam add_1098_21.INJECT1_0 = "NO";
    defparam add_1098_21.INJECT1_1 = "NO";
    CCU2D add_1098_19 (.A0(d9[17]), .B0(d_d9[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[18]), .B1(d_d9[18]), .C1(GND_net), .D1(GND_net), .CIN(n11632), 
          .COUT(n11633));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1098_19.INIT0 = 16'h5999;
    defparam add_1098_19.INIT1 = 16'h5999;
    defparam add_1098_19.INJECT1_0 = "NO";
    defparam add_1098_19.INJECT1_1 = "NO";
    CCU2D add_1098_17 (.A0(d9[15]), .B0(d_d9[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[16]), .B1(d_d9[16]), .C1(GND_net), .D1(GND_net), .CIN(n11631), 
          .COUT(n11632));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1098_17.INIT0 = 16'h5999;
    defparam add_1098_17.INIT1 = 16'h5999;
    defparam add_1098_17.INJECT1_0 = "NO";
    defparam add_1098_17.INJECT1_1 = "NO";
    CCU2D add_1098_15 (.A0(d9[13]), .B0(d_d9[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[14]), .B1(d_d9[14]), .C1(GND_net), .D1(GND_net), .CIN(n11630), 
          .COUT(n11631));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1098_15.INIT0 = 16'h5999;
    defparam add_1098_15.INIT1 = 16'h5999;
    defparam add_1098_15.INJECT1_0 = "NO";
    defparam add_1098_15.INJECT1_1 = "NO";
    CCU2D add_1098_13 (.A0(d9[11]), .B0(d_d9[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[12]), .B1(d_d9[12]), .C1(GND_net), .D1(GND_net), .CIN(n11629), 
          .COUT(n11630));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1098_13.INIT0 = 16'h5999;
    defparam add_1098_13.INIT1 = 16'h5999;
    defparam add_1098_13.INJECT1_0 = "NO";
    defparam add_1098_13.INJECT1_1 = "NO";
    CCU2D add_1133_31 (.A0(d6[29]), .B0(d_d6[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[30]), .B1(d_d6[30]), .C1(GND_net), .D1(GND_net), .CIN(n12421), 
          .COUT(n12422), .S0(d7_71__N_1531[29]), .S1(d7_71__N_1531[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1133_31.INIT0 = 16'h5999;
    defparam add_1133_31.INIT1 = 16'h5999;
    defparam add_1133_31.INJECT1_0 = "NO";
    defparam add_1133_31.INJECT1_1 = "NO";
    CCU2D add_1133_29 (.A0(d6[27]), .B0(d_d6[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[28]), .B1(d_d6[28]), .C1(GND_net), .D1(GND_net), .CIN(n12420), 
          .COUT(n12421), .S0(d7_71__N_1531[27]), .S1(d7_71__N_1531[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1133_29.INIT0 = 16'h5999;
    defparam add_1133_29.INIT1 = 16'h5999;
    defparam add_1133_29.INJECT1_0 = "NO";
    defparam add_1133_29.INJECT1_1 = "NO";
    CCU2D add_1133_27 (.A0(d6[25]), .B0(d_d6[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[26]), .B1(d_d6[26]), .C1(GND_net), .D1(GND_net), .CIN(n12419), 
          .COUT(n12420), .S0(d7_71__N_1531[25]), .S1(d7_71__N_1531[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1133_27.INIT0 = 16'h5999;
    defparam add_1133_27.INIT1 = 16'h5999;
    defparam add_1133_27.INJECT1_0 = "NO";
    defparam add_1133_27.INJECT1_1 = "NO";
    CCU2D add_1133_25 (.A0(d6[23]), .B0(d_d6[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[24]), .B1(d_d6[24]), .C1(GND_net), .D1(GND_net), .CIN(n12418), 
          .COUT(n12419), .S0(d7_71__N_1531[23]), .S1(d7_71__N_1531[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1133_25.INIT0 = 16'h5999;
    defparam add_1133_25.INIT1 = 16'h5999;
    defparam add_1133_25.INJECT1_0 = "NO";
    defparam add_1133_25.INJECT1_1 = "NO";
    LUT4 shift_right_31_i70_3_lut (.A(d10[69]), .B(d10[70]), .C(\CICGain[0] ), 
         .Z(n70_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i70_3_lut.init = 16'hcaca;
    LUT4 i4_4_lut (.A(n7), .B(count[15]), .C(count[11]), .D(count[14]), 
         .Z(n12793)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i4_4_lut.init = 16'hffef;
    CCU2D add_1133_23 (.A0(d6[21]), .B0(d_d6[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[22]), .B1(d_d6[22]), .C1(GND_net), .D1(GND_net), .CIN(n12417), 
          .COUT(n12418), .S0(d7_71__N_1531[21]), .S1(d7_71__N_1531[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1133_23.INIT0 = 16'h5999;
    defparam add_1133_23.INIT1 = 16'h5999;
    defparam add_1133_23.INJECT1_0 = "NO";
    defparam add_1133_23.INJECT1_1 = "NO";
    CCU2D add_1133_21 (.A0(d6[19]), .B0(d_d6[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[20]), .B1(d_d6[20]), .C1(GND_net), .D1(GND_net), .CIN(n12416), 
          .COUT(n12417), .S0(d7_71__N_1531[19]), .S1(d7_71__N_1531[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1133_21.INIT0 = 16'h5999;
    defparam add_1133_21.INIT1 = 16'h5999;
    defparam add_1133_21.INJECT1_0 = "NO";
    defparam add_1133_21.INJECT1_1 = "NO";
    CCU2D add_1133_19 (.A0(d6[17]), .B0(d_d6[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[18]), .B1(d_d6[18]), .C1(GND_net), .D1(GND_net), .CIN(n12415), 
          .COUT(n12416), .S0(d7_71__N_1531[17]), .S1(d7_71__N_1531[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1133_19.INIT0 = 16'h5999;
    defparam add_1133_19.INIT1 = 16'h5999;
    defparam add_1133_19.INJECT1_0 = "NO";
    defparam add_1133_19.INJECT1_1 = "NO";
    CCU2D add_1133_17 (.A0(d6[15]), .B0(d_d6[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[16]), .B1(d_d6[16]), .C1(GND_net), .D1(GND_net), .CIN(n12414), 
          .COUT(n12415), .S0(d7_71__N_1531[15]), .S1(d7_71__N_1531[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1133_17.INIT0 = 16'h5999;
    defparam add_1133_17.INIT1 = 16'h5999;
    defparam add_1133_17.INJECT1_0 = "NO";
    defparam add_1133_17.INJECT1_1 = "NO";
    CCU2D add_1133_15 (.A0(d6[13]), .B0(d_d6[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[14]), .B1(d_d6[14]), .C1(GND_net), .D1(GND_net), .CIN(n12413), 
          .COUT(n12414), .S0(d7_71__N_1531[13]), .S1(d7_71__N_1531[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1133_15.INIT0 = 16'h5999;
    defparam add_1133_15.INIT1 = 16'h5999;
    defparam add_1133_15.INJECT1_0 = "NO";
    defparam add_1133_15.INJECT1_1 = "NO";
    CCU2D add_1133_13 (.A0(d6[11]), .B0(d_d6[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[12]), .B1(d_d6[12]), .C1(GND_net), .D1(GND_net), .CIN(n12412), 
          .COUT(n12413), .S0(d7_71__N_1531[11]), .S1(d7_71__N_1531[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1133_13.INIT0 = 16'h5999;
    defparam add_1133_13.INIT1 = 16'h5999;
    defparam add_1133_13.INJECT1_0 = "NO";
    defparam add_1133_13.INJECT1_1 = "NO";
    CCU2D add_1133_11 (.A0(d6[9]), .B0(d_d6[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[10]), .B1(d_d6[10]), .C1(GND_net), .D1(GND_net), .CIN(n12411), 
          .COUT(n12412), .S0(d7_71__N_1531[9]), .S1(d7_71__N_1531[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1133_11.INIT0 = 16'h5999;
    defparam add_1133_11.INIT1 = 16'h5999;
    defparam add_1133_11.INJECT1_0 = "NO";
    defparam add_1133_11.INJECT1_1 = "NO";
    CCU2D add_1133_9 (.A0(d6[7]), .B0(d_d6[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[8]), .B1(d_d6[8]), .C1(GND_net), .D1(GND_net), .CIN(n12410), 
          .COUT(n12411), .S0(d7_71__N_1531[7]), .S1(d7_71__N_1531[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1133_9.INIT0 = 16'h5999;
    defparam add_1133_9.INIT1 = 16'h5999;
    defparam add_1133_9.INJECT1_0 = "NO";
    defparam add_1133_9.INJECT1_1 = "NO";
    CCU2D add_1133_7 (.A0(d6[5]), .B0(d_d6[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[6]), .B1(d_d6[6]), .C1(GND_net), .D1(GND_net), .CIN(n12409), 
          .COUT(n12410), .S0(d7_71__N_1531[5]), .S1(d7_71__N_1531[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1133_7.INIT0 = 16'h5999;
    defparam add_1133_7.INIT1 = 16'h5999;
    defparam add_1133_7.INJECT1_0 = "NO";
    defparam add_1133_7.INJECT1_1 = "NO";
    CCU2D add_1133_5 (.A0(d6[3]), .B0(d_d6[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[4]), .B1(d_d6[4]), .C1(GND_net), .D1(GND_net), .CIN(n12408), 
          .COUT(n12409), .S0(d7_71__N_1531[3]), .S1(d7_71__N_1531[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1133_5.INIT0 = 16'h5999;
    defparam add_1133_5.INIT1 = 16'h5999;
    defparam add_1133_5.INJECT1_0 = "NO";
    defparam add_1133_5.INJECT1_1 = "NO";
    CCU2D add_1133_3 (.A0(d6[1]), .B0(d_d6[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[2]), .B1(d_d6[2]), .C1(GND_net), .D1(GND_net), .CIN(n12407), 
          .COUT(n12408), .S0(d7_71__N_1531[1]), .S1(d7_71__N_1531[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1133_3.INIT0 = 16'h5999;
    defparam add_1133_3.INIT1 = 16'h5999;
    defparam add_1133_3.INJECT1_0 = "NO";
    defparam add_1133_3.INJECT1_1 = "NO";
    CCU2D add_1133_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d6[0]), .B1(d_d6[0]), .C1(GND_net), .D1(GND_net), .COUT(n12407), 
          .S1(d7_71__N_1531[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1133_1.INIT0 = 16'h0000;
    defparam add_1133_1.INIT1 = 16'h5999;
    defparam add_1133_1.INJECT1_0 = "NO";
    defparam add_1133_1.INJECT1_1 = "NO";
    CCU2D add_1054_32 (.A0(d2[66]), .B0(d3[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[67]), .B1(d3[67]), .C1(GND_net), .D1(GND_net), .CIN(n12205), 
          .COUT(n12206), .S0(n4581[30]), .S1(n4581[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1054_32.INIT0 = 16'h5666;
    defparam add_1054_32.INIT1 = 16'h5666;
    defparam add_1054_32.INJECT1_0 = "NO";
    defparam add_1054_32.INJECT1_1 = "NO";
    CCU2D add_1054_30 (.A0(d2[64]), .B0(d3[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[65]), .B1(d3[65]), .C1(GND_net), .D1(GND_net), .CIN(n12204), 
          .COUT(n12205), .S0(n4581[28]), .S1(n4581[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1054_30.INIT0 = 16'h5666;
    defparam add_1054_30.INIT1 = 16'h5666;
    defparam add_1054_30.INJECT1_0 = "NO";
    defparam add_1054_30.INJECT1_1 = "NO";
    CCU2D add_1054_28 (.A0(d2[62]), .B0(d3[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[63]), .B1(d3[63]), .C1(GND_net), .D1(GND_net), .CIN(n12203), 
          .COUT(n12204), .S0(n4581[26]), .S1(n4581[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1054_28.INIT0 = 16'h5666;
    defparam add_1054_28.INIT1 = 16'h5666;
    defparam add_1054_28.INJECT1_0 = "NO";
    defparam add_1054_28.INJECT1_1 = "NO";
    LUT4 i2905_2_lut (.A(n375[11]), .B(n31), .Z(count_15__N_1442[11])) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(86[13] 89[16])
    defparam i2905_2_lut.init = 16'hbbbb;
    LUT4 i2_2_lut (.A(count[13]), .B(count[12]), .Z(n7)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i5706_2_lut (.A(n31), .B(n13505), .Z(n8376)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam i5706_2_lut.init = 16'hdddd;
    CCU2D add_1054_26 (.A0(d2[60]), .B0(d3[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[61]), .B1(d3[61]), .C1(GND_net), .D1(GND_net), .CIN(n12202), 
          .COUT(n12203), .S0(n4581[24]), .S1(n4581[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1054_26.INIT0 = 16'h5666;
    defparam add_1054_26.INIT1 = 16'h5666;
    defparam add_1054_26.INJECT1_0 = "NO";
    defparam add_1054_26.INJECT1_1 = "NO";
    CCU2D add_1054_24 (.A0(d2[58]), .B0(d3[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[59]), .B1(d3[59]), .C1(GND_net), .D1(GND_net), .CIN(n12201), 
          .COUT(n12202), .S0(n4581[22]), .S1(n4581[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1054_24.INIT0 = 16'h5666;
    defparam add_1054_24.INIT1 = 16'h5666;
    defparam add_1054_24.INJECT1_0 = "NO";
    defparam add_1054_24.INJECT1_1 = "NO";
    CCU2D add_1054_22 (.A0(d2[56]), .B0(d3[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[57]), .B1(d3[57]), .C1(GND_net), .D1(GND_net), .CIN(n12200), 
          .COUT(n12201), .S0(n4581[20]), .S1(n4581[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1054_22.INIT0 = 16'h5666;
    defparam add_1054_22.INIT1 = 16'h5666;
    defparam add_1054_22.INJECT1_0 = "NO";
    defparam add_1054_22.INJECT1_1 = "NO";
    CCU2D add_1054_20 (.A0(d2[54]), .B0(d3[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[55]), .B1(d3[55]), .C1(GND_net), .D1(GND_net), .CIN(n12199), 
          .COUT(n12200), .S0(n4581[18]), .S1(n4581[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1054_20.INIT0 = 16'h5666;
    defparam add_1054_20.INIT1 = 16'h5666;
    defparam add_1054_20.INJECT1_0 = "NO";
    defparam add_1054_20.INJECT1_1 = "NO";
    CCU2D add_1054_18 (.A0(d2[52]), .B0(d3[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[53]), .B1(d3[53]), .C1(GND_net), .D1(GND_net), .CIN(n12198), 
          .COUT(n12199), .S0(n4581[16]), .S1(n4581[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1054_18.INIT0 = 16'h5666;
    defparam add_1054_18.INIT1 = 16'h5666;
    defparam add_1054_18.INJECT1_0 = "NO";
    defparam add_1054_18.INJECT1_1 = "NO";
    CCU2D add_1054_16 (.A0(d2[50]), .B0(d3[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[51]), .B1(d3[51]), .C1(GND_net), .D1(GND_net), .CIN(n12197), 
          .COUT(n12198), .S0(n4581[14]), .S1(n4581[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1054_16.INIT0 = 16'h5666;
    defparam add_1054_16.INIT1 = 16'h5666;
    defparam add_1054_16.INJECT1_0 = "NO";
    defparam add_1054_16.INJECT1_1 = "NO";
    CCU2D add_1054_14 (.A0(d2[48]), .B0(d3[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[49]), .B1(d3[49]), .C1(GND_net), .D1(GND_net), .CIN(n12196), 
          .COUT(n12197), .S0(n4581[12]), .S1(n4581[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1054_14.INIT0 = 16'h5666;
    defparam add_1054_14.INIT1 = 16'h5666;
    defparam add_1054_14.INJECT1_0 = "NO";
    defparam add_1054_14.INJECT1_1 = "NO";
    CCU2D add_1054_12 (.A0(d2[46]), .B0(d3[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[47]), .B1(d3[47]), .C1(GND_net), .D1(GND_net), .CIN(n12195), 
          .COUT(n12196), .S0(n4581[10]), .S1(n4581[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1054_12.INIT0 = 16'h5666;
    defparam add_1054_12.INIT1 = 16'h5666;
    defparam add_1054_12.INJECT1_0 = "NO";
    defparam add_1054_12.INJECT1_1 = "NO";
    CCU2D add_1054_10 (.A0(d2[44]), .B0(d3[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[45]), .B1(d3[45]), .C1(GND_net), .D1(GND_net), .CIN(n12194), 
          .COUT(n12195), .S0(n4581[8]), .S1(n4581[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1054_10.INIT0 = 16'h5666;
    defparam add_1054_10.INIT1 = 16'h5666;
    defparam add_1054_10.INJECT1_0 = "NO";
    defparam add_1054_10.INJECT1_1 = "NO";
    CCU2D add_1054_8 (.A0(d2[42]), .B0(d3[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[43]), .B1(d3[43]), .C1(GND_net), .D1(GND_net), .CIN(n12193), 
          .COUT(n12194), .S0(n4581[6]), .S1(n4581[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1054_8.INIT0 = 16'h5666;
    defparam add_1054_8.INIT1 = 16'h5666;
    defparam add_1054_8.INJECT1_0 = "NO";
    defparam add_1054_8.INJECT1_1 = "NO";
    CCU2D add_1054_6 (.A0(d2[40]), .B0(d3[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[41]), .B1(d3[41]), .C1(GND_net), .D1(GND_net), .CIN(n12192), 
          .COUT(n12193), .S0(n4581[4]), .S1(n4581[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1054_6.INIT0 = 16'h5666;
    defparam add_1054_6.INIT1 = 16'h5666;
    defparam add_1054_6.INJECT1_0 = "NO";
    defparam add_1054_6.INJECT1_1 = "NO";
    CCU2D add_1054_4 (.A0(d2[38]), .B0(d3[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[39]), .B1(d3[39]), .C1(GND_net), .D1(GND_net), .CIN(n12191), 
          .COUT(n12192), .S0(n4581[2]), .S1(n4581[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1054_4.INIT0 = 16'h5666;
    defparam add_1054_4.INIT1 = 16'h5666;
    defparam add_1054_4.INJECT1_0 = "NO";
    defparam add_1054_4.INJECT1_1 = "NO";
    CCU2D add_1054_2 (.A0(d2[36]), .B0(d3[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[37]), .B1(d3[37]), .C1(GND_net), .D1(GND_net), .COUT(n12191), 
          .S1(n4581[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1054_2.INIT0 = 16'h7000;
    defparam add_1054_2.INIT1 = 16'h5666;
    defparam add_1054_2.INJECT1_0 = "NO";
    defparam add_1054_2.INJECT1_1 = "NO";
    CCU2D add_1055_37 (.A0(d3[70]), .B0(n4580), .C0(n4581[34]), .D0(d2[70]), 
          .A1(d3[71]), .B1(n4580), .C1(n4581[35]), .D1(d2[71]), .CIN(n12188), 
          .S0(d3_71__N_562[70]), .S1(d3_71__N_562[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1055_37.INIT0 = 16'h74b8;
    defparam add_1055_37.INIT1 = 16'h74b8;
    defparam add_1055_37.INJECT1_0 = "NO";
    defparam add_1055_37.INJECT1_1 = "NO";
    CCU2D add_1055_35 (.A0(d3[68]), .B0(n4580), .C0(n4581[32]), .D0(d2[68]), 
          .A1(d3[69]), .B1(n4580), .C1(n4581[33]), .D1(d2[69]), .CIN(n12187), 
          .COUT(n12188), .S0(d3_71__N_562[68]), .S1(d3_71__N_562[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1055_35.INIT0 = 16'h74b8;
    defparam add_1055_35.INIT1 = 16'h74b8;
    defparam add_1055_35.INJECT1_0 = "NO";
    defparam add_1055_35.INJECT1_1 = "NO";
    CCU2D add_1055_33 (.A0(d3[66]), .B0(n4580), .C0(n4581[30]), .D0(d2[66]), 
          .A1(d3[67]), .B1(n4580), .C1(n4581[31]), .D1(d2[67]), .CIN(n12186), 
          .COUT(n12187), .S0(d3_71__N_562[66]), .S1(d3_71__N_562[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1055_33.INIT0 = 16'h74b8;
    defparam add_1055_33.INIT1 = 16'h74b8;
    defparam add_1055_33.INJECT1_0 = "NO";
    defparam add_1055_33.INJECT1_1 = "NO";
    CCU2D add_1055_31 (.A0(d3[64]), .B0(n4580), .C0(n4581[28]), .D0(d2[64]), 
          .A1(d3[65]), .B1(n4580), .C1(n4581[29]), .D1(d2[65]), .CIN(n12185), 
          .COUT(n12186), .S0(d3_71__N_562[64]), .S1(d3_71__N_562[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1055_31.INIT0 = 16'h74b8;
    defparam add_1055_31.INIT1 = 16'h74b8;
    defparam add_1055_31.INJECT1_0 = "NO";
    defparam add_1055_31.INJECT1_1 = "NO";
    CCU2D add_1055_29 (.A0(d3[62]), .B0(n4580), .C0(n4581[26]), .D0(d2[62]), 
          .A1(d3[63]), .B1(n4580), .C1(n4581[27]), .D1(d2[63]), .CIN(n12184), 
          .COUT(n12185), .S0(d3_71__N_562[62]), .S1(d3_71__N_562[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1055_29.INIT0 = 16'h74b8;
    defparam add_1055_29.INIT1 = 16'h74b8;
    defparam add_1055_29.INJECT1_0 = "NO";
    defparam add_1055_29.INJECT1_1 = "NO";
    CCU2D add_1055_27 (.A0(d3[60]), .B0(n4580), .C0(n4581[24]), .D0(d2[60]), 
          .A1(d3[61]), .B1(n4580), .C1(n4581[25]), .D1(d2[61]), .CIN(n12183), 
          .COUT(n12184), .S0(d3_71__N_562[60]), .S1(d3_71__N_562[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1055_27.INIT0 = 16'h74b8;
    defparam add_1055_27.INIT1 = 16'h74b8;
    defparam add_1055_27.INJECT1_0 = "NO";
    defparam add_1055_27.INJECT1_1 = "NO";
    CCU2D add_1055_25 (.A0(d3[58]), .B0(n4580), .C0(n4581[22]), .D0(d2[58]), 
          .A1(d3[59]), .B1(n4580), .C1(n4581[23]), .D1(d2[59]), .CIN(n12182), 
          .COUT(n12183), .S0(d3_71__N_562[58]), .S1(d3_71__N_562[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1055_25.INIT0 = 16'h74b8;
    defparam add_1055_25.INIT1 = 16'h74b8;
    defparam add_1055_25.INJECT1_0 = "NO";
    defparam add_1055_25.INJECT1_1 = "NO";
    CCU2D add_1055_23 (.A0(d3[56]), .B0(n4580), .C0(n4581[20]), .D0(d2[56]), 
          .A1(d3[57]), .B1(n4580), .C1(n4581[21]), .D1(d2[57]), .CIN(n12181), 
          .COUT(n12182), .S0(d3_71__N_562[56]), .S1(d3_71__N_562[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1055_23.INIT0 = 16'h74b8;
    defparam add_1055_23.INIT1 = 16'h74b8;
    defparam add_1055_23.INJECT1_0 = "NO";
    defparam add_1055_23.INJECT1_1 = "NO";
    CCU2D add_1055_21 (.A0(d3[54]), .B0(n4580), .C0(n4581[18]), .D0(d2[54]), 
          .A1(d3[55]), .B1(n4580), .C1(n4581[19]), .D1(d2[55]), .CIN(n12180), 
          .COUT(n12181), .S0(d3_71__N_562[54]), .S1(d3_71__N_562[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1055_21.INIT0 = 16'h74b8;
    defparam add_1055_21.INIT1 = 16'h74b8;
    defparam add_1055_21.INJECT1_0 = "NO";
    defparam add_1055_21.INJECT1_1 = "NO";
    CCU2D add_1055_19 (.A0(d3[52]), .B0(n4580), .C0(n4581[16]), .D0(d2[52]), 
          .A1(d3[53]), .B1(n4580), .C1(n4581[17]), .D1(d2[53]), .CIN(n12179), 
          .COUT(n12180), .S0(d3_71__N_562[52]), .S1(d3_71__N_562[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1055_19.INIT0 = 16'h74b8;
    defparam add_1055_19.INIT1 = 16'h74b8;
    defparam add_1055_19.INJECT1_0 = "NO";
    defparam add_1055_19.INJECT1_1 = "NO";
    CCU2D add_1055_17 (.A0(d3[50]), .B0(n4580), .C0(n4581[14]), .D0(d2[50]), 
          .A1(d3[51]), .B1(n4580), .C1(n4581[15]), .D1(d2[51]), .CIN(n12178), 
          .COUT(n12179), .S0(d3_71__N_562[50]), .S1(d3_71__N_562[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1055_17.INIT0 = 16'h74b8;
    defparam add_1055_17.INIT1 = 16'h74b8;
    defparam add_1055_17.INJECT1_0 = "NO";
    defparam add_1055_17.INJECT1_1 = "NO";
    CCU2D add_1055_15 (.A0(d3[48]), .B0(n4580), .C0(n4581[12]), .D0(d2[48]), 
          .A1(d3[49]), .B1(n4580), .C1(n4581[13]), .D1(d2[49]), .CIN(n12177), 
          .COUT(n12178), .S0(d3_71__N_562[48]), .S1(d3_71__N_562[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1055_15.INIT0 = 16'h74b8;
    defparam add_1055_15.INIT1 = 16'h74b8;
    defparam add_1055_15.INJECT1_0 = "NO";
    defparam add_1055_15.INJECT1_1 = "NO";
    CCU2D add_1055_13 (.A0(d3[46]), .B0(n4580), .C0(n4581[10]), .D0(d2[46]), 
          .A1(d3[47]), .B1(n4580), .C1(n4581[11]), .D1(d2[47]), .CIN(n12176), 
          .COUT(n12177), .S0(d3_71__N_562[46]), .S1(d3_71__N_562[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1055_13.INIT0 = 16'h74b8;
    defparam add_1055_13.INIT1 = 16'h74b8;
    defparam add_1055_13.INJECT1_0 = "NO";
    defparam add_1055_13.INJECT1_1 = "NO";
    CCU2D add_1055_11 (.A0(d3[44]), .B0(n4580), .C0(n4581[8]), .D0(d2[44]), 
          .A1(d3[45]), .B1(n4580), .C1(n4581[9]), .D1(d2[45]), .CIN(n12175), 
          .COUT(n12176), .S0(d3_71__N_562[44]), .S1(d3_71__N_562[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1055_11.INIT0 = 16'h74b8;
    defparam add_1055_11.INIT1 = 16'h74b8;
    defparam add_1055_11.INJECT1_0 = "NO";
    defparam add_1055_11.INJECT1_1 = "NO";
    CCU2D add_1055_9 (.A0(d3[42]), .B0(n4580), .C0(n4581[6]), .D0(d2[42]), 
          .A1(d3[43]), .B1(n4580), .C1(n4581[7]), .D1(d2[43]), .CIN(n12174), 
          .COUT(n12175), .S0(d3_71__N_562[42]), .S1(d3_71__N_562[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1055_9.INIT0 = 16'h74b8;
    defparam add_1055_9.INIT1 = 16'h74b8;
    defparam add_1055_9.INJECT1_0 = "NO";
    defparam add_1055_9.INJECT1_1 = "NO";
    CCU2D add_1055_7 (.A0(d3[40]), .B0(n4580), .C0(n4581[4]), .D0(d2[40]), 
          .A1(d3[41]), .B1(n4580), .C1(n4581[5]), .D1(d2[41]), .CIN(n12173), 
          .COUT(n12174), .S0(d3_71__N_562[40]), .S1(d3_71__N_562[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1055_7.INIT0 = 16'h74b8;
    defparam add_1055_7.INIT1 = 16'h74b8;
    defparam add_1055_7.INJECT1_0 = "NO";
    defparam add_1055_7.INJECT1_1 = "NO";
    CCU2D add_1055_5 (.A0(d3[38]), .B0(n4580), .C0(n4581[2]), .D0(d2[38]), 
          .A1(d3[39]), .B1(n4580), .C1(n4581[3]), .D1(d2[39]), .CIN(n12172), 
          .COUT(n12173), .S0(d3_71__N_562[38]), .S1(d3_71__N_562[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1055_5.INIT0 = 16'h74b8;
    defparam add_1055_5.INIT1 = 16'h74b8;
    defparam add_1055_5.INJECT1_0 = "NO";
    defparam add_1055_5.INJECT1_1 = "NO";
    CCU2D add_1055_3 (.A0(d3[36]), .B0(n4580), .C0(n4581[0]), .D0(d2[36]), 
          .A1(d3[37]), .B1(n4580), .C1(n4581[1]), .D1(d2[37]), .CIN(n12171), 
          .COUT(n12172), .S0(d3_71__N_562[36]), .S1(d3_71__N_562[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1055_3.INIT0 = 16'h74b8;
    defparam add_1055_3.INIT1 = 16'h74b8;
    defparam add_1055_3.INJECT1_0 = "NO";
    defparam add_1055_3.INJECT1_1 = "NO";
    CCU2D add_1055_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n4580), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n12171));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1055_1.INIT0 = 16'hF000;
    defparam add_1055_1.INIT1 = 16'h0555;
    defparam add_1055_1.INJECT1_0 = "NO";
    defparam add_1055_1.INJECT1_1 = "NO";
    CCU2D add_1059_36 (.A0(d3[70]), .B0(d4[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[71]), .B1(d4[71]), .C1(GND_net), .D1(GND_net), .CIN(n12166), 
          .S0(n4733[34]), .S1(n4733[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1059_36.INIT0 = 16'h5666;
    defparam add_1059_36.INIT1 = 16'h5666;
    defparam add_1059_36.INJECT1_0 = "NO";
    defparam add_1059_36.INJECT1_1 = "NO";
    CCU2D add_1059_34 (.A0(d3[68]), .B0(d4[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[69]), .B1(d4[69]), .C1(GND_net), .D1(GND_net), .CIN(n12165), 
          .COUT(n12166), .S0(n4733[32]), .S1(n4733[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1059_34.INIT0 = 16'h5666;
    defparam add_1059_34.INIT1 = 16'h5666;
    defparam add_1059_34.INJECT1_0 = "NO";
    defparam add_1059_34.INJECT1_1 = "NO";
    CCU2D add_1059_32 (.A0(d3[66]), .B0(d4[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[67]), .B1(d4[67]), .C1(GND_net), .D1(GND_net), .CIN(n12164), 
          .COUT(n12165), .S0(n4733[30]), .S1(n4733[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1059_32.INIT0 = 16'h5666;
    defparam add_1059_32.INIT1 = 16'h5666;
    defparam add_1059_32.INJECT1_0 = "NO";
    defparam add_1059_32.INJECT1_1 = "NO";
    CCU2D add_1059_30 (.A0(d3[64]), .B0(d4[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[65]), .B1(d4[65]), .C1(GND_net), .D1(GND_net), .CIN(n12163), 
          .COUT(n12164), .S0(n4733[28]), .S1(n4733[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1059_30.INIT0 = 16'h5666;
    defparam add_1059_30.INIT1 = 16'h5666;
    defparam add_1059_30.INJECT1_0 = "NO";
    defparam add_1059_30.INJECT1_1 = "NO";
    CCU2D add_1059_28 (.A0(d3[62]), .B0(d4[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[63]), .B1(d4[63]), .C1(GND_net), .D1(GND_net), .CIN(n12162), 
          .COUT(n12163), .S0(n4733[26]), .S1(n4733[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1059_28.INIT0 = 16'h5666;
    defparam add_1059_28.INIT1 = 16'h5666;
    defparam add_1059_28.INJECT1_0 = "NO";
    defparam add_1059_28.INJECT1_1 = "NO";
    CCU2D add_1059_26 (.A0(d3[60]), .B0(d4[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[61]), .B1(d4[61]), .C1(GND_net), .D1(GND_net), .CIN(n12161), 
          .COUT(n12162), .S0(n4733[24]), .S1(n4733[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1059_26.INIT0 = 16'h5666;
    defparam add_1059_26.INIT1 = 16'h5666;
    defparam add_1059_26.INJECT1_0 = "NO";
    defparam add_1059_26.INJECT1_1 = "NO";
    CCU2D add_1059_24 (.A0(d3[58]), .B0(d4[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[59]), .B1(d4[59]), .C1(GND_net), .D1(GND_net), .CIN(n12160), 
          .COUT(n12161), .S0(n4733[22]), .S1(n4733[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1059_24.INIT0 = 16'h5666;
    defparam add_1059_24.INIT1 = 16'h5666;
    defparam add_1059_24.INJECT1_0 = "NO";
    defparam add_1059_24.INJECT1_1 = "NO";
    CCU2D add_1059_22 (.A0(d3[56]), .B0(d4[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[57]), .B1(d4[57]), .C1(GND_net), .D1(GND_net), .CIN(n12159), 
          .COUT(n12160), .S0(n4733[20]), .S1(n4733[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1059_22.INIT0 = 16'h5666;
    defparam add_1059_22.INIT1 = 16'h5666;
    defparam add_1059_22.INJECT1_0 = "NO";
    defparam add_1059_22.INJECT1_1 = "NO";
    CCU2D add_1059_20 (.A0(d3[54]), .B0(d4[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[55]), .B1(d4[55]), .C1(GND_net), .D1(GND_net), .CIN(n12158), 
          .COUT(n12159), .S0(n4733[18]), .S1(n4733[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1059_20.INIT0 = 16'h5666;
    defparam add_1059_20.INIT1 = 16'h5666;
    defparam add_1059_20.INJECT1_0 = "NO";
    defparam add_1059_20.INJECT1_1 = "NO";
    CCU2D add_1059_18 (.A0(d3[52]), .B0(d4[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[53]), .B1(d4[53]), .C1(GND_net), .D1(GND_net), .CIN(n12157), 
          .COUT(n12158), .S0(n4733[16]), .S1(n4733[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1059_18.INIT0 = 16'h5666;
    defparam add_1059_18.INIT1 = 16'h5666;
    defparam add_1059_18.INJECT1_0 = "NO";
    defparam add_1059_18.INJECT1_1 = "NO";
    CCU2D add_1059_16 (.A0(d3[50]), .B0(d4[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[51]), .B1(d4[51]), .C1(GND_net), .D1(GND_net), .CIN(n12156), 
          .COUT(n12157), .S0(n4733[14]), .S1(n4733[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1059_16.INIT0 = 16'h5666;
    defparam add_1059_16.INIT1 = 16'h5666;
    defparam add_1059_16.INJECT1_0 = "NO";
    defparam add_1059_16.INJECT1_1 = "NO";
    CCU2D add_1059_14 (.A0(d3[48]), .B0(d4[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[49]), .B1(d4[49]), .C1(GND_net), .D1(GND_net), .CIN(n12155), 
          .COUT(n12156), .S0(n4733[12]), .S1(n4733[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1059_14.INIT0 = 16'h5666;
    defparam add_1059_14.INIT1 = 16'h5666;
    defparam add_1059_14.INJECT1_0 = "NO";
    defparam add_1059_14.INJECT1_1 = "NO";
    CCU2D add_1059_12 (.A0(d3[46]), .B0(d4[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[47]), .B1(d4[47]), .C1(GND_net), .D1(GND_net), .CIN(n12154), 
          .COUT(n12155), .S0(n4733[10]), .S1(n4733[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1059_12.INIT0 = 16'h5666;
    defparam add_1059_12.INIT1 = 16'h5666;
    defparam add_1059_12.INJECT1_0 = "NO";
    defparam add_1059_12.INJECT1_1 = "NO";
    CCU2D add_1059_10 (.A0(d3[44]), .B0(d4[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[45]), .B1(d4[45]), .C1(GND_net), .D1(GND_net), .CIN(n12153), 
          .COUT(n12154), .S0(n4733[8]), .S1(n4733[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1059_10.INIT0 = 16'h5666;
    defparam add_1059_10.INIT1 = 16'h5666;
    defparam add_1059_10.INJECT1_0 = "NO";
    defparam add_1059_10.INJECT1_1 = "NO";
    CCU2D add_1059_8 (.A0(d3[42]), .B0(d4[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[43]), .B1(d4[43]), .C1(GND_net), .D1(GND_net), .CIN(n12152), 
          .COUT(n12153), .S0(n4733[6]), .S1(n4733[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1059_8.INIT0 = 16'h5666;
    defparam add_1059_8.INIT1 = 16'h5666;
    defparam add_1059_8.INJECT1_0 = "NO";
    defparam add_1059_8.INJECT1_1 = "NO";
    CCU2D add_1059_6 (.A0(d3[40]), .B0(d4[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[41]), .B1(d4[41]), .C1(GND_net), .D1(GND_net), .CIN(n12151), 
          .COUT(n12152), .S0(n4733[4]), .S1(n4733[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1059_6.INIT0 = 16'h5666;
    defparam add_1059_6.INIT1 = 16'h5666;
    defparam add_1059_6.INJECT1_0 = "NO";
    defparam add_1059_6.INJECT1_1 = "NO";
    CCU2D add_1059_4 (.A0(d3[38]), .B0(d4[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[39]), .B1(d4[39]), .C1(GND_net), .D1(GND_net), .CIN(n12150), 
          .COUT(n12151), .S0(n4733[2]), .S1(n4733[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1059_4.INIT0 = 16'h5666;
    defparam add_1059_4.INIT1 = 16'h5666;
    defparam add_1059_4.INJECT1_0 = "NO";
    defparam add_1059_4.INJECT1_1 = "NO";
    CCU2D add_1059_2 (.A0(d3[36]), .B0(d4[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[37]), .B1(d4[37]), .C1(GND_net), .D1(GND_net), .COUT(n12150), 
          .S1(n4733[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1059_2.INIT0 = 16'h7000;
    defparam add_1059_2.INIT1 = 16'h5666;
    defparam add_1059_2.INJECT1_0 = "NO";
    defparam add_1059_2.INJECT1_1 = "NO";
    LUT4 i4969_2_lut (.A(MixerOutSin[11]), .B(d1[36]), .Z(n4277[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4969_2_lut.init = 16'h6666;
    FD1S3AX v_comb_66_rep_90 (.D(osc_clk_enable_1458), .CK(osc_clk), .Q(osc_clk_enable_497)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_90.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_89 (.D(osc_clk_enable_1458), .CK(osc_clk), .Q(osc_clk_enable_447)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_89.GSR = "ENABLED";
    LUT4 i5777_else_3_lut (.A(n62_c), .B(\CICGain[1] ), .C(d10[59]), .Z(n13391)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i5777_else_3_lut.init = 16'he2e2;
    LUT4 i5774_then_3_lut (.A(\CICGain[1] ), .B(d10[59]), .C(d10[57]), 
         .Z(n13395)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i5774_then_3_lut.init = 16'he4e4;
    LUT4 i5774_else_3_lut (.A(n61_adj_2521), .B(\CICGain[1] ), .C(d10[58]), 
         .Z(n13394)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i5774_else_3_lut.init = 16'he2e2;
    LUT4 i11_3_lut_4_lut_then_3_lut (.A(\CICGain[0] ), .B(\d10[67] ), .C(\d10[68] ), 
         .Z(n13398)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam i11_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 i11_3_lut_4_lut_else_3_lut (.A(\CICGain[0] ), .B(\d10[69] ), .C(\d10[70] ), 
         .Z(n13397)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam i11_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 i11_3_lut_4_lut_else_3_lut_adj_43 (.A(\CICGain[0] ), .B(d10[69]), 
         .C(d10[70]), .Z(n13400)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam i11_3_lut_4_lut_else_3_lut_adj_43.init = 16'hd8d8;
    LUT4 shift_right_31_i67_3_lut_rep_80 (.A(d10[66]), .B(d10[67]), .C(\CICGain[0] ), 
         .Z(n13488)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i67_3_lut_rep_80.init = 16'hcaca;
    LUT4 i4908_2_lut (.A(d1[0]), .B(d2[0]), .Z(d2_71__N_490[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4908_2_lut.init = 16'h6666;
    LUT4 i5704_4_lut (.A(n13125), .B(n13), .C(n13127), .D(n13113), .Z(d_clk_tmp_N_1831)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i5704_4_lut.init = 16'h2000;
    LUT4 i4909_2_lut (.A(d2[0]), .B(d3[0]), .Z(d3_71__N_562[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4909_2_lut.init = 16'h6666;
    LUT4 i4910_2_lut (.A(d3[0]), .B(d4[0]), .Z(d4_71__N_634[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4910_2_lut.init = 16'h6666;
    LUT4 i4911_2_lut (.A(d4[0]), .B(d5[0]), .Z(d5_71__N_706[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4911_2_lut.init = 16'h6666;
    FD1S3AX v_comb_66_rep_88 (.D(osc_clk_enable_1458), .CK(osc_clk), .Q(osc_clk_enable_397)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_88.GSR = "ENABLED";
    LUT4 i2321_2_lut (.A(n31), .B(d_clk_tmp), .Z(n8356)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam i2321_2_lut.init = 16'h8888;
    CCU2D add_1060_37 (.A0(d4[70]), .B0(n4732), .C0(n4733[34]), .D0(d3[70]), 
          .A1(d4[71]), .B1(n4732), .C1(n4733[35]), .D1(d3[71]), .CIN(n12147), 
          .S0(d4_71__N_634[70]), .S1(d4_71__N_634[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1060_37.INIT0 = 16'h74b8;
    defparam add_1060_37.INIT1 = 16'h74b8;
    defparam add_1060_37.INJECT1_0 = "NO";
    defparam add_1060_37.INJECT1_1 = "NO";
    CCU2D add_1060_35 (.A0(d4[68]), .B0(n4732), .C0(n4733[32]), .D0(d3[68]), 
          .A1(d4[69]), .B1(n4732), .C1(n4733[33]), .D1(d3[69]), .CIN(n12146), 
          .COUT(n12147), .S0(d4_71__N_634[68]), .S1(d4_71__N_634[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1060_35.INIT0 = 16'h74b8;
    defparam add_1060_35.INIT1 = 16'h74b8;
    defparam add_1060_35.INJECT1_0 = "NO";
    defparam add_1060_35.INJECT1_1 = "NO";
    CCU2D add_1039_37 (.A0(d_tmp[71]), .B0(d_d_tmp[71]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12330), .S0(n4125[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1039_37.INIT0 = 16'h5999;
    defparam add_1039_37.INIT1 = 16'h0000;
    defparam add_1039_37.INJECT1_0 = "NO";
    defparam add_1039_37.INJECT1_1 = "NO";
    CCU2D add_1039_35 (.A0(d_tmp[69]), .B0(d_d_tmp[69]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[70]), .B1(d_d_tmp[70]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12329), .COUT(n12330), .S0(n4125[33]), 
          .S1(n4125[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1039_35.INIT0 = 16'h5999;
    defparam add_1039_35.INIT1 = 16'h5999;
    defparam add_1039_35.INJECT1_0 = "NO";
    defparam add_1039_35.INJECT1_1 = "NO";
    CCU2D add_1060_33 (.A0(d4[66]), .B0(n4732), .C0(n4733[30]), .D0(d3[66]), 
          .A1(d4[67]), .B1(n4732), .C1(n4733[31]), .D1(d3[67]), .CIN(n12145), 
          .COUT(n12146), .S0(d4_71__N_634[66]), .S1(d4_71__N_634[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1060_33.INIT0 = 16'h74b8;
    defparam add_1060_33.INIT1 = 16'h74b8;
    defparam add_1060_33.INJECT1_0 = "NO";
    defparam add_1060_33.INJECT1_1 = "NO";
    CCU2D add_1039_33 (.A0(d_tmp[67]), .B0(d_d_tmp[67]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[68]), .B1(d_d_tmp[68]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12328), .COUT(n12329), .S0(n4125[31]), 
          .S1(n4125[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1039_33.INIT0 = 16'h5999;
    defparam add_1039_33.INIT1 = 16'h5999;
    defparam add_1039_33.INJECT1_0 = "NO";
    defparam add_1039_33.INJECT1_1 = "NO";
    CCU2D add_1039_31 (.A0(d_tmp[65]), .B0(d_d_tmp[65]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[66]), .B1(d_d_tmp[66]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12327), .COUT(n12328), .S0(n4125[29]), 
          .S1(n4125[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1039_31.INIT0 = 16'h5999;
    defparam add_1039_31.INIT1 = 16'h5999;
    defparam add_1039_31.INJECT1_0 = "NO";
    defparam add_1039_31.INJECT1_1 = "NO";
    CCU2D add_1039_29 (.A0(d_tmp[63]), .B0(d_d_tmp[63]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[64]), .B1(d_d_tmp[64]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12326), .COUT(n12327), .S0(n4125[27]), 
          .S1(n4125[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1039_29.INIT0 = 16'h5999;
    defparam add_1039_29.INIT1 = 16'h5999;
    defparam add_1039_29.INJECT1_0 = "NO";
    defparam add_1039_29.INJECT1_1 = "NO";
    CCU2D add_1060_31 (.A0(d4[64]), .B0(n4732), .C0(n4733[28]), .D0(d3[64]), 
          .A1(d4[65]), .B1(n4732), .C1(n4733[29]), .D1(d3[65]), .CIN(n12144), 
          .COUT(n12145), .S0(d4_71__N_634[64]), .S1(d4_71__N_634[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1060_31.INIT0 = 16'h74b8;
    defparam add_1060_31.INIT1 = 16'h74b8;
    defparam add_1060_31.INJECT1_0 = "NO";
    defparam add_1060_31.INJECT1_1 = "NO";
    CCU2D add_1060_29 (.A0(d4[62]), .B0(n4732), .C0(n4733[26]), .D0(d3[62]), 
          .A1(d4[63]), .B1(n4732), .C1(n4733[27]), .D1(d3[63]), .CIN(n12143), 
          .COUT(n12144), .S0(d4_71__N_634[62]), .S1(d4_71__N_634[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1060_29.INIT0 = 16'h74b8;
    defparam add_1060_29.INIT1 = 16'h74b8;
    defparam add_1060_29.INJECT1_0 = "NO";
    defparam add_1060_29.INJECT1_1 = "NO";
    CCU2D add_1039_27 (.A0(d_tmp[61]), .B0(d_d_tmp[61]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[62]), .B1(d_d_tmp[62]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12325), .COUT(n12326), .S0(n4125[25]), 
          .S1(n4125[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1039_27.INIT0 = 16'h5999;
    defparam add_1039_27.INIT1 = 16'h5999;
    defparam add_1039_27.INJECT1_0 = "NO";
    defparam add_1039_27.INJECT1_1 = "NO";
    CCU2D add_1039_25 (.A0(d_tmp[59]), .B0(d_d_tmp[59]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[60]), .B1(d_d_tmp[60]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12324), .COUT(n12325), .S0(n4125[23]), 
          .S1(n4125[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1039_25.INIT0 = 16'h5999;
    defparam add_1039_25.INIT1 = 16'h5999;
    defparam add_1039_25.INJECT1_0 = "NO";
    defparam add_1039_25.INJECT1_1 = "NO";
    CCU2D add_1039_23 (.A0(d_tmp[57]), .B0(d_d_tmp[57]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[58]), .B1(d_d_tmp[58]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12323), .COUT(n12324), .S0(n4125[21]), 
          .S1(n4125[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1039_23.INIT0 = 16'h5999;
    defparam add_1039_23.INIT1 = 16'h5999;
    defparam add_1039_23.INJECT1_0 = "NO";
    defparam add_1039_23.INJECT1_1 = "NO";
    CCU2D add_1060_27 (.A0(d4[60]), .B0(n4732), .C0(n4733[24]), .D0(d3[60]), 
          .A1(d4[61]), .B1(n4732), .C1(n4733[25]), .D1(d3[61]), .CIN(n12142), 
          .COUT(n12143), .S0(d4_71__N_634[60]), .S1(d4_71__N_634[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1060_27.INIT0 = 16'h74b8;
    defparam add_1060_27.INIT1 = 16'h74b8;
    defparam add_1060_27.INJECT1_0 = "NO";
    defparam add_1060_27.INJECT1_1 = "NO";
    CCU2D add_1039_21 (.A0(d_tmp[55]), .B0(d_d_tmp[55]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[56]), .B1(d_d_tmp[56]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12322), .COUT(n12323), .S0(n4125[19]), 
          .S1(n4125[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1039_21.INIT0 = 16'h5999;
    defparam add_1039_21.INIT1 = 16'h5999;
    defparam add_1039_21.INJECT1_0 = "NO";
    defparam add_1039_21.INJECT1_1 = "NO";
    CCU2D add_1039_19 (.A0(d_tmp[53]), .B0(d_d_tmp[53]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[54]), .B1(d_d_tmp[54]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12321), .COUT(n12322), .S0(n4125[17]), 
          .S1(n4125[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1039_19.INIT0 = 16'h5999;
    defparam add_1039_19.INIT1 = 16'h5999;
    defparam add_1039_19.INJECT1_0 = "NO";
    defparam add_1039_19.INJECT1_1 = "NO";
    CCU2D add_1039_17 (.A0(d_tmp[51]), .B0(d_d_tmp[51]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[52]), .B1(d_d_tmp[52]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12320), .COUT(n12321), .S0(n4125[15]), 
          .S1(n4125[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1039_17.INIT0 = 16'h5999;
    defparam add_1039_17.INIT1 = 16'h5999;
    defparam add_1039_17.INJECT1_0 = "NO";
    defparam add_1039_17.INJECT1_1 = "NO";
    CCU2D add_1060_25 (.A0(d4[58]), .B0(n4732), .C0(n4733[22]), .D0(d3[58]), 
          .A1(d4[59]), .B1(n4732), .C1(n4733[23]), .D1(d3[59]), .CIN(n12141), 
          .COUT(n12142), .S0(d4_71__N_634[58]), .S1(d4_71__N_634[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1060_25.INIT0 = 16'h74b8;
    defparam add_1060_25.INIT1 = 16'h74b8;
    defparam add_1060_25.INJECT1_0 = "NO";
    defparam add_1060_25.INJECT1_1 = "NO";
    CCU2D add_1060_23 (.A0(d4[56]), .B0(n4732), .C0(n4733[20]), .D0(d3[56]), 
          .A1(d4[57]), .B1(n4732), .C1(n4733[21]), .D1(d3[57]), .CIN(n12140), 
          .COUT(n12141), .S0(d4_71__N_634[56]), .S1(d4_71__N_634[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1060_23.INIT0 = 16'h74b8;
    defparam add_1060_23.INIT1 = 16'h74b8;
    defparam add_1060_23.INJECT1_0 = "NO";
    defparam add_1060_23.INJECT1_1 = "NO";
    CCU2D add_1039_15 (.A0(d_tmp[49]), .B0(d_d_tmp[49]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[50]), .B1(d_d_tmp[50]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12319), .COUT(n12320), .S0(n4125[13]), 
          .S1(n4125[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1039_15.INIT0 = 16'h5999;
    defparam add_1039_15.INIT1 = 16'h5999;
    defparam add_1039_15.INJECT1_0 = "NO";
    defparam add_1039_15.INJECT1_1 = "NO";
    CCU2D add_1039_13 (.A0(d_tmp[47]), .B0(d_d_tmp[47]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[48]), .B1(d_d_tmp[48]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12318), .COUT(n12319), .S0(n4125[11]), 
          .S1(n4125[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1039_13.INIT0 = 16'h5999;
    defparam add_1039_13.INIT1 = 16'h5999;
    defparam add_1039_13.INJECT1_0 = "NO";
    defparam add_1039_13.INJECT1_1 = "NO";
    CCU2D add_1039_11 (.A0(d_tmp[45]), .B0(d_d_tmp[45]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[46]), .B1(d_d_tmp[46]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12317), .COUT(n12318), .S0(n4125[9]), 
          .S1(n4125[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1039_11.INIT0 = 16'h5999;
    defparam add_1039_11.INIT1 = 16'h5999;
    defparam add_1039_11.INJECT1_0 = "NO";
    defparam add_1039_11.INJECT1_1 = "NO";
    CCU2D add_1039_9 (.A0(d_tmp[43]), .B0(d_d_tmp[43]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[44]), .B1(d_d_tmp[44]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12316), .COUT(n12317), .S0(n4125[7]), 
          .S1(n4125[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1039_9.INIT0 = 16'h5999;
    defparam add_1039_9.INIT1 = 16'h5999;
    defparam add_1039_9.INJECT1_0 = "NO";
    defparam add_1039_9.INJECT1_1 = "NO";
    CCU2D add_1039_7 (.A0(d_tmp[41]), .B0(d_d_tmp[41]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[42]), .B1(d_d_tmp[42]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12315), .COUT(n12316), .S0(n4125[5]), 
          .S1(n4125[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1039_7.INIT0 = 16'h5999;
    defparam add_1039_7.INIT1 = 16'h5999;
    defparam add_1039_7.INJECT1_0 = "NO";
    defparam add_1039_7.INJECT1_1 = "NO";
    CCU2D add_1039_5 (.A0(d_tmp[39]), .B0(d_d_tmp[39]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[40]), .B1(d_d_tmp[40]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12314), .COUT(n12315), .S0(n4125[3]), 
          .S1(n4125[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1039_5.INIT0 = 16'h5999;
    defparam add_1039_5.INIT1 = 16'h5999;
    defparam add_1039_5.INJECT1_0 = "NO";
    defparam add_1039_5.INJECT1_1 = "NO";
    LUT4 i11_4_lut (.A(n21), .B(n19), .C(n15), .D(n16), .Z(n31)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i11_4_lut.init = 16'hfffe;
    CCU2D add_1039_3 (.A0(d_tmp[37]), .B0(d_d_tmp[37]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[38]), .B1(d_d_tmp[38]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12313), .COUT(n12314), .S0(n4125[1]), 
          .S1(n4125[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1039_3.INIT0 = 16'h5999;
    defparam add_1039_3.INIT1 = 16'h5999;
    defparam add_1039_3.INJECT1_0 = "NO";
    defparam add_1039_3.INJECT1_1 = "NO";
    CCU2D add_1039_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[36]), .B1(d_d_tmp[36]), .C1(GND_net), .D1(GND_net), 
          .COUT(n12313), .S1(n4125[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1039_1.INIT0 = 16'hF000;
    defparam add_1039_1.INIT1 = 16'h5999;
    defparam add_1039_1.INJECT1_0 = "NO";
    defparam add_1039_1.INJECT1_1 = "NO";
    CCU2D add_1040_37 (.A0(d_d_tmp[70]), .B0(n4124), .C0(n4125[34]), .D0(d_tmp[70]), 
          .A1(d_d_tmp[71]), .B1(n4124), .C1(n4125[35]), .D1(d_tmp[71]), 
          .CIN(n12311), .S0(d6_71__N_1459[70]), .S1(d6_71__N_1459[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1040_37.INIT0 = 16'hb874;
    defparam add_1040_37.INIT1 = 16'hb874;
    defparam add_1040_37.INJECT1_0 = "NO";
    defparam add_1040_37.INJECT1_1 = "NO";
    CCU2D add_1040_35 (.A0(d_d_tmp[68]), .B0(n4124), .C0(n4125[32]), .D0(d_tmp[68]), 
          .A1(d_d_tmp[69]), .B1(n4124), .C1(n4125[33]), .D1(d_tmp[69]), 
          .CIN(n12310), .COUT(n12311), .S0(d6_71__N_1459[68]), .S1(d6_71__N_1459[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1040_35.INIT0 = 16'hb874;
    defparam add_1040_35.INIT1 = 16'hb874;
    defparam add_1040_35.INJECT1_0 = "NO";
    defparam add_1040_35.INJECT1_1 = "NO";
    CCU2D add_1040_33 (.A0(d_d_tmp[66]), .B0(n4124), .C0(n4125[30]), .D0(d_tmp[66]), 
          .A1(d_d_tmp[67]), .B1(n4124), .C1(n4125[31]), .D1(d_tmp[67]), 
          .CIN(n12309), .COUT(n12310), .S0(d6_71__N_1459[66]), .S1(d6_71__N_1459[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1040_33.INIT0 = 16'hb874;
    defparam add_1040_33.INIT1 = 16'hb874;
    defparam add_1040_33.INJECT1_0 = "NO";
    defparam add_1040_33.INJECT1_1 = "NO";
    CCU2D add_1040_31 (.A0(d_d_tmp[64]), .B0(n4124), .C0(n4125[28]), .D0(d_tmp[64]), 
          .A1(d_d_tmp[65]), .B1(n4124), .C1(n4125[29]), .D1(d_tmp[65]), 
          .CIN(n12308), .COUT(n12309), .S0(d6_71__N_1459[64]), .S1(d6_71__N_1459[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1040_31.INIT0 = 16'hb874;
    defparam add_1040_31.INIT1 = 16'hb874;
    defparam add_1040_31.INJECT1_0 = "NO";
    defparam add_1040_31.INJECT1_1 = "NO";
    CCU2D add_1040_29 (.A0(d_d_tmp[62]), .B0(n4124), .C0(n4125[26]), .D0(d_tmp[62]), 
          .A1(d_d_tmp[63]), .B1(n4124), .C1(n4125[27]), .D1(d_tmp[63]), 
          .CIN(n12307), .COUT(n12308), .S0(d6_71__N_1459[62]), .S1(d6_71__N_1459[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1040_29.INIT0 = 16'hb874;
    defparam add_1040_29.INIT1 = 16'hb874;
    defparam add_1040_29.INJECT1_0 = "NO";
    defparam add_1040_29.INJECT1_1 = "NO";
    CCU2D add_1040_27 (.A0(d_d_tmp[60]), .B0(n4124), .C0(n4125[24]), .D0(d_tmp[60]), 
          .A1(d_d_tmp[61]), .B1(n4124), .C1(n4125[25]), .D1(d_tmp[61]), 
          .CIN(n12306), .COUT(n12307), .S0(d6_71__N_1459[60]), .S1(d6_71__N_1459[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1040_27.INIT0 = 16'hb874;
    defparam add_1040_27.INIT1 = 16'hb874;
    defparam add_1040_27.INJECT1_0 = "NO";
    defparam add_1040_27.INJECT1_1 = "NO";
    LUT4 i9_4_lut (.A(count[9]), .B(count[3]), .C(count[4]), .D(count[0]), 
         .Z(n21)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i9_4_lut.init = 16'hfffe;
    CCU2D add_1040_25 (.A0(d_d_tmp[58]), .B0(n4124), .C0(n4125[22]), .D0(d_tmp[58]), 
          .A1(d_d_tmp[59]), .B1(n4124), .C1(n4125[23]), .D1(d_tmp[59]), 
          .CIN(n12305), .COUT(n12306), .S0(d6_71__N_1459[58]), .S1(d6_71__N_1459[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1040_25.INIT0 = 16'hb874;
    defparam add_1040_25.INIT1 = 16'hb874;
    defparam add_1040_25.INJECT1_0 = "NO";
    defparam add_1040_25.INJECT1_1 = "NO";
    CCU2D add_1040_23 (.A0(d_d_tmp[56]), .B0(n4124), .C0(n4125[20]), .D0(d_tmp[56]), 
          .A1(d_d_tmp[57]), .B1(n4124), .C1(n4125[21]), .D1(d_tmp[57]), 
          .CIN(n12304), .COUT(n12305), .S0(d6_71__N_1459[56]), .S1(d6_71__N_1459[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1040_23.INIT0 = 16'hb874;
    defparam add_1040_23.INIT1 = 16'hb874;
    defparam add_1040_23.INJECT1_0 = "NO";
    defparam add_1040_23.INJECT1_1 = "NO";
    CCU2D add_1040_21 (.A0(d_d_tmp[54]), .B0(n4124), .C0(n4125[18]), .D0(d_tmp[54]), 
          .A1(d_d_tmp[55]), .B1(n4124), .C1(n4125[19]), .D1(d_tmp[55]), 
          .CIN(n12303), .COUT(n12304), .S0(d6_71__N_1459[54]), .S1(d6_71__N_1459[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1040_21.INIT0 = 16'hb874;
    defparam add_1040_21.INIT1 = 16'hb874;
    defparam add_1040_21.INJECT1_0 = "NO";
    defparam add_1040_21.INJECT1_1 = "NO";
    FD1S3AX v_comb_66_rep_87 (.D(osc_clk_enable_1458), .CK(osc_clk), .Q(osc_clk_enable_347)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_87.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_82 (.D(osc_clk_enable_1458), .CK(osc_clk), .Q(osc_clk_enable_75)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_82.GSR = "ENABLED";
    CCU2D add_1060_21 (.A0(d4[54]), .B0(n4732), .C0(n4733[18]), .D0(d3[54]), 
          .A1(d4[55]), .B1(n4732), .C1(n4733[19]), .D1(d3[55]), .CIN(n12139), 
          .COUT(n12140), .S0(d4_71__N_634[54]), .S1(d4_71__N_634[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1060_21.INIT0 = 16'h74b8;
    defparam add_1060_21.INIT1 = 16'h74b8;
    defparam add_1060_21.INJECT1_0 = "NO";
    defparam add_1060_21.INJECT1_1 = "NO";
    CCU2D add_1040_19 (.A0(d_d_tmp[52]), .B0(n4124), .C0(n4125[16]), .D0(d_tmp[52]), 
          .A1(d_d_tmp[53]), .B1(n4124), .C1(n4125[17]), .D1(d_tmp[53]), 
          .CIN(n12302), .COUT(n12303), .S0(d6_71__N_1459[52]), .S1(d6_71__N_1459[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1040_19.INIT0 = 16'hb874;
    defparam add_1040_19.INIT1 = 16'hb874;
    defparam add_1040_19.INJECT1_0 = "NO";
    defparam add_1040_19.INJECT1_1 = "NO";
    CCU2D add_1040_17 (.A0(d_d_tmp[50]), .B0(n4124), .C0(n4125[14]), .D0(d_tmp[50]), 
          .A1(d_d_tmp[51]), .B1(n4124), .C1(n4125[15]), .D1(d_tmp[51]), 
          .CIN(n12301), .COUT(n12302), .S0(d6_71__N_1459[50]), .S1(d6_71__N_1459[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1040_17.INIT0 = 16'hb874;
    defparam add_1040_17.INIT1 = 16'hb874;
    defparam add_1040_17.INJECT1_0 = "NO";
    defparam add_1040_17.INJECT1_1 = "NO";
    CCU2D add_1040_15 (.A0(d_d_tmp[48]), .B0(n4124), .C0(n4125[12]), .D0(d_tmp[48]), 
          .A1(d_d_tmp[49]), .B1(n4124), .C1(n4125[13]), .D1(d_tmp[49]), 
          .CIN(n12300), .COUT(n12301), .S0(d6_71__N_1459[48]), .S1(d6_71__N_1459[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1040_15.INIT0 = 16'hb874;
    defparam add_1040_15.INIT1 = 16'hb874;
    defparam add_1040_15.INJECT1_0 = "NO";
    defparam add_1040_15.INJECT1_1 = "NO";
    CCU2D add_1040_13 (.A0(d_d_tmp[46]), .B0(n4124), .C0(n4125[10]), .D0(d_tmp[46]), 
          .A1(d_d_tmp[47]), .B1(n4124), .C1(n4125[11]), .D1(d_tmp[47]), 
          .CIN(n12299), .COUT(n12300), .S0(d6_71__N_1459[46]), .S1(d6_71__N_1459[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1040_13.INIT0 = 16'hb874;
    defparam add_1040_13.INIT1 = 16'hb874;
    defparam add_1040_13.INJECT1_0 = "NO";
    defparam add_1040_13.INJECT1_1 = "NO";
    CCU2D add_1040_11 (.A0(d_d_tmp[44]), .B0(n4124), .C0(n4125[8]), .D0(d_tmp[44]), 
          .A1(d_d_tmp[45]), .B1(n4124), .C1(n4125[9]), .D1(d_tmp[45]), 
          .CIN(n12298), .COUT(n12299), .S0(d6_71__N_1459[44]), .S1(d6_71__N_1459[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1040_11.INIT0 = 16'hb874;
    defparam add_1040_11.INIT1 = 16'hb874;
    defparam add_1040_11.INJECT1_0 = "NO";
    defparam add_1040_11.INJECT1_1 = "NO";
    CCU2D add_1040_9 (.A0(d_d_tmp[42]), .B0(n4124), .C0(n4125[6]), .D0(d_tmp[42]), 
          .A1(d_d_tmp[43]), .B1(n4124), .C1(n4125[7]), .D1(d_tmp[43]), 
          .CIN(n12297), .COUT(n12298), .S0(d6_71__N_1459[42]), .S1(d6_71__N_1459[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1040_9.INIT0 = 16'hb874;
    defparam add_1040_9.INIT1 = 16'hb874;
    defparam add_1040_9.INJECT1_0 = "NO";
    defparam add_1040_9.INJECT1_1 = "NO";
    CCU2D add_1060_19 (.A0(d4[52]), .B0(n4732), .C0(n4733[16]), .D0(d3[52]), 
          .A1(d4[53]), .B1(n4732), .C1(n4733[17]), .D1(d3[53]), .CIN(n12138), 
          .COUT(n12139), .S0(d4_71__N_634[52]), .S1(d4_71__N_634[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1060_19.INIT0 = 16'h74b8;
    defparam add_1060_19.INIT1 = 16'h74b8;
    defparam add_1060_19.INJECT1_0 = "NO";
    defparam add_1060_19.INJECT1_1 = "NO";
    CCU2D add_1040_7 (.A0(d_d_tmp[40]), .B0(n4124), .C0(n4125[4]), .D0(d_tmp[40]), 
          .A1(d_d_tmp[41]), .B1(n4124), .C1(n4125[5]), .D1(d_tmp[41]), 
          .CIN(n12296), .COUT(n12297), .S0(d6_71__N_1459[40]), .S1(d6_71__N_1459[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1040_7.INIT0 = 16'hb874;
    defparam add_1040_7.INIT1 = 16'hb874;
    defparam add_1040_7.INJECT1_0 = "NO";
    defparam add_1040_7.INJECT1_1 = "NO";
    CCU2D add_1040_5 (.A0(d_d_tmp[38]), .B0(n4124), .C0(n4125[2]), .D0(d_tmp[38]), 
          .A1(d_d_tmp[39]), .B1(n4124), .C1(n4125[3]), .D1(d_tmp[39]), 
          .CIN(n12295), .COUT(n12296), .S0(d6_71__N_1459[38]), .S1(d6_71__N_1459[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1040_5.INIT0 = 16'hb874;
    defparam add_1040_5.INIT1 = 16'hb874;
    defparam add_1040_5.INJECT1_0 = "NO";
    defparam add_1040_5.INJECT1_1 = "NO";
    CCU2D add_1040_3 (.A0(d_d_tmp[36]), .B0(n4124), .C0(n4125[0]), .D0(d_tmp[36]), 
          .A1(d_d_tmp[37]), .B1(n4124), .C1(n4125[1]), .D1(d_tmp[37]), 
          .CIN(n12294), .COUT(n12295), .S0(d6_71__N_1459[36]), .S1(d6_71__N_1459[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1040_3.INIT0 = 16'hb874;
    defparam add_1040_3.INIT1 = 16'hb874;
    defparam add_1040_3.INJECT1_0 = "NO";
    defparam add_1040_3.INJECT1_1 = "NO";
    CCU2D add_1040_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n4124), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n12294));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1040_1.INIT0 = 16'hF000;
    defparam add_1040_1.INIT1 = 16'h0555;
    defparam add_1040_1.INJECT1_0 = "NO";
    defparam add_1040_1.INJECT1_1 = "NO";
    CCU2D add_1044_36 (.A0(MixerOutSin[11]), .B0(d1[70]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[71]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12289), .S0(n4277[34]), .S1(n4277[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1044_36.INIT0 = 16'h5666;
    defparam add_1044_36.INIT1 = 16'h5666;
    defparam add_1044_36.INJECT1_0 = "NO";
    defparam add_1044_36.INJECT1_1 = "NO";
    CCU2D add_1060_17 (.A0(d4[50]), .B0(n4732), .C0(n4733[14]), .D0(d3[50]), 
          .A1(d4[51]), .B1(n4732), .C1(n4733[15]), .D1(d3[51]), .CIN(n12137), 
          .COUT(n12138), .S0(d4_71__N_634[50]), .S1(d4_71__N_634[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1060_17.INIT0 = 16'h74b8;
    defparam add_1060_17.INIT1 = 16'h74b8;
    defparam add_1060_17.INJECT1_0 = "NO";
    defparam add_1060_17.INJECT1_1 = "NO";
    CCU2D add_1044_34 (.A0(MixerOutSin[11]), .B0(d1[68]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[69]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12288), .COUT(n12289), .S0(n4277[32]), 
          .S1(n4277[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1044_34.INIT0 = 16'h5666;
    defparam add_1044_34.INIT1 = 16'h5666;
    defparam add_1044_34.INJECT1_0 = "NO";
    defparam add_1044_34.INJECT1_1 = "NO";
    CCU2D add_1044_32 (.A0(MixerOutSin[11]), .B0(d1[66]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[67]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12287), .COUT(n12288), .S0(n4277[30]), 
          .S1(n4277[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1044_32.INIT0 = 16'h5666;
    defparam add_1044_32.INIT1 = 16'h5666;
    defparam add_1044_32.INJECT1_0 = "NO";
    defparam add_1044_32.INJECT1_1 = "NO";
    CCU2D add_1044_30 (.A0(MixerOutSin[11]), .B0(d1[64]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[65]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12286), .COUT(n12287), .S0(n4277[28]), 
          .S1(n4277[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1044_30.INIT0 = 16'h5666;
    defparam add_1044_30.INIT1 = 16'h5666;
    defparam add_1044_30.INJECT1_0 = "NO";
    defparam add_1044_30.INJECT1_1 = "NO";
    CCU2D add_1044_28 (.A0(MixerOutSin[11]), .B0(d1[62]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[63]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12285), .COUT(n12286), .S0(n4277[26]), 
          .S1(n4277[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1044_28.INIT0 = 16'h5666;
    defparam add_1044_28.INIT1 = 16'h5666;
    defparam add_1044_28.INJECT1_0 = "NO";
    defparam add_1044_28.INJECT1_1 = "NO";
    CCU2D add_1099_21 (.A0(d9[55]), .B0(d_d9[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[56]), .B1(d_d9[56]), .C1(GND_net), .D1(GND_net), .CIN(n11832), 
          .COUT(n11833));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1099_21.INIT0 = 16'h5999;
    defparam add_1099_21.INIT1 = 16'h5999;
    defparam add_1099_21.INJECT1_0 = "NO";
    defparam add_1099_21.INJECT1_1 = "NO";
    FD1P3AX d_tmp_i0_i0 (.D(d5[0]), .SP(osc_clk_enable_1458), .CK(osc_clk), 
            .Q(d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i0.GSR = "ENABLED";
    CCU2D add_1095_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5796), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11844));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1095_1.INIT0 = 16'hF000;
    defparam add_1095_1.INIT1 = 16'h0555;
    defparam add_1095_1.INJECT1_0 = "NO";
    defparam add_1095_1.INJECT1_1 = "NO";
    CCU2D add_1099_37 (.A0(d9[71]), .B0(d_d9[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11840), 
          .S0(n5949[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1099_37.INIT0 = 16'h5999;
    defparam add_1099_37.INIT1 = 16'h0000;
    defparam add_1099_37.INJECT1_0 = "NO";
    defparam add_1099_37.INJECT1_1 = "NO";
    CCU2D add_1044_26 (.A0(MixerOutSin[11]), .B0(d1[60]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[61]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12284), .COUT(n12285), .S0(n4277[24]), 
          .S1(n4277[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1044_26.INIT0 = 16'h5666;
    defparam add_1044_26.INIT1 = 16'h5666;
    defparam add_1044_26.INJECT1_0 = "NO";
    defparam add_1044_26.INJECT1_1 = "NO";
    CCU2D add_1044_24 (.A0(MixerOutSin[11]), .B0(d1[58]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[59]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12283), .COUT(n12284), .S0(n4277[22]), 
          .S1(n4277[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1044_24.INIT0 = 16'h5666;
    defparam add_1044_24.INIT1 = 16'h5666;
    defparam add_1044_24.INJECT1_0 = "NO";
    defparam add_1044_24.INJECT1_1 = "NO";
    CCU2D add_1044_22 (.A0(MixerOutSin[11]), .B0(d1[56]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[57]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12282), .COUT(n12283), .S0(n4277[20]), 
          .S1(n4277[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1044_22.INIT0 = 16'h5666;
    defparam add_1044_22.INIT1 = 16'h5666;
    defparam add_1044_22.INJECT1_0 = "NO";
    defparam add_1044_22.INJECT1_1 = "NO";
    CCU2D add_1044_20 (.A0(MixerOutSin[11]), .B0(d1[54]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[55]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12281), .COUT(n12282), .S0(n4277[18]), 
          .S1(n4277[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1044_20.INIT0 = 16'h5666;
    defparam add_1044_20.INIT1 = 16'h5666;
    defparam add_1044_20.INJECT1_0 = "NO";
    defparam add_1044_20.INJECT1_1 = "NO";
    CCU2D add_1044_18 (.A0(MixerOutSin[11]), .B0(d1[52]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[53]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12280), .COUT(n12281), .S0(n4277[16]), 
          .S1(n4277[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1044_18.INIT0 = 16'h5666;
    defparam add_1044_18.INIT1 = 16'h5666;
    defparam add_1044_18.INJECT1_0 = "NO";
    defparam add_1044_18.INJECT1_1 = "NO";
    CCU2D add_1044_16 (.A0(MixerOutSin[11]), .B0(d1[50]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[51]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12279), .COUT(n12280), .S0(n4277[14]), 
          .S1(n4277[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1044_16.INIT0 = 16'h5666;
    defparam add_1044_16.INIT1 = 16'h5666;
    defparam add_1044_16.INJECT1_0 = "NO";
    defparam add_1044_16.INJECT1_1 = "NO";
    CCU2D add_1044_14 (.A0(MixerOutSin[11]), .B0(d1[48]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[49]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12278), .COUT(n12279), .S0(n4277[12]), 
          .S1(n4277[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1044_14.INIT0 = 16'h5666;
    defparam add_1044_14.INIT1 = 16'h5666;
    defparam add_1044_14.INJECT1_0 = "NO";
    defparam add_1044_14.INJECT1_1 = "NO";
    CCU2D add_1044_12 (.A0(MixerOutSin[11]), .B0(d1[46]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[47]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12277), .COUT(n12278), .S0(n4277[10]), 
          .S1(n4277[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1044_12.INIT0 = 16'h5666;
    defparam add_1044_12.INIT1 = 16'h5666;
    defparam add_1044_12.INJECT1_0 = "NO";
    defparam add_1044_12.INJECT1_1 = "NO";
    CCU2D add_1044_10 (.A0(MixerOutSin[11]), .B0(d1[44]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[45]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12276), .COUT(n12277), .S0(n4277[8]), 
          .S1(n4277[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1044_10.INIT0 = 16'h5666;
    defparam add_1044_10.INIT1 = 16'h5666;
    defparam add_1044_10.INJECT1_0 = "NO";
    defparam add_1044_10.INJECT1_1 = "NO";
    CCU2D add_1044_8 (.A0(MixerOutSin[11]), .B0(d1[42]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[43]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12275), .COUT(n12276), .S0(n4277[6]), 
          .S1(n4277[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1044_8.INIT0 = 16'h5666;
    defparam add_1044_8.INIT1 = 16'h5666;
    defparam add_1044_8.INJECT1_0 = "NO";
    defparam add_1044_8.INJECT1_1 = "NO";
    CCU2D add_1060_15 (.A0(d4[48]), .B0(n4732), .C0(n4733[12]), .D0(d3[48]), 
          .A1(d4[49]), .B1(n4732), .C1(n4733[13]), .D1(d3[49]), .CIN(n12136), 
          .COUT(n12137), .S0(d4_71__N_634[48]), .S1(d4_71__N_634[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1060_15.INIT0 = 16'h74b8;
    defparam add_1060_15.INIT1 = 16'h74b8;
    defparam add_1060_15.INJECT1_0 = "NO";
    defparam add_1060_15.INJECT1_1 = "NO";
    CCU2D add_1060_13 (.A0(d4[46]), .B0(n4732), .C0(n4733[10]), .D0(d3[46]), 
          .A1(d4[47]), .B1(n4732), .C1(n4733[11]), .D1(d3[47]), .CIN(n12135), 
          .COUT(n12136), .S0(d4_71__N_634[46]), .S1(d4_71__N_634[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1060_13.INIT0 = 16'h74b8;
    defparam add_1060_13.INIT1 = 16'h74b8;
    defparam add_1060_13.INJECT1_0 = "NO";
    defparam add_1060_13.INJECT1_1 = "NO";
    LUT4 i5777_then_3_lut (.A(\CICGain[1] ), .B(d10[60]), .C(d10[58]), 
         .Z(n13392)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i5777_then_3_lut.init = 16'he4e4;
    CCU2D add_1060_11 (.A0(d4[44]), .B0(n4732), .C0(n4733[8]), .D0(d3[44]), 
          .A1(d4[45]), .B1(n4732), .C1(n4733[9]), .D1(d3[45]), .CIN(n12134), 
          .COUT(n12135), .S0(d4_71__N_634[44]), .S1(d4_71__N_634[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1060_11.INIT0 = 16'h74b8;
    defparam add_1060_11.INIT1 = 16'h74b8;
    defparam add_1060_11.INJECT1_0 = "NO";
    defparam add_1060_11.INJECT1_1 = "NO";
    LUT4 i7_4_lut (.A(count[10]), .B(count[1]), .C(count[5]), .D(count[6]), 
         .Z(n19)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i7_4_lut.init = 16'hfffe;
    CCU2D add_1060_9 (.A0(d4[42]), .B0(n4732), .C0(n4733[6]), .D0(d3[42]), 
          .A1(d4[43]), .B1(n4732), .C1(n4733[7]), .D1(d3[43]), .CIN(n12133), 
          .COUT(n12134), .S0(d4_71__N_634[42]), .S1(d4_71__N_634[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1060_9.INIT0 = 16'h74b8;
    defparam add_1060_9.INIT1 = 16'h74b8;
    defparam add_1060_9.INJECT1_0 = "NO";
    defparam add_1060_9.INJECT1_1 = "NO";
    LUT4 i4966_2_lut (.A(d1[36]), .B(d2[36]), .Z(n4429[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4966_2_lut.init = 16'h6666;
    LUT4 i3_2_lut (.A(count[8]), .B(count[7]), .Z(n15)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i4_2_lut (.A(n12793), .B(count[2]), .Z(n16)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i4_2_lut.init = 16'heeee;
    LUT4 i4963_2_lut (.A(d2[36]), .B(d3[36]), .Z(n4581[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4963_2_lut.init = 16'h6666;
    CCU2D add_1060_7 (.A0(d4[40]), .B0(n4732), .C0(n4733[4]), .D0(d3[40]), 
          .A1(d4[41]), .B1(n4732), .C1(n4733[5]), .D1(d3[41]), .CIN(n12132), 
          .COUT(n12133), .S0(d4_71__N_634[40]), .S1(d4_71__N_634[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1060_7.INIT0 = 16'h74b8;
    defparam add_1060_7.INIT1 = 16'h74b8;
    defparam add_1060_7.INJECT1_0 = "NO";
    defparam add_1060_7.INJECT1_1 = "NO";
    LUT4 i5657_4_lut (.A(count[6]), .B(count[1]), .C(count[0]), .D(count[8]), 
         .Z(n13125)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5657_4_lut.init = 16'h8000;
    CCU2D add_1060_5 (.A0(d4[38]), .B0(n4732), .C0(n4733[2]), .D0(d3[38]), 
          .A1(d4[39]), .B1(n4732), .C1(n4733[3]), .D1(d3[39]), .CIN(n12131), 
          .COUT(n12132), .S0(d4_71__N_634[38]), .S1(d4_71__N_634[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1060_5.INIT0 = 16'h74b8;
    defparam add_1060_5.INIT1 = 16'h74b8;
    defparam add_1060_5.INJECT1_0 = "NO";
    defparam add_1060_5.INJECT1_1 = "NO";
    CCU2D add_1060_3 (.A0(d4[36]), .B0(n4732), .C0(n4733[0]), .D0(d3[36]), 
          .A1(d4[37]), .B1(n4732), .C1(n4733[1]), .D1(d3[37]), .CIN(n12130), 
          .COUT(n12131), .S0(d4_71__N_634[36]), .S1(d4_71__N_634[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1060_3.INIT0 = 16'h74b8;
    defparam add_1060_3.INIT1 = 16'h74b8;
    defparam add_1060_3.INJECT1_0 = "NO";
    defparam add_1060_3.INJECT1_1 = "NO";
    LUT4 i1_2_lut (.A(n12793), .B(count[3]), .Z(n13)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut.init = 16'hbbbb;
    CCU2D add_1060_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n4732), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n12130));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1060_1.INIT0 = 16'hF000;
    defparam add_1060_1.INIT1 = 16'h0555;
    defparam add_1060_1.INJECT1_0 = "NO";
    defparam add_1060_1.INJECT1_1 = "NO";
    CCU2D add_1064_36 (.A0(d4[70]), .B0(d5[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[71]), .B1(d5[71]), .C1(GND_net), .D1(GND_net), .CIN(n12125), 
          .S0(n4885[34]), .S1(n4885[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1064_36.INIT0 = 16'h5666;
    defparam add_1064_36.INIT1 = 16'h5666;
    defparam add_1064_36.INJECT1_0 = "NO";
    defparam add_1064_36.INJECT1_1 = "NO";
    CCU2D add_1064_34 (.A0(d4[68]), .B0(d5[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[69]), .B1(d5[69]), .C1(GND_net), .D1(GND_net), .CIN(n12124), 
          .COUT(n12125), .S0(n4885[32]), .S1(n4885[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1064_34.INIT0 = 16'h5666;
    defparam add_1064_34.INIT1 = 16'h5666;
    defparam add_1064_34.INJECT1_0 = "NO";
    defparam add_1064_34.INJECT1_1 = "NO";
    CCU2D add_1064_32 (.A0(d4[66]), .B0(d5[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[67]), .B1(d5[67]), .C1(GND_net), .D1(GND_net), .CIN(n12123), 
          .COUT(n12124), .S0(n4885[30]), .S1(n4885[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1064_32.INIT0 = 16'h5666;
    defparam add_1064_32.INIT1 = 16'h5666;
    defparam add_1064_32.INJECT1_0 = "NO";
    defparam add_1064_32.INJECT1_1 = "NO";
    LUT4 i4960_2_lut (.A(d3[36]), .B(d4[36]), .Z(n4733[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4960_2_lut.init = 16'h6666;
    CCU2D add_1064_30 (.A0(d4[64]), .B0(d5[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[65]), .B1(d5[65]), .C1(GND_net), .D1(GND_net), .CIN(n12122), 
          .COUT(n12123), .S0(n4885[28]), .S1(n4885[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1064_30.INIT0 = 16'h5666;
    defparam add_1064_30.INIT1 = 16'h5666;
    defparam add_1064_30.INJECT1_0 = "NO";
    defparam add_1064_30.INJECT1_1 = "NO";
    FD1S3AX v_comb_66_rep_92 (.D(osc_clk_enable_1458), .CK(osc_clk), .Q(osc_clk_enable_597)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_92.GSR = "ENABLED";
    CCU2D add_1064_28 (.A0(d4[62]), .B0(d5[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[63]), .B1(d5[63]), .C1(GND_net), .D1(GND_net), .CIN(n12121), 
          .COUT(n12122), .S0(n4885[26]), .S1(n4885[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1064_28.INIT0 = 16'h5666;
    defparam add_1064_28.INIT1 = 16'h5666;
    defparam add_1064_28.INJECT1_0 = "NO";
    defparam add_1064_28.INJECT1_1 = "NO";
    CCU2D add_1064_26 (.A0(d4[60]), .B0(d5[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[61]), .B1(d5[61]), .C1(GND_net), .D1(GND_net), .CIN(n12120), 
          .COUT(n12121), .S0(n4885[24]), .S1(n4885[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1064_26.INIT0 = 16'h5666;
    defparam add_1064_26.INIT1 = 16'h5666;
    defparam add_1064_26.INJECT1_0 = "NO";
    defparam add_1064_26.INJECT1_1 = "NO";
    CCU2D add_1064_24 (.A0(d4[58]), .B0(d5[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[59]), .B1(d5[59]), .C1(GND_net), .D1(GND_net), .CIN(n12119), 
          .COUT(n12120), .S0(n4885[22]), .S1(n4885[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1064_24.INIT0 = 16'h5666;
    defparam add_1064_24.INIT1 = 16'h5666;
    defparam add_1064_24.INJECT1_0 = "NO";
    defparam add_1064_24.INJECT1_1 = "NO";
    CCU2D add_1064_22 (.A0(d4[56]), .B0(d5[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[57]), .B1(d5[57]), .C1(GND_net), .D1(GND_net), .CIN(n12118), 
          .COUT(n12119), .S0(n4885[20]), .S1(n4885[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1064_22.INIT0 = 16'h5666;
    defparam add_1064_22.INIT1 = 16'h5666;
    defparam add_1064_22.INJECT1_0 = "NO";
    defparam add_1064_22.INJECT1_1 = "NO";
    CCU2D add_1064_20 (.A0(d4[54]), .B0(d5[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[55]), .B1(d5[55]), .C1(GND_net), .D1(GND_net), .CIN(n12117), 
          .COUT(n12118), .S0(n4885[18]), .S1(n4885[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1064_20.INIT0 = 16'h5666;
    defparam add_1064_20.INIT1 = 16'h5666;
    defparam add_1064_20.INJECT1_0 = "NO";
    defparam add_1064_20.INJECT1_1 = "NO";
    CCU2D add_1064_18 (.A0(d4[52]), .B0(d5[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[53]), .B1(d5[53]), .C1(GND_net), .D1(GND_net), .CIN(n12116), 
          .COUT(n12117), .S0(n4885[16]), .S1(n4885[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1064_18.INIT0 = 16'h5666;
    defparam add_1064_18.INIT1 = 16'h5666;
    defparam add_1064_18.INJECT1_0 = "NO";
    defparam add_1064_18.INJECT1_1 = "NO";
    CCU2D add_1064_16 (.A0(d4[50]), .B0(d5[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[51]), .B1(d5[51]), .C1(GND_net), .D1(GND_net), .CIN(n12115), 
          .COUT(n12116), .S0(n4885[14]), .S1(n4885[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1064_16.INIT0 = 16'h5666;
    defparam add_1064_16.INIT1 = 16'h5666;
    defparam add_1064_16.INJECT1_0 = "NO";
    defparam add_1064_16.INJECT1_1 = "NO";
    CCU2D add_1064_14 (.A0(d4[48]), .B0(d5[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[49]), .B1(d5[49]), .C1(GND_net), .D1(GND_net), .CIN(n12114), 
          .COUT(n12115), .S0(n4885[12]), .S1(n4885[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1064_14.INIT0 = 16'h5666;
    defparam add_1064_14.INIT1 = 16'h5666;
    defparam add_1064_14.INJECT1_0 = "NO";
    defparam add_1064_14.INJECT1_1 = "NO";
    CCU2D add_1064_12 (.A0(d4[46]), .B0(d5[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[47]), .B1(d5[47]), .C1(GND_net), .D1(GND_net), .CIN(n12113), 
          .COUT(n12114), .S0(n4885[10]), .S1(n4885[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1064_12.INIT0 = 16'h5666;
    defparam add_1064_12.INIT1 = 16'h5666;
    defparam add_1064_12.INJECT1_0 = "NO";
    defparam add_1064_12.INJECT1_1 = "NO";
    CCU2D add_1064_10 (.A0(d4[44]), .B0(d5[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[45]), .B1(d5[45]), .C1(GND_net), .D1(GND_net), .CIN(n12112), 
          .COUT(n12113), .S0(n4885[8]), .S1(n4885[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1064_10.INIT0 = 16'h5666;
    defparam add_1064_10.INIT1 = 16'h5666;
    defparam add_1064_10.INJECT1_0 = "NO";
    defparam add_1064_10.INJECT1_1 = "NO";
    CCU2D add_1064_8 (.A0(d4[42]), .B0(d5[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[43]), .B1(d5[43]), .C1(GND_net), .D1(GND_net), .CIN(n12111), 
          .COUT(n12112), .S0(n4885[6]), .S1(n4885[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1064_8.INIT0 = 16'h5666;
    defparam add_1064_8.INIT1 = 16'h5666;
    defparam add_1064_8.INJECT1_0 = "NO";
    defparam add_1064_8.INJECT1_1 = "NO";
    CCU2D add_1064_6 (.A0(d4[40]), .B0(d5[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[41]), .B1(d5[41]), .C1(GND_net), .D1(GND_net), .CIN(n12110), 
          .COUT(n12111), .S0(n4885[4]), .S1(n4885[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1064_6.INIT0 = 16'h5666;
    defparam add_1064_6.INIT1 = 16'h5666;
    defparam add_1064_6.INJECT1_0 = "NO";
    defparam add_1064_6.INJECT1_1 = "NO";
    FD1S3AX v_comb_66_rep_94 (.D(osc_clk_enable_1458), .CK(osc_clk), .Q(osc_clk_enable_697)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_94.GSR = "ENABLED";
    CCU2D add_1064_4 (.A0(d4[38]), .B0(d5[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[39]), .B1(d5[39]), .C1(GND_net), .D1(GND_net), .CIN(n12109), 
          .COUT(n12110), .S0(n4885[2]), .S1(n4885[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1064_4.INIT0 = 16'h5666;
    defparam add_1064_4.INIT1 = 16'h5666;
    defparam add_1064_4.INJECT1_0 = "NO";
    defparam add_1064_4.INJECT1_1 = "NO";
    CCU2D add_1064_2 (.A0(d4[36]), .B0(d5[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[37]), .B1(d5[37]), .C1(GND_net), .D1(GND_net), .COUT(n12109), 
          .S1(n4885[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1064_2.INIT0 = 16'h7000;
    defparam add_1064_2.INIT1 = 16'h5666;
    defparam add_1064_2.INJECT1_0 = "NO";
    defparam add_1064_2.INJECT1_1 = "NO";
    CCU2D add_1044_6 (.A0(MixerOutSin[11]), .B0(d1[40]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[41]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12274), .COUT(n12275), .S0(n4277[4]), 
          .S1(n4277[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1044_6.INIT0 = 16'h5666;
    defparam add_1044_6.INIT1 = 16'h5666;
    defparam add_1044_6.INJECT1_0 = "NO";
    defparam add_1044_6.INJECT1_1 = "NO";
    LUT4 i4957_2_lut (.A(d4[36]), .B(d5[36]), .Z(n4885[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4957_2_lut.init = 16'h6666;
    CCU2D add_1044_4 (.A0(MixerOutSin[11]), .B0(d1[38]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[39]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12273), .COUT(n12274), .S0(n4277[2]), 
          .S1(n4277[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1044_4.INIT0 = 16'h5666;
    defparam add_1044_4.INIT1 = 16'h5666;
    defparam add_1044_4.INJECT1_0 = "NO";
    defparam add_1044_4.INJECT1_1 = "NO";
    CCU2D add_1044_2 (.A0(MixerOutSin[11]), .B0(d1[36]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[37]), .C1(GND_net), 
          .D1(GND_net), .COUT(n12273), .S1(n4277[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1044_2.INIT0 = 16'h7000;
    defparam add_1044_2.INIT1 = 16'h5666;
    defparam add_1044_2.INJECT1_0 = "NO";
    defparam add_1044_2.INJECT1_1 = "NO";
    CCU2D add_1065_37 (.A0(d5[70]), .B0(n4884), .C0(n4885[34]), .D0(d4[70]), 
          .A1(d5[71]), .B1(n4884), .C1(n4885[35]), .D1(d4[71]), .CIN(n12106), 
          .S0(d5_71__N_706[70]), .S1(d5_71__N_706[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1065_37.INIT0 = 16'h74b8;
    defparam add_1065_37.INIT1 = 16'h74b8;
    defparam add_1065_37.INJECT1_0 = "NO";
    defparam add_1065_37.INJECT1_1 = "NO";
    PFUMX i5798 (.BLUT(n13400), .ALUT(n13401), .C0(\CICGain[1] ), .Z(d_out_11__N_1819[10]));
    CCU2D add_1065_35 (.A0(d5[68]), .B0(n4884), .C0(n4885[32]), .D0(d4[68]), 
          .A1(d5[69]), .B1(n4884), .C1(n4885[33]), .D1(d4[69]), .CIN(n12105), 
          .COUT(n12106), .S0(d5_71__N_706[68]), .S1(d5_71__N_706[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1065_35.INIT0 = 16'h74b8;
    defparam add_1065_35.INIT1 = 16'h74b8;
    defparam add_1065_35.INJECT1_0 = "NO";
    defparam add_1065_35.INJECT1_1 = "NO";
    CCU2D add_1065_33 (.A0(d5[66]), .B0(n4884), .C0(n4885[30]), .D0(d4[66]), 
          .A1(d5[67]), .B1(n4884), .C1(n4885[31]), .D1(d4[67]), .CIN(n12104), 
          .COUT(n12105), .S0(d5_71__N_706[66]), .S1(d5_71__N_706[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1065_33.INIT0 = 16'h74b8;
    defparam add_1065_33.INIT1 = 16'h74b8;
    defparam add_1065_33.INJECT1_0 = "NO";
    defparam add_1065_33.INJECT1_1 = "NO";
    CCU2D add_1065_31 (.A0(d5[64]), .B0(n4884), .C0(n4885[28]), .D0(d4[64]), 
          .A1(d5[65]), .B1(n4884), .C1(n4885[29]), .D1(d4[65]), .CIN(n12103), 
          .COUT(n12104), .S0(d5_71__N_706[64]), .S1(d5_71__N_706[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1065_31.INIT0 = 16'h74b8;
    defparam add_1065_31.INIT1 = 16'h74b8;
    defparam add_1065_31.INJECT1_0 = "NO";
    defparam add_1065_31.INJECT1_1 = "NO";
    FD1S3AX v_comb_66_rep_84 (.D(osc_clk_enable_1458), .CK(osc_clk), .Q(osc_clk_enable_197)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_84.GSR = "ENABLED";
    PFUMX i5796 (.BLUT(n13397), .ALUT(n13398), .C0(\CICGain[1] ), .Z(\d_out_11__N_1819[10] ));
    CCU2D add_1065_29 (.A0(d5[62]), .B0(n4884), .C0(n4885[26]), .D0(d4[62]), 
          .A1(d5[63]), .B1(n4884), .C1(n4885[27]), .D1(d4[63]), .CIN(n12102), 
          .COUT(n12103), .S0(d5_71__N_706[62]), .S1(d5_71__N_706[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1065_29.INIT0 = 16'h74b8;
    defparam add_1065_29.INIT1 = 16'h74b8;
    defparam add_1065_29.INJECT1_0 = "NO";
    defparam add_1065_29.INJECT1_1 = "NO";
    CCU2D add_1065_27 (.A0(d5[60]), .B0(n4884), .C0(n4885[24]), .D0(d4[60]), 
          .A1(d5[61]), .B1(n4884), .C1(n4885[25]), .D1(d4[61]), .CIN(n12101), 
          .COUT(n12102), .S0(d5_71__N_706[60]), .S1(d5_71__N_706[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1065_27.INIT0 = 16'h74b8;
    defparam add_1065_27.INIT1 = 16'h74b8;
    defparam add_1065_27.INJECT1_0 = "NO";
    defparam add_1065_27.INJECT1_1 = "NO";
    CCU2D add_1065_25 (.A0(d5[58]), .B0(n4884), .C0(n4885[22]), .D0(d4[58]), 
          .A1(d5[59]), .B1(n4884), .C1(n4885[23]), .D1(d4[59]), .CIN(n12100), 
          .COUT(n12101), .S0(d5_71__N_706[58]), .S1(d5_71__N_706[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1065_25.INIT0 = 16'h74b8;
    defparam add_1065_25.INIT1 = 16'h74b8;
    defparam add_1065_25.INJECT1_0 = "NO";
    defparam add_1065_25.INJECT1_1 = "NO";
    CCU2D add_1065_23 (.A0(d5[56]), .B0(n4884), .C0(n4885[20]), .D0(d4[56]), 
          .A1(d5[57]), .B1(n4884), .C1(n4885[21]), .D1(d4[57]), .CIN(n12099), 
          .COUT(n12100), .S0(d5_71__N_706[56]), .S1(d5_71__N_706[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1065_23.INIT0 = 16'h74b8;
    defparam add_1065_23.INIT1 = 16'h74b8;
    defparam add_1065_23.INJECT1_0 = "NO";
    defparam add_1065_23.INJECT1_1 = "NO";
    CCU2D add_1065_21 (.A0(d5[54]), .B0(n4884), .C0(n4885[18]), .D0(d4[54]), 
          .A1(d5[55]), .B1(n4884), .C1(n4885[19]), .D1(d4[55]), .CIN(n12098), 
          .COUT(n12099), .S0(d5_71__N_706[54]), .S1(d5_71__N_706[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1065_21.INIT0 = 16'h74b8;
    defparam add_1065_21.INIT1 = 16'h74b8;
    defparam add_1065_21.INJECT1_0 = "NO";
    defparam add_1065_21.INJECT1_1 = "NO";
    PFUMX i5794 (.BLUT(n13394), .ALUT(n13395), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[0]));
    CCU2D add_1065_19 (.A0(d5[52]), .B0(n4884), .C0(n4885[16]), .D0(d4[52]), 
          .A1(d5[53]), .B1(n4884), .C1(n4885[17]), .D1(d4[53]), .CIN(n12097), 
          .COUT(n12098), .S0(d5_71__N_706[52]), .S1(d5_71__N_706[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1065_19.INIT0 = 16'h74b8;
    defparam add_1065_19.INIT1 = 16'h74b8;
    defparam add_1065_19.INJECT1_0 = "NO";
    defparam add_1065_19.INJECT1_1 = "NO";
    CCU2D add_1065_17 (.A0(d5[50]), .B0(n4884), .C0(n4885[14]), .D0(d4[50]), 
          .A1(d5[51]), .B1(n4884), .C1(n4885[15]), .D1(d4[51]), .CIN(n12096), 
          .COUT(n12097), .S0(d5_71__N_706[50]), .S1(d5_71__N_706[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1065_17.INIT0 = 16'h74b8;
    defparam add_1065_17.INIT1 = 16'h74b8;
    defparam add_1065_17.INJECT1_0 = "NO";
    defparam add_1065_17.INJECT1_1 = "NO";
    CCU2D add_1065_15 (.A0(d5[48]), .B0(n4884), .C0(n4885[12]), .D0(d4[48]), 
          .A1(d5[49]), .B1(n4884), .C1(n4885[13]), .D1(d4[49]), .CIN(n12095), 
          .COUT(n12096), .S0(d5_71__N_706[48]), .S1(d5_71__N_706[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1065_15.INIT0 = 16'h74b8;
    defparam add_1065_15.INIT1 = 16'h74b8;
    defparam add_1065_15.INJECT1_0 = "NO";
    defparam add_1065_15.INJECT1_1 = "NO";
    CCU2D add_1065_13 (.A0(d5[46]), .B0(n4884), .C0(n4885[10]), .D0(d4[46]), 
          .A1(d5[47]), .B1(n4884), .C1(n4885[11]), .D1(d4[47]), .CIN(n12094), 
          .COUT(n12095), .S0(d5_71__N_706[46]), .S1(d5_71__N_706[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1065_13.INIT0 = 16'h74b8;
    defparam add_1065_13.INIT1 = 16'h74b8;
    defparam add_1065_13.INJECT1_0 = "NO";
    defparam add_1065_13.INJECT1_1 = "NO";
    CCU2D add_1065_11 (.A0(d5[44]), .B0(n4884), .C0(n4885[8]), .D0(d4[44]), 
          .A1(d5[45]), .B1(n4884), .C1(n4885[9]), .D1(d4[45]), .CIN(n12093), 
          .COUT(n12094), .S0(d5_71__N_706[44]), .S1(d5_71__N_706[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1065_11.INIT0 = 16'h74b8;
    defparam add_1065_11.INIT1 = 16'h74b8;
    defparam add_1065_11.INJECT1_0 = "NO";
    defparam add_1065_11.INJECT1_1 = "NO";
    CCU2D add_1065_9 (.A0(d5[42]), .B0(n4884), .C0(n4885[6]), .D0(d4[42]), 
          .A1(d5[43]), .B1(n4884), .C1(n4885[7]), .D1(d4[43]), .CIN(n12092), 
          .COUT(n12093), .S0(d5_71__N_706[42]), .S1(d5_71__N_706[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1065_9.INIT0 = 16'h74b8;
    defparam add_1065_9.INIT1 = 16'h74b8;
    defparam add_1065_9.INJECT1_0 = "NO";
    defparam add_1065_9.INJECT1_1 = "NO";
    CCU2D add_1065_7 (.A0(d5[40]), .B0(n4884), .C0(n4885[4]), .D0(d4[40]), 
          .A1(d5[41]), .B1(n4884), .C1(n4885[5]), .D1(d4[41]), .CIN(n12091), 
          .COUT(n12092), .S0(d5_71__N_706[40]), .S1(d5_71__N_706[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1065_7.INIT0 = 16'h74b8;
    defparam add_1065_7.INIT1 = 16'h74b8;
    defparam add_1065_7.INJECT1_0 = "NO";
    defparam add_1065_7.INJECT1_1 = "NO";
    PFUMX i5792 (.BLUT(n13391), .ALUT(n13392), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[1]));
    CCU2D add_1065_5 (.A0(d5[38]), .B0(n4884), .C0(n4885[2]), .D0(d4[38]), 
          .A1(d5[39]), .B1(n4884), .C1(n4885[3]), .D1(d4[39]), .CIN(n12090), 
          .COUT(n12091), .S0(d5_71__N_706[38]), .S1(d5_71__N_706[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1065_5.INIT0 = 16'h74b8;
    defparam add_1065_5.INIT1 = 16'h74b8;
    defparam add_1065_5.INJECT1_0 = "NO";
    defparam add_1065_5.INJECT1_1 = "NO";
    CCU2D add_1065_3 (.A0(d5[36]), .B0(n4884), .C0(n4885[0]), .D0(d4[36]), 
          .A1(d5[37]), .B1(n4884), .C1(n4885[1]), .D1(d4[37]), .CIN(n12089), 
          .COUT(n12090), .S0(d5_71__N_706[36]), .S1(d5_71__N_706[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1065_3.INIT0 = 16'h74b8;
    defparam add_1065_3.INIT1 = 16'h74b8;
    defparam add_1065_3.INJECT1_0 = "NO";
    defparam add_1065_3.INJECT1_1 = "NO";
    CCU2D add_1065_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n4884), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n12089));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1065_1.INIT0 = 16'hF000;
    defparam add_1065_1.INIT1 = 16'h0555;
    defparam add_1065_1.INJECT1_0 = "NO";
    defparam add_1065_1.INJECT1_1 = "NO";
    CCU2D add_1045_37 (.A0(d1[70]), .B0(n4276), .C0(n4277[34]), .D0(MixerOutSin[11]), 
          .A1(d1[71]), .B1(n4276), .C1(n4277[35]), .D1(MixerOutSin[11]), 
          .CIN(n12270), .S0(d1_71__N_418[70]), .S1(d1_71__N_418[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1045_37.INIT0 = 16'h74b8;
    defparam add_1045_37.INIT1 = 16'h74b8;
    defparam add_1045_37.INJECT1_0 = "NO";
    defparam add_1045_37.INJECT1_1 = "NO";
    CCU2D add_1045_35 (.A0(d1[68]), .B0(n4276), .C0(n4277[32]), .D0(MixerOutSin[11]), 
          .A1(d1[69]), .B1(n4276), .C1(n4277[33]), .D1(MixerOutSin[11]), 
          .CIN(n12269), .COUT(n12270), .S0(d1_71__N_418[68]), .S1(d1_71__N_418[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1045_35.INIT0 = 16'h74b8;
    defparam add_1045_35.INIT1 = 16'h74b8;
    defparam add_1045_35.INJECT1_0 = "NO";
    defparam add_1045_35.INJECT1_1 = "NO";
    CCU2D add_1045_33 (.A0(d1[66]), .B0(n4276), .C0(n4277[30]), .D0(MixerOutSin[11]), 
          .A1(d1[67]), .B1(n4276), .C1(n4277[31]), .D1(MixerOutSin[11]), 
          .CIN(n12268), .COUT(n12269), .S0(d1_71__N_418[66]), .S1(d1_71__N_418[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1045_33.INIT0 = 16'h74b8;
    defparam add_1045_33.INIT1 = 16'h74b8;
    defparam add_1045_33.INJECT1_0 = "NO";
    defparam add_1045_33.INJECT1_1 = "NO";
    CCU2D add_1045_31 (.A0(d1[64]), .B0(n4276), .C0(n4277[28]), .D0(MixerOutSin[11]), 
          .A1(d1[65]), .B1(n4276), .C1(n4277[29]), .D1(MixerOutSin[11]), 
          .CIN(n12267), .COUT(n12268), .S0(d1_71__N_418[64]), .S1(d1_71__N_418[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1045_31.INIT0 = 16'h74b8;
    defparam add_1045_31.INIT1 = 16'h74b8;
    defparam add_1045_31.INJECT1_0 = "NO";
    defparam add_1045_31.INJECT1_1 = "NO";
    CCU2D add_1045_29 (.A0(d1[62]), .B0(n4276), .C0(n4277[26]), .D0(MixerOutSin[11]), 
          .A1(d1[63]), .B1(n4276), .C1(n4277[27]), .D1(MixerOutSin[11]), 
          .CIN(n12266), .COUT(n12267), .S0(d1_71__N_418[62]), .S1(d1_71__N_418[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1045_29.INIT0 = 16'h74b8;
    defparam add_1045_29.INIT1 = 16'h74b8;
    defparam add_1045_29.INJECT1_0 = "NO";
    defparam add_1045_29.INJECT1_1 = "NO";
    FD1S3AX v_comb_66_rep_93 (.D(osc_clk_enable_1458), .CK(osc_clk), .Q(osc_clk_enable_647)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=168, LSE_RLINE=174 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_93.GSR = "ENABLED";
    CCU2D add_1045_27 (.A0(d1[60]), .B0(n4276), .C0(n4277[24]), .D0(MixerOutSin[11]), 
          .A1(d1[61]), .B1(n4276), .C1(n4277[25]), .D1(MixerOutSin[11]), 
          .CIN(n12265), .COUT(n12266), .S0(d1_71__N_418[60]), .S1(d1_71__N_418[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1045_27.INIT0 = 16'h74b8;
    defparam add_1045_27.INIT1 = 16'h74b8;
    defparam add_1045_27.INJECT1_0 = "NO";
    defparam add_1045_27.INJECT1_1 = "NO";
    CCU2D add_1045_25 (.A0(d1[58]), .B0(n4276), .C0(n4277[22]), .D0(MixerOutSin[11]), 
          .A1(d1[59]), .B1(n4276), .C1(n4277[23]), .D1(MixerOutSin[11]), 
          .CIN(n12264), .COUT(n12265), .S0(d1_71__N_418[58]), .S1(d1_71__N_418[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1045_25.INIT0 = 16'h74b8;
    defparam add_1045_25.INIT1 = 16'h74b8;
    defparam add_1045_25.INJECT1_0 = "NO";
    defparam add_1045_25.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \CIC(width=72,decimation_ratio=4096)_U1 
//

module \CIC(width=72,decimation_ratio=4096)_U1  (GND_net, MixerOutCos, osc_clk, 
            CIC1_outCos, \d10[59] , \d10[60] , \d10[61] , \d10[62] , 
            \d10[63] , \d10[64] , \d10[65] , \d10[66] , \d10[67] , 
            \d10[68] , \d10[69] , \d10[70] , \d10[71] , \d_out_11__N_1819[2] , 
            \d_out_11__N_1819[3] , \d_out_11__N_1819[4] , \d_out_11__N_1819[5] , 
            \d_out_11__N_1819[6] , \d_out_11__N_1819[7] , \d_out_11__N_1819[8] , 
            \d_out_11__N_1819[9] , \d_out_11__N_1819[10] , \d_out_11__N_1819[11] , 
            \CICGain[0] , n61, n70, \CICGain[1] , n62, n63, n64, 
            n65, n66, n67, n68) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input [11:0]MixerOutCos;
    input osc_clk;
    output [11:0]CIC1_outCos;
    output \d10[59] ;
    output \d10[60] ;
    output \d10[61] ;
    output \d10[62] ;
    output \d10[63] ;
    output \d10[64] ;
    output \d10[65] ;
    output \d10[66] ;
    output \d10[67] ;
    output \d10[68] ;
    output \d10[69] ;
    output \d10[70] ;
    output \d10[71] ;
    input \d_out_11__N_1819[2] ;
    input \d_out_11__N_1819[3] ;
    input \d_out_11__N_1819[4] ;
    input \d_out_11__N_1819[5] ;
    input \d_out_11__N_1819[6] ;
    input \d_out_11__N_1819[7] ;
    input \d_out_11__N_1819[8] ;
    input \d_out_11__N_1819[9] ;
    input \d_out_11__N_1819[10] ;
    input \d_out_11__N_1819[11] ;
    input \CICGain[0] ;
    output n61;
    output n70;
    input \CICGain[1] ;
    output n62;
    output n63;
    output n64;
    output n65;
    output n66;
    output n67;
    output n68;
    
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(71[8:15])
    
    wire n12035;
    wire [71:0]d1;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(35[26:28])
    wire [71:0]d2;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(36[26:28])
    wire [35:0]n5189;
    
    wire n12036, n12034, n12033, n11976;
    wire [71:0]d3;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(37[26:28])
    
    wire n5340;
    wire [35:0]n5341;
    wire [71:0]d3_71__N_562;
    
    wire n11977, n13121, n13, n13123, n13103, osc_clk_enable_744, 
        n11898;
    wire [71:0]d5;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(39[26:28])
    
    wire n5644;
    wire [35:0]n5645;
    wire [71:0]d4;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(38[26:28])
    wire [71:0]d5_71__N_706;
    
    wire n11899, n12054, n5036;
    wire [35:0]n5037;
    wire [71:0]d1_71__N_418;
    
    wire n12055, n11975, n12053, n12052, n12050, n12051;
    wire [71:0]d_tmp;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(30[26:31])
    wire [71:0]d_d_tmp;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(30[33:40])
    
    wire osc_clk_enable_784;
    wire [71:0]d2_71__N_490;
    wire [71:0]d4_71__N_634;
    wire [71:0]d6;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(43[26:28])
    wire [71:0]d6_71__N_1459;
    wire [71:0]d_d6;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(43[30:34])
    
    wire v_comb;
    wire [71:0]d7;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(44[26:28])
    wire [71:0]d7_71__N_1531;
    wire [71:0]d_d7;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(44[30:34])
    wire [71:0]d8;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(45[26:28])
    wire [71:0]d8_71__N_1603;
    wire [71:0]d_d8;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(45[30:34])
    wire [71:0]d9;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(46[26:28])
    wire [71:0]d9_71__N_1675;
    wire [71:0]d_d9;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(46[30:34])
    wire [71:0]d_out_11__N_1819;
    
    wire n11909, n11910, n12042, n12043, n11901, n12041, n12040, 
        n12039, n12038, n11974, n12037, n11973, n11897, n12019, 
        n5188, n12020, n12028, n12029, n11896, n11895, n11908, 
        n11972, n12017, n12018, n12016, n12013, n12014, n12010, 
        n12011, n12012, n12015, n12009, n11971, n11970, n11907, 
        n11623;
    wire [35:0]n6101;
    wire [15:0]count;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(50[14:19])
    wire [15:0]count_15__N_1442;
    
    wire n11969, n11968, n11967, n11906, n11966, n11905, n12008, 
        n12002, n11894, n11992, n11993, n11991, n11990, n11988, 
        n11989, n11987, n11904;
    wire [15:0]n375;
    
    wire n31, n11986, n11983, n11978, n11982, n11981, n11980, 
        n11979, n11893, n12021, n12022, n12032, n21, n19, n15, 
        n16, n11892, n11891, n11890, n11889, n11888, n11887, n11886, 
        n11885, n11884, n12031, n12030, n12027, n12024, n12023, 
        n11622, n11621, n11620, n11619, n11618, n11617, n11616, 
        n11615, n11614, n11996, n11997, n11613, n11612, n11611, 
        n11961;
    wire [35:0]n5493;
    
    wire n11995, n11960, n12001, n11994, n12000, n12007, n11999, 
        n11959, n11998, n12049, n12048, n11900, count_15__N_1458, 
        n12790, n11958, n11957, n11956, n11955, n11954, n11953, 
        n11952, n11951, n11610, n11950, n11949, n11948, n11947, 
        n11946, n11945, n11942, n5492, n11941, n11940, n7, n11939, 
        n11938, n11937, n11936, n13507, n11935, n11934, n11933, 
        n11932, n11931, n11930, n11929, n11928, n11927, n11926, 
        n11925, n11920, n11919, n11918, n11917, n11916, n11915, 
        n11914, n11913, n11912, osc_clk_enable_834, osc_clk_enable_884, 
        osc_clk_enable_934, osc_clk_enable_984, osc_clk_enable_1034, osc_clk_enable_1084, 
        osc_clk_enable_1134, osc_clk_enable_1184, osc_clk_enable_1234, 
        osc_clk_enable_1284, osc_clk_enable_1334, osc_clk_enable_1384;
    wire [71:0]d10;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(47[26:29])
    wire [71:0]d10_71__N_1747;
    
    wire n11609, n11608, n11607, n11606, n11604, n6100, n11603, 
        n11602, n11601, n11600, n11599, n11598, n11597, n11596, 
        n11595, n11594, n11593, n11592, n11591, n11590, n11589, 
        n11588, n11587, n11583;
    wire [35:0]n6253;
    
    wire n11582, n11581, n11580, n11579, n11578, n11577, n11576, 
        n11575, n11574, n11573, n11572, n11571, n11570, n11569, 
        n11568, n11567, n11566, n11564, n6252, n11563, n11562, 
        n11561, n11560, n11559, n11558, n11557, n11556, n11555, 
        n11554, n11553, n11552, n11551, n11550, n11549, n11548, 
        n11547, n11543;
    wire [35:0]n6405;
    
    wire n11542, n11541, n11540, n11539, n11538, n11537, n11536, 
        n11535, n11534, n11533, n11532, n11531, n11530, n11529, 
        n11528, n11527, n11526, n11524, n6404, n11523, n11522, 
        n11521, n11520, n11519, n11518, n11517, n11516, n11515, 
        n11514, n11513, n11512, n11511, n11510, n11509, n11508, 
        n11507, n11503;
    wire [35:0]n6557;
    
    wire n11502, n11501, n11500, n11499, n11498, n11497, n11496, 
        n11495, n11494, n11493, n11492, n11491, n11490, n11489, 
        n11488, n11487, n11486, n11484, n6556, n11483, n11482, 
        n11481, n11480, n11479, n11478, n11477, n11476, n11475, 
        n11474, n11473, n11472, n11471, n11470, n11469, n11468, 
        n11467, n11463;
    wire [35:0]n6709;
    
    wire n11462, n11461, n11460, n11459, n11458, n11457, n11456, 
        n11455, n11454, n11453, n11452, n11451, n11450, n11449, 
        n11448, n11447, n11446, n11445;
    wire [35:0]n6747;
    
    wire n11444, n11443, n11442, n11441, n11440, n11439, n11438, 
        n11437, n11436, n11435, n11434, n11433, n11432, n11431, 
        n11430, n11429, n11428, n8387, n11231, n11230, n11229, 
        n11228, n11227, n11226, n11225, n11224, n11205, n11204, 
        n11203, n11202, n11201, n11200, n11199, n11198, n11197, 
        n11196, n11195, n11194, n11193, n11192, n11191, n11190, 
        n11189, n11188, n11186, n11185, n11184, n11183, n11182, 
        n11181, n11180, n11179, n11178, n11177, n11176, n11175, 
        n11174, n11173, n11172, n11171, n11170, n11169, n11167, 
        n11166, n11165, n11164, n11163, n11162, n11161, n11160, 
        n11159, n11158, n11157, n11156, n11155, n11154, n11153, 
        n11152, n11151, n11150, n11148, n11147, n11146, n11145, 
        n11144, n11143, n11142, n11141, n11140, n11139, n11138, 
        n11137, n11136, n11135, n11134, n11133, n11132, n11131, 
        n11091, n11090, n11089, n11088, n11087, n11086, n11085, 
        n11084, n11083, n11082, n11081, n11080, n11079, n11078, 
        n11077, n11076, n11075, n11074, n11745, n6708, n11744, 
        n11743, n11742, n11741, n11740, n11739, n11738, n11737, 
        n11736, n11735, n11734, n11733, n11732, n11731, n11730, 
        n11729, n11728, n11727, n11726, n11725, n11724, n11723, 
        n11722, n11721, n11720, n11719, n11718, n11717, n11716, 
        n11715, n11714, n11713, n11712, n11711, n11710, n11709, 
        n11708, n11707, n11706, n11705, n11704, n11703, n11702, 
        n11701, n11700, n11699, n11698, n11697, n11696, n11695, 
        n11694, n11693, n11692, n11691, n11690, n11689, n11688, 
        n11687, n11686, n11685, n11684, n11683, n11682, n11681, 
        n11680, n11679, n11678, n11677, n11676, n11675, n11674, 
        n11673, n11672, n11671, n11670, n11669, n11668, n11667, 
        n11666, n11665, n11664, n11663, n11662, n11661, n11660, 
        n11659, n11658, n11657, n11656, n13404, n13403, n13407, 
        n13406, n12056, n11911, n12059, n12060, n12071, n12072, 
        n12070, n12069, n12068, n12065, n12064, n12063, n12062, 
        n12058, n12057, n12061, n12084, n12083, n12082, n12081, 
        n12080, n12079, n12078, n12077, n12076, n12075, n12074, 
        n12073;
    
    CCU2D add_1074_20 (.A0(d1[54]), .B0(d2[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[55]), .B1(d2[55]), .C1(GND_net), .D1(GND_net), .CIN(n12035), 
          .COUT(n12036), .S0(n5189[18]), .S1(n5189[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1074_20.INIT0 = 16'h5666;
    defparam add_1074_20.INIT1 = 16'h5666;
    defparam add_1074_20.INJECT1_0 = "NO";
    defparam add_1074_20.INJECT1_1 = "NO";
    CCU2D add_1074_18 (.A0(d1[52]), .B0(d2[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[53]), .B1(d2[53]), .C1(GND_net), .D1(GND_net), .CIN(n12034), 
          .COUT(n12035), .S0(n5189[16]), .S1(n5189[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1074_18.INIT0 = 16'h5666;
    defparam add_1074_18.INIT1 = 16'h5666;
    defparam add_1074_18.INJECT1_0 = "NO";
    defparam add_1074_18.INJECT1_1 = "NO";
    CCU2D add_1074_16 (.A0(d1[50]), .B0(d2[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[51]), .B1(d2[51]), .C1(GND_net), .D1(GND_net), .CIN(n12033), 
          .COUT(n12034), .S0(n5189[14]), .S1(n5189[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1074_16.INIT0 = 16'h5666;
    defparam add_1074_16.INIT1 = 16'h5666;
    defparam add_1074_16.INJECT1_0 = "NO";
    defparam add_1074_16.INJECT1_1 = "NO";
    CCU2D add_1080_23 (.A0(d3[56]), .B0(n5340), .C0(n5341[20]), .D0(d2[56]), 
          .A1(d3[57]), .B1(n5340), .C1(n5341[21]), .D1(d2[57]), .CIN(n11976), 
          .COUT(n11977), .S0(d3_71__N_562[56]), .S1(d3_71__N_562[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1080_23.INIT0 = 16'h74b8;
    defparam add_1080_23.INIT1 = 16'h74b8;
    defparam add_1080_23.INJECT1_0 = "NO";
    defparam add_1080_23.INJECT1_1 = "NO";
    LUT4 i5686_4_lut_rep_98 (.A(n13121), .B(n13), .C(n13123), .D(n13103), 
         .Z(osc_clk_enable_744)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i5686_4_lut_rep_98.init = 16'h2000;
    CCU2D add_1090_31 (.A0(d5[64]), .B0(n5644), .C0(n5645[28]), .D0(d4[64]), 
          .A1(d5[65]), .B1(n5644), .C1(n5645[29]), .D1(d4[65]), .CIN(n11898), 
          .COUT(n11899), .S0(d5_71__N_706[64]), .S1(d5_71__N_706[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1090_31.INIT0 = 16'h74b8;
    defparam add_1090_31.INIT1 = 16'h74b8;
    defparam add_1090_31.INJECT1_0 = "NO";
    defparam add_1090_31.INJECT1_1 = "NO";
    CCU2D add_1070_15 (.A0(d1[48]), .B0(n5036), .C0(n5037[12]), .D0(MixerOutCos[11]), 
          .A1(d1[49]), .B1(n5036), .C1(n5037[13]), .D1(MixerOutCos[11]), 
          .CIN(n12054), .COUT(n12055), .S0(d1_71__N_418[48]), .S1(d1_71__N_418[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1070_15.INIT0 = 16'h74b8;
    defparam add_1070_15.INIT1 = 16'h74b8;
    defparam add_1070_15.INJECT1_0 = "NO";
    defparam add_1070_15.INJECT1_1 = "NO";
    CCU2D add_1080_21 (.A0(d3[54]), .B0(n5340), .C0(n5341[18]), .D0(d2[54]), 
          .A1(d3[55]), .B1(n5340), .C1(n5341[19]), .D1(d2[55]), .CIN(n11975), 
          .COUT(n11976), .S0(d3_71__N_562[54]), .S1(d3_71__N_562[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1080_21.INIT0 = 16'h74b8;
    defparam add_1080_21.INIT1 = 16'h74b8;
    defparam add_1080_21.INJECT1_0 = "NO";
    defparam add_1080_21.INJECT1_1 = "NO";
    CCU2D add_1070_13 (.A0(d1[46]), .B0(n5036), .C0(n5037[10]), .D0(MixerOutCos[11]), 
          .A1(d1[47]), .B1(n5036), .C1(n5037[11]), .D1(MixerOutCos[11]), 
          .CIN(n12053), .COUT(n12054), .S0(d1_71__N_418[46]), .S1(d1_71__N_418[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1070_13.INIT0 = 16'h74b8;
    defparam add_1070_13.INIT1 = 16'h74b8;
    defparam add_1070_13.INJECT1_0 = "NO";
    defparam add_1070_13.INJECT1_1 = "NO";
    CCU2D add_1070_11 (.A0(d1[44]), .B0(n5036), .C0(n5037[8]), .D0(MixerOutCos[11]), 
          .A1(d1[45]), .B1(n5036), .C1(n5037[9]), .D1(MixerOutCos[11]), 
          .CIN(n12052), .COUT(n12053), .S0(d1_71__N_418[44]), .S1(d1_71__N_418[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1070_11.INIT0 = 16'h74b8;
    defparam add_1070_11.INIT1 = 16'h74b8;
    defparam add_1070_11.INJECT1_0 = "NO";
    defparam add_1070_11.INJECT1_1 = "NO";
    CCU2D add_1070_7 (.A0(d1[40]), .B0(n5036), .C0(n5037[4]), .D0(MixerOutCos[11]), 
          .A1(d1[41]), .B1(n5036), .C1(n5037[5]), .D1(MixerOutCos[11]), 
          .CIN(n12050), .COUT(n12051), .S0(d1_71__N_418[40]), .S1(d1_71__N_418[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1070_7.INIT0 = 16'h74b8;
    defparam add_1070_7.INIT1 = 16'h74b8;
    defparam add_1070_7.INJECT1_0 = "NO";
    defparam add_1070_7.INJECT1_1 = "NO";
    FD1P3AX d_tmp_i0_i0 (.D(d5[0]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i0 (.D(d_tmp[0]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i0.GSR = "ENABLED";
    FD1S3AX d2_i0 (.D(d2_71__N_490[0]), .CK(osc_clk), .Q(d2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i0.GSR = "ENABLED";
    FD1S3AX d3_i0 (.D(d3_71__N_562[0]), .CK(osc_clk), .Q(d3[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i0.GSR = "ENABLED";
    FD1S3AX d4_i0 (.D(d4_71__N_634[0]), .CK(osc_clk), .Q(d4[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i0.GSR = "ENABLED";
    FD1S3AX d5_i0 (.D(d5_71__N_706[0]), .CK(osc_clk), .Q(d5[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i0.GSR = "ENABLED";
    FD1P3AX d6_i0_i0 (.D(d6_71__N_1459[0]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i0 (.D(d6[0]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i0.GSR = "ENABLED";
    FD1S3AX v_comb_66 (.D(osc_clk_enable_744), .CK(osc_clk), .Q(v_comb)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66.GSR = "ENABLED";
    FD1P3AX d7_i0_i0 (.D(d7_71__N_1531[0]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i0 (.D(d7[0]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d8_i0_i0 (.D(d8_71__N_1603[0]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i0 (.D(d8[0]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d9_i0_i0 (.D(d9_71__N_1675[0]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i0 (.D(d9[0]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_out_i0_i0 (.D(d_out_11__N_1819[0]), .SP(osc_clk_enable_784), 
            .CK(osc_clk), .Q(CIC1_outCos[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i0.GSR = "ENABLED";
    FD1S3AX d1_i0 (.D(d1_71__N_418[0]), .CK(osc_clk), .Q(d1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i0.GSR = "ENABLED";
    CCU2D add_1070_9 (.A0(d1[42]), .B0(n5036), .C0(n5037[6]), .D0(MixerOutCos[11]), 
          .A1(d1[43]), .B1(n5036), .C1(n5037[7]), .D1(MixerOutCos[11]), 
          .CIN(n12051), .COUT(n12052), .S0(d1_71__N_418[42]), .S1(d1_71__N_418[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1070_9.INIT0 = 16'h74b8;
    defparam add_1070_9.INIT1 = 16'h74b8;
    defparam add_1070_9.INJECT1_0 = "NO";
    defparam add_1070_9.INJECT1_1 = "NO";
    CCU2D add_1089_14 (.A0(d4[48]), .B0(d5[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[49]), .B1(d5[49]), .C1(GND_net), .D1(GND_net), .CIN(n11909), 
          .COUT(n11910), .S0(n5645[12]), .S1(n5645[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1089_14.INIT0 = 16'h5666;
    defparam add_1089_14.INIT1 = 16'h5666;
    defparam add_1089_14.INJECT1_0 = "NO";
    defparam add_1089_14.INJECT1_1 = "NO";
    CCU2D add_1074_34 (.A0(d1[68]), .B0(d2[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[69]), .B1(d2[69]), .C1(GND_net), .D1(GND_net), .CIN(n12042), 
          .COUT(n12043), .S0(n5189[32]), .S1(n5189[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1074_34.INIT0 = 16'h5666;
    defparam add_1074_34.INIT1 = 16'h5666;
    defparam add_1074_34.INJECT1_0 = "NO";
    defparam add_1074_34.INJECT1_1 = "NO";
    CCU2D add_1090_37 (.A0(d5[70]), .B0(n5644), .C0(n5645[34]), .D0(d4[70]), 
          .A1(d5[71]), .B1(n5644), .C1(n5645[35]), .D1(d4[71]), .CIN(n11901), 
          .S0(d5_71__N_706[70]), .S1(d5_71__N_706[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1090_37.INIT0 = 16'h74b8;
    defparam add_1090_37.INIT1 = 16'h74b8;
    defparam add_1090_37.INJECT1_0 = "NO";
    defparam add_1090_37.INJECT1_1 = "NO";
    CCU2D add_1074_32 (.A0(d1[66]), .B0(d2[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[67]), .B1(d2[67]), .C1(GND_net), .D1(GND_net), .CIN(n12041), 
          .COUT(n12042), .S0(n5189[30]), .S1(n5189[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1074_32.INIT0 = 16'h5666;
    defparam add_1074_32.INIT1 = 16'h5666;
    defparam add_1074_32.INJECT1_0 = "NO";
    defparam add_1074_32.INJECT1_1 = "NO";
    CCU2D add_1074_30 (.A0(d1[64]), .B0(d2[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[65]), .B1(d2[65]), .C1(GND_net), .D1(GND_net), .CIN(n12040), 
          .COUT(n12041), .S0(n5189[28]), .S1(n5189[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1074_30.INIT0 = 16'h5666;
    defparam add_1074_30.INIT1 = 16'h5666;
    defparam add_1074_30.INJECT1_0 = "NO";
    defparam add_1074_30.INJECT1_1 = "NO";
    CCU2D add_1074_28 (.A0(d1[62]), .B0(d2[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[63]), .B1(d2[63]), .C1(GND_net), .D1(GND_net), .CIN(n12039), 
          .COUT(n12040), .S0(n5189[26]), .S1(n5189[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1074_28.INIT0 = 16'h5666;
    defparam add_1074_28.INIT1 = 16'h5666;
    defparam add_1074_28.INJECT1_0 = "NO";
    defparam add_1074_28.INJECT1_1 = "NO";
    CCU2D add_1074_26 (.A0(d1[60]), .B0(d2[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[61]), .B1(d2[61]), .C1(GND_net), .D1(GND_net), .CIN(n12038), 
          .COUT(n12039), .S0(n5189[24]), .S1(n5189[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1074_26.INIT0 = 16'h5666;
    defparam add_1074_26.INIT1 = 16'h5666;
    defparam add_1074_26.INJECT1_0 = "NO";
    defparam add_1074_26.INJECT1_1 = "NO";
    CCU2D add_1080_19 (.A0(d3[52]), .B0(n5340), .C0(n5341[16]), .D0(d2[52]), 
          .A1(d3[53]), .B1(n5340), .C1(n5341[17]), .D1(d2[53]), .CIN(n11974), 
          .COUT(n11975), .S0(d3_71__N_562[52]), .S1(d3_71__N_562[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1080_19.INIT0 = 16'h74b8;
    defparam add_1080_19.INIT1 = 16'h74b8;
    defparam add_1080_19.INJECT1_0 = "NO";
    defparam add_1080_19.INJECT1_1 = "NO";
    CCU2D add_1074_24 (.A0(d1[58]), .B0(d2[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[59]), .B1(d2[59]), .C1(GND_net), .D1(GND_net), .CIN(n12037), 
          .COUT(n12038), .S0(n5189[22]), .S1(n5189[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1074_24.INIT0 = 16'h5666;
    defparam add_1074_24.INIT1 = 16'h5666;
    defparam add_1074_24.INJECT1_0 = "NO";
    defparam add_1074_24.INJECT1_1 = "NO";
    CCU2D add_1080_17 (.A0(d3[50]), .B0(n5340), .C0(n5341[14]), .D0(d2[50]), 
          .A1(d3[51]), .B1(n5340), .C1(n5341[15]), .D1(d2[51]), .CIN(n11973), 
          .COUT(n11974), .S0(d3_71__N_562[50]), .S1(d3_71__N_562[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1080_17.INIT0 = 16'h74b8;
    defparam add_1080_17.INIT1 = 16'h74b8;
    defparam add_1080_17.INJECT1_0 = "NO";
    defparam add_1080_17.INJECT1_1 = "NO";
    CCU2D add_1074_22 (.A0(d1[56]), .B0(d2[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[57]), .B1(d2[57]), .C1(GND_net), .D1(GND_net), .CIN(n12036), 
          .COUT(n12037), .S0(n5189[20]), .S1(n5189[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1074_22.INIT0 = 16'h5666;
    defparam add_1074_22.INIT1 = 16'h5666;
    defparam add_1074_22.INJECT1_0 = "NO";
    defparam add_1074_22.INJECT1_1 = "NO";
    CCU2D add_1090_29 (.A0(d5[62]), .B0(n5644), .C0(n5645[26]), .D0(d4[62]), 
          .A1(d5[63]), .B1(n5644), .C1(n5645[27]), .D1(d4[63]), .CIN(n11897), 
          .COUT(n11898), .S0(d5_71__N_706[62]), .S1(d5_71__N_706[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1090_29.INIT0 = 16'h74b8;
    defparam add_1090_29.INIT1 = 16'h74b8;
    defparam add_1090_29.INJECT1_0 = "NO";
    defparam add_1090_29.INJECT1_1 = "NO";
    CCU2D add_1075_27 (.A0(d2[60]), .B0(n5188), .C0(n5189[24]), .D0(d1[60]), 
          .A1(d2[61]), .B1(n5188), .C1(n5189[25]), .D1(d1[61]), .CIN(n12019), 
          .COUT(n12020), .S0(d2_71__N_490[60]), .S1(d2_71__N_490[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1075_27.INIT0 = 16'h74b8;
    defparam add_1075_27.INIT1 = 16'h74b8;
    defparam add_1075_27.INJECT1_0 = "NO";
    defparam add_1075_27.INJECT1_1 = "NO";
    CCU2D add_1074_6 (.A0(d1[40]), .B0(d2[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[41]), .B1(d2[41]), .C1(GND_net), .D1(GND_net), .CIN(n12028), 
          .COUT(n12029), .S0(n5189[4]), .S1(n5189[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1074_6.INIT0 = 16'h5666;
    defparam add_1074_6.INIT1 = 16'h5666;
    defparam add_1074_6.INJECT1_0 = "NO";
    defparam add_1074_6.INJECT1_1 = "NO";
    CCU2D add_1090_27 (.A0(d5[60]), .B0(n5644), .C0(n5645[24]), .D0(d4[60]), 
          .A1(d5[61]), .B1(n5644), .C1(n5645[25]), .D1(d4[61]), .CIN(n11896), 
          .COUT(n11897), .S0(d5_71__N_706[60]), .S1(d5_71__N_706[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1090_27.INIT0 = 16'h74b8;
    defparam add_1090_27.INIT1 = 16'h74b8;
    defparam add_1090_27.INJECT1_0 = "NO";
    defparam add_1090_27.INJECT1_1 = "NO";
    CCU2D add_1090_25 (.A0(d5[58]), .B0(n5644), .C0(n5645[22]), .D0(d4[58]), 
          .A1(d5[59]), .B1(n5644), .C1(n5645[23]), .D1(d4[59]), .CIN(n11895), 
          .COUT(n11896), .S0(d5_71__N_706[58]), .S1(d5_71__N_706[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1090_25.INIT0 = 16'h74b8;
    defparam add_1090_25.INIT1 = 16'h74b8;
    defparam add_1090_25.INJECT1_0 = "NO";
    defparam add_1090_25.INJECT1_1 = "NO";
    CCU2D add_1089_12 (.A0(d4[46]), .B0(d5[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[47]), .B1(d5[47]), .C1(GND_net), .D1(GND_net), .CIN(n11908), 
          .COUT(n11909), .S0(n5645[10]), .S1(n5645[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1089_12.INIT0 = 16'h5666;
    defparam add_1089_12.INIT1 = 16'h5666;
    defparam add_1089_12.INJECT1_0 = "NO";
    defparam add_1089_12.INJECT1_1 = "NO";
    CCU2D add_1080_15 (.A0(d3[48]), .B0(n5340), .C0(n5341[12]), .D0(d2[48]), 
          .A1(d3[49]), .B1(n5340), .C1(n5341[13]), .D1(d2[49]), .CIN(n11972), 
          .COUT(n11973), .S0(d3_71__N_562[48]), .S1(d3_71__N_562[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1080_15.INIT0 = 16'h74b8;
    defparam add_1080_15.INIT1 = 16'h74b8;
    defparam add_1080_15.INJECT1_0 = "NO";
    defparam add_1080_15.INJECT1_1 = "NO";
    CCU2D add_1075_23 (.A0(d2[56]), .B0(n5188), .C0(n5189[20]), .D0(d1[56]), 
          .A1(d2[57]), .B1(n5188), .C1(n5189[21]), .D1(d1[57]), .CIN(n12017), 
          .COUT(n12018), .S0(d2_71__N_490[56]), .S1(d2_71__N_490[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1075_23.INIT0 = 16'h74b8;
    defparam add_1075_23.INIT1 = 16'h74b8;
    defparam add_1075_23.INJECT1_0 = "NO";
    defparam add_1075_23.INJECT1_1 = "NO";
    CCU2D add_1075_21 (.A0(d2[54]), .B0(n5188), .C0(n5189[18]), .D0(d1[54]), 
          .A1(d2[55]), .B1(n5188), .C1(n5189[19]), .D1(d1[55]), .CIN(n12016), 
          .COUT(n12017), .S0(d2_71__N_490[54]), .S1(d2_71__N_490[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1075_21.INIT0 = 16'h74b8;
    defparam add_1075_21.INIT1 = 16'h74b8;
    defparam add_1075_21.INJECT1_0 = "NO";
    defparam add_1075_21.INJECT1_1 = "NO";
    CCU2D add_1075_15 (.A0(d2[48]), .B0(n5188), .C0(n5189[12]), .D0(d1[48]), 
          .A1(d2[49]), .B1(n5188), .C1(n5189[13]), .D1(d1[49]), .CIN(n12013), 
          .COUT(n12014), .S0(d2_71__N_490[48]), .S1(d2_71__N_490[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1075_15.INIT0 = 16'h74b8;
    defparam add_1075_15.INIT1 = 16'h74b8;
    defparam add_1075_15.INJECT1_0 = "NO";
    defparam add_1075_15.INJECT1_1 = "NO";
    CCU2D add_1075_9 (.A0(d2[42]), .B0(n5188), .C0(n5189[6]), .D0(d1[42]), 
          .A1(d2[43]), .B1(n5188), .C1(n5189[7]), .D1(d1[43]), .CIN(n12010), 
          .COUT(n12011), .S0(d2_71__N_490[42]), .S1(d2_71__N_490[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1075_9.INIT0 = 16'h74b8;
    defparam add_1075_9.INIT1 = 16'h74b8;
    defparam add_1075_9.INJECT1_0 = "NO";
    defparam add_1075_9.INJECT1_1 = "NO";
    CCU2D add_1075_13 (.A0(d2[46]), .B0(n5188), .C0(n5189[10]), .D0(d1[46]), 
          .A1(d2[47]), .B1(n5188), .C1(n5189[11]), .D1(d1[47]), .CIN(n12012), 
          .COUT(n12013), .S0(d2_71__N_490[46]), .S1(d2_71__N_490[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1075_13.INIT0 = 16'h74b8;
    defparam add_1075_13.INIT1 = 16'h74b8;
    defparam add_1075_13.INJECT1_0 = "NO";
    defparam add_1075_13.INJECT1_1 = "NO";
    CCU2D add_1075_19 (.A0(d2[52]), .B0(n5188), .C0(n5189[16]), .D0(d1[52]), 
          .A1(d2[53]), .B1(n5188), .C1(n5189[17]), .D1(d1[53]), .CIN(n12015), 
          .COUT(n12016), .S0(d2_71__N_490[52]), .S1(d2_71__N_490[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1075_19.INIT0 = 16'h74b8;
    defparam add_1075_19.INIT1 = 16'h74b8;
    defparam add_1075_19.INJECT1_0 = "NO";
    defparam add_1075_19.INJECT1_1 = "NO";
    CCU2D add_1075_11 (.A0(d2[44]), .B0(n5188), .C0(n5189[8]), .D0(d1[44]), 
          .A1(d2[45]), .B1(n5188), .C1(n5189[9]), .D1(d1[45]), .CIN(n12011), 
          .COUT(n12012), .S0(d2_71__N_490[44]), .S1(d2_71__N_490[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1075_11.INIT0 = 16'h74b8;
    defparam add_1075_11.INIT1 = 16'h74b8;
    defparam add_1075_11.INJECT1_0 = "NO";
    defparam add_1075_11.INJECT1_1 = "NO";
    CCU2D add_1075_7 (.A0(d2[40]), .B0(n5188), .C0(n5189[4]), .D0(d1[40]), 
          .A1(d2[41]), .B1(n5188), .C1(n5189[5]), .D1(d1[41]), .CIN(n12009), 
          .COUT(n12010), .S0(d2_71__N_490[40]), .S1(d2_71__N_490[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1075_7.INIT0 = 16'h74b8;
    defparam add_1075_7.INIT1 = 16'h74b8;
    defparam add_1075_7.INJECT1_0 = "NO";
    defparam add_1075_7.INJECT1_1 = "NO";
    CCU2D add_1075_17 (.A0(d2[50]), .B0(n5188), .C0(n5189[14]), .D0(d1[50]), 
          .A1(d2[51]), .B1(n5188), .C1(n5189[15]), .D1(d1[51]), .CIN(n12014), 
          .COUT(n12015), .S0(d2_71__N_490[50]), .S1(d2_71__N_490[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1075_17.INIT0 = 16'h74b8;
    defparam add_1075_17.INIT1 = 16'h74b8;
    defparam add_1075_17.INJECT1_0 = "NO";
    defparam add_1075_17.INJECT1_1 = "NO";
    CCU2D add_1080_13 (.A0(d3[46]), .B0(n5340), .C0(n5341[10]), .D0(d2[46]), 
          .A1(d3[47]), .B1(n5340), .C1(n5341[11]), .D1(d2[47]), .CIN(n11971), 
          .COUT(n11972), .S0(d3_71__N_562[46]), .S1(d3_71__N_562[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1080_13.INIT0 = 16'h74b8;
    defparam add_1080_13.INIT1 = 16'h74b8;
    defparam add_1080_13.INJECT1_0 = "NO";
    defparam add_1080_13.INJECT1_1 = "NO";
    CCU2D add_1080_11 (.A0(d3[44]), .B0(n5340), .C0(n5341[8]), .D0(d2[44]), 
          .A1(d3[45]), .B1(n5340), .C1(n5341[9]), .D1(d2[45]), .CIN(n11970), 
          .COUT(n11971), .S0(d3_71__N_562[44]), .S1(d3_71__N_562[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1080_11.INIT0 = 16'h74b8;
    defparam add_1080_11.INIT1 = 16'h74b8;
    defparam add_1080_11.INJECT1_0 = "NO";
    defparam add_1080_11.INJECT1_1 = "NO";
    CCU2D add_1089_10 (.A0(d4[44]), .B0(d5[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[45]), .B1(d5[45]), .C1(GND_net), .D1(GND_net), .CIN(n11907), 
          .COUT(n11908), .S0(n5645[8]), .S1(n5645[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1089_10.INIT0 = 16'h5666;
    defparam add_1089_10.INIT1 = 16'h5666;
    defparam add_1089_10.INJECT1_0 = "NO";
    defparam add_1089_10.INJECT1_1 = "NO";
    CCU2D add_1104_37 (.A0(d_tmp[71]), .B0(d_d_tmp[71]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11623), .S0(n6101[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1104_37.INIT0 = 16'h5999;
    defparam add_1104_37.INIT1 = 16'h0000;
    defparam add_1104_37.INJECT1_0 = "NO";
    defparam add_1104_37.INJECT1_1 = "NO";
    FD1S3IX count__i0 (.D(count_15__N_1442[0]), .CK(osc_clk), .CD(osc_clk_enable_744), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i0.GSR = "ENABLED";
    CCU2D add_1080_9 (.A0(d3[42]), .B0(n5340), .C0(n5341[6]), .D0(d2[42]), 
          .A1(d3[43]), .B1(n5340), .C1(n5341[7]), .D1(d2[43]), .CIN(n11969), 
          .COUT(n11970), .S0(d3_71__N_562[42]), .S1(d3_71__N_562[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1080_9.INIT0 = 16'h74b8;
    defparam add_1080_9.INIT1 = 16'h74b8;
    defparam add_1080_9.INJECT1_0 = "NO";
    defparam add_1080_9.INJECT1_1 = "NO";
    CCU2D add_1080_7 (.A0(d3[40]), .B0(n5340), .C0(n5341[4]), .D0(d2[40]), 
          .A1(d3[41]), .B1(n5340), .C1(n5341[5]), .D1(d2[41]), .CIN(n11968), 
          .COUT(n11969), .S0(d3_71__N_562[40]), .S1(d3_71__N_562[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1080_7.INIT0 = 16'h74b8;
    defparam add_1080_7.INIT1 = 16'h74b8;
    defparam add_1080_7.INJECT1_0 = "NO";
    defparam add_1080_7.INJECT1_1 = "NO";
    CCU2D add_1080_5 (.A0(d3[38]), .B0(n5340), .C0(n5341[2]), .D0(d2[38]), 
          .A1(d3[39]), .B1(n5340), .C1(n5341[3]), .D1(d2[39]), .CIN(n11967), 
          .COUT(n11968), .S0(d3_71__N_562[38]), .S1(d3_71__N_562[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1080_5.INIT0 = 16'h74b8;
    defparam add_1080_5.INIT1 = 16'h74b8;
    defparam add_1080_5.INJECT1_0 = "NO";
    defparam add_1080_5.INJECT1_1 = "NO";
    CCU2D add_1089_8 (.A0(d4[42]), .B0(d5[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[43]), .B1(d5[43]), .C1(GND_net), .D1(GND_net), .CIN(n11906), 
          .COUT(n11907), .S0(n5645[6]), .S1(n5645[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1089_8.INIT0 = 16'h5666;
    defparam add_1089_8.INIT1 = 16'h5666;
    defparam add_1089_8.INJECT1_0 = "NO";
    defparam add_1089_8.INJECT1_1 = "NO";
    CCU2D add_1080_3 (.A0(d3[36]), .B0(n5340), .C0(n5341[0]), .D0(d2[36]), 
          .A1(d3[37]), .B1(n5340), .C1(n5341[1]), .D1(d2[37]), .CIN(n11966), 
          .COUT(n11967), .S0(d3_71__N_562[36]), .S1(d3_71__N_562[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1080_3.INIT0 = 16'h74b8;
    defparam add_1080_3.INIT1 = 16'h74b8;
    defparam add_1080_3.INJECT1_0 = "NO";
    defparam add_1080_3.INJECT1_1 = "NO";
    CCU2D add_1089_6 (.A0(d4[40]), .B0(d5[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[41]), .B1(d5[41]), .C1(GND_net), .D1(GND_net), .CIN(n11905), 
          .COUT(n11906), .S0(n5645[4]), .S1(n5645[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1089_6.INIT0 = 16'h5666;
    defparam add_1089_6.INIT1 = 16'h5666;
    defparam add_1089_6.INJECT1_0 = "NO";
    defparam add_1089_6.INJECT1_1 = "NO";
    CCU2D add_1075_5 (.A0(d2[38]), .B0(n5188), .C0(n5189[2]), .D0(d1[38]), 
          .A1(d2[39]), .B1(n5188), .C1(n5189[3]), .D1(d1[39]), .CIN(n12008), 
          .COUT(n12009), .S0(d2_71__N_490[38]), .S1(d2_71__N_490[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1075_5.INIT0 = 16'h74b8;
    defparam add_1075_5.INIT1 = 16'h74b8;
    defparam add_1075_5.INJECT1_0 = "NO";
    defparam add_1075_5.INJECT1_1 = "NO";
    CCU2D add_1079_36 (.A0(d2[70]), .B0(d3[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[71]), .B1(d3[71]), .C1(GND_net), .D1(GND_net), .CIN(n12002), 
          .S0(n5341[34]), .S1(n5341[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1079_36.INIT0 = 16'h5666;
    defparam add_1079_36.INIT1 = 16'h5666;
    defparam add_1079_36.INJECT1_0 = "NO";
    defparam add_1079_36.INJECT1_1 = "NO";
    CCU2D add_1090_23 (.A0(d5[56]), .B0(n5644), .C0(n5645[20]), .D0(d4[56]), 
          .A1(d5[57]), .B1(n5644), .C1(n5645[21]), .D1(d4[57]), .CIN(n11894), 
          .COUT(n11895), .S0(d5_71__N_706[56]), .S1(d5_71__N_706[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1090_23.INIT0 = 16'h74b8;
    defparam add_1090_23.INIT1 = 16'h74b8;
    defparam add_1090_23.INJECT1_0 = "NO";
    defparam add_1090_23.INJECT1_1 = "NO";
    CCU2D add_1079_16 (.A0(d2[50]), .B0(d3[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[51]), .B1(d3[51]), .C1(GND_net), .D1(GND_net), .CIN(n11992), 
          .COUT(n11993), .S0(n5341[14]), .S1(n5341[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1079_16.INIT0 = 16'h5666;
    defparam add_1079_16.INIT1 = 16'h5666;
    defparam add_1079_16.INJECT1_0 = "NO";
    defparam add_1079_16.INJECT1_1 = "NO";
    CCU2D add_1079_14 (.A0(d2[48]), .B0(d3[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[49]), .B1(d3[49]), .C1(GND_net), .D1(GND_net), .CIN(n11991), 
          .COUT(n11992), .S0(n5341[12]), .S1(n5341[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1079_14.INIT0 = 16'h5666;
    defparam add_1079_14.INIT1 = 16'h5666;
    defparam add_1079_14.INJECT1_0 = "NO";
    defparam add_1079_14.INJECT1_1 = "NO";
    CCU2D add_1079_12 (.A0(d2[46]), .B0(d3[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[47]), .B1(d3[47]), .C1(GND_net), .D1(GND_net), .CIN(n11990), 
          .COUT(n11991), .S0(n5341[10]), .S1(n5341[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1079_12.INIT0 = 16'h5666;
    defparam add_1079_12.INIT1 = 16'h5666;
    defparam add_1079_12.INJECT1_0 = "NO";
    defparam add_1079_12.INJECT1_1 = "NO";
    CCU2D add_1079_8 (.A0(d2[42]), .B0(d3[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[43]), .B1(d3[43]), .C1(GND_net), .D1(GND_net), .CIN(n11988), 
          .COUT(n11989), .S0(n5341[6]), .S1(n5341[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1079_8.INIT0 = 16'h5666;
    defparam add_1079_8.INIT1 = 16'h5666;
    defparam add_1079_8.INJECT1_0 = "NO";
    defparam add_1079_8.INJECT1_1 = "NO";
    CCU2D add_1079_6 (.A0(d2[40]), .B0(d3[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[41]), .B1(d3[41]), .C1(GND_net), .D1(GND_net), .CIN(n11987), 
          .COUT(n11988), .S0(n5341[4]), .S1(n5341[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1079_6.INIT0 = 16'h5666;
    defparam add_1079_6.INIT1 = 16'h5666;
    defparam add_1079_6.INJECT1_0 = "NO";
    defparam add_1079_6.INJECT1_1 = "NO";
    CCU2D add_1089_4 (.A0(d4[38]), .B0(d5[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[39]), .B1(d5[39]), .C1(GND_net), .D1(GND_net), .CIN(n11904), 
          .COUT(n11905), .S0(n5645[2]), .S1(n5645[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1089_4.INIT0 = 16'h5666;
    defparam add_1089_4.INIT1 = 16'h5666;
    defparam add_1089_4.INJECT1_0 = "NO";
    defparam add_1089_4.INJECT1_1 = "NO";
    CCU2D add_1079_10 (.A0(d2[44]), .B0(d3[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[45]), .B1(d3[45]), .C1(GND_net), .D1(GND_net), .CIN(n11989), 
          .COUT(n11990), .S0(n5341[8]), .S1(n5341[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1079_10.INIT0 = 16'h5666;
    defparam add_1079_10.INIT1 = 16'h5666;
    defparam add_1079_10.INJECT1_0 = "NO";
    defparam add_1079_10.INJECT1_1 = "NO";
    LUT4 i2851_2_lut (.A(n375[0]), .B(n31), .Z(count_15__N_1442[0])) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(86[13] 89[16])
    defparam i2851_2_lut.init = 16'hbbbb;
    LUT4 i4912_2_lut (.A(MixerOutCos[0]), .B(d1[0]), .Z(d1_71__N_418[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4912_2_lut.init = 16'h6666;
    CCU2D add_1079_4 (.A0(d2[38]), .B0(d3[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[39]), .B1(d3[39]), .C1(GND_net), .D1(GND_net), .CIN(n11986), 
          .COUT(n11987), .S0(n5341[2]), .S1(n5341[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1079_4.INIT0 = 16'h5666;
    defparam add_1079_4.INIT1 = 16'h5666;
    defparam add_1079_4.INJECT1_0 = "NO";
    defparam add_1079_4.INJECT1_1 = "NO";
    CCU2D add_1080_37 (.A0(d3[70]), .B0(n5340), .C0(n5341[34]), .D0(d2[70]), 
          .A1(d3[71]), .B1(n5340), .C1(n5341[35]), .D1(d2[71]), .CIN(n11983), 
          .S0(d3_71__N_562[70]), .S1(d3_71__N_562[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1080_37.INIT0 = 16'h74b8;
    defparam add_1080_37.INIT1 = 16'h74b8;
    defparam add_1080_37.INJECT1_0 = "NO";
    defparam add_1080_37.INJECT1_1 = "NO";
    CCU2D add_1080_25 (.A0(d3[58]), .B0(n5340), .C0(n5341[22]), .D0(d2[58]), 
          .A1(d3[59]), .B1(n5340), .C1(n5341[23]), .D1(d2[59]), .CIN(n11977), 
          .COUT(n11978), .S0(d3_71__N_562[58]), .S1(d3_71__N_562[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1080_25.INIT0 = 16'h74b8;
    defparam add_1080_25.INIT1 = 16'h74b8;
    defparam add_1080_25.INJECT1_0 = "NO";
    defparam add_1080_25.INJECT1_1 = "NO";
    CCU2D add_1080_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5340), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11966));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1080_1.INIT0 = 16'hF000;
    defparam add_1080_1.INIT1 = 16'h0555;
    defparam add_1080_1.INJECT1_0 = "NO";
    defparam add_1080_1.INJECT1_1 = "NO";
    CCU2D add_1080_35 (.A0(d3[68]), .B0(n5340), .C0(n5341[32]), .D0(d2[68]), 
          .A1(d3[69]), .B1(n5340), .C1(n5341[33]), .D1(d2[69]), .CIN(n11982), 
          .COUT(n11983), .S0(d3_71__N_562[68]), .S1(d3_71__N_562[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1080_35.INIT0 = 16'h74b8;
    defparam add_1080_35.INIT1 = 16'h74b8;
    defparam add_1080_35.INJECT1_0 = "NO";
    defparam add_1080_35.INJECT1_1 = "NO";
    CCU2D add_1080_33 (.A0(d3[66]), .B0(n5340), .C0(n5341[30]), .D0(d2[66]), 
          .A1(d3[67]), .B1(n5340), .C1(n5341[31]), .D1(d2[67]), .CIN(n11981), 
          .COUT(n11982), .S0(d3_71__N_562[66]), .S1(d3_71__N_562[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1080_33.INIT0 = 16'h74b8;
    defparam add_1080_33.INIT1 = 16'h74b8;
    defparam add_1080_33.INJECT1_0 = "NO";
    defparam add_1080_33.INJECT1_1 = "NO";
    CCU2D add_1079_2 (.A0(d2[36]), .B0(d3[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[37]), .B1(d3[37]), .C1(GND_net), .D1(GND_net), .COUT(n11986), 
          .S1(n5341[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1079_2.INIT0 = 16'h7000;
    defparam add_1079_2.INIT1 = 16'h5666;
    defparam add_1079_2.INJECT1_0 = "NO";
    defparam add_1079_2.INJECT1_1 = "NO";
    CCU2D add_1080_31 (.A0(d3[64]), .B0(n5340), .C0(n5341[28]), .D0(d2[64]), 
          .A1(d3[65]), .B1(n5340), .C1(n5341[29]), .D1(d2[65]), .CIN(n11980), 
          .COUT(n11981), .S0(d3_71__N_562[64]), .S1(d3_71__N_562[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1080_31.INIT0 = 16'h74b8;
    defparam add_1080_31.INIT1 = 16'h74b8;
    defparam add_1080_31.INJECT1_0 = "NO";
    defparam add_1080_31.INJECT1_1 = "NO";
    CCU2D add_1080_29 (.A0(d3[62]), .B0(n5340), .C0(n5341[26]), .D0(d2[62]), 
          .A1(d3[63]), .B1(n5340), .C1(n5341[27]), .D1(d2[63]), .CIN(n11979), 
          .COUT(n11980), .S0(d3_71__N_562[62]), .S1(d3_71__N_562[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1080_29.INIT0 = 16'h74b8;
    defparam add_1080_29.INIT1 = 16'h74b8;
    defparam add_1080_29.INJECT1_0 = "NO";
    defparam add_1080_29.INJECT1_1 = "NO";
    CCU2D add_1080_27 (.A0(d3[60]), .B0(n5340), .C0(n5341[24]), .D0(d2[60]), 
          .A1(d3[61]), .B1(n5340), .C1(n5341[25]), .D1(d2[61]), .CIN(n11978), 
          .COUT(n11979), .S0(d3_71__N_562[60]), .S1(d3_71__N_562[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1080_27.INIT0 = 16'h74b8;
    defparam add_1080_27.INIT1 = 16'h74b8;
    defparam add_1080_27.INJECT1_0 = "NO";
    defparam add_1080_27.INJECT1_1 = "NO";
    CCU2D add_1090_21 (.A0(d5[54]), .B0(n5644), .C0(n5645[18]), .D0(d4[54]), 
          .A1(d5[55]), .B1(n5644), .C1(n5645[19]), .D1(d4[55]), .CIN(n11893), 
          .COUT(n11894), .S0(d5_71__N_706[54]), .S1(d5_71__N_706[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1090_21.INIT0 = 16'h74b8;
    defparam add_1090_21.INIT1 = 16'h74b8;
    defparam add_1090_21.INJECT1_0 = "NO";
    defparam add_1090_21.INJECT1_1 = "NO";
    CCU2D add_1075_31 (.A0(d2[64]), .B0(n5188), .C0(n5189[28]), .D0(d1[64]), 
          .A1(d2[65]), .B1(n5188), .C1(n5189[29]), .D1(d1[65]), .CIN(n12021), 
          .COUT(n12022), .S0(d2_71__N_490[64]), .S1(d2_71__N_490[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1075_31.INIT0 = 16'h74b8;
    defparam add_1075_31.INIT1 = 16'h74b8;
    defparam add_1075_31.INJECT1_0 = "NO";
    defparam add_1075_31.INJECT1_1 = "NO";
    CCU2D add_1074_14 (.A0(d1[48]), .B0(d2[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[49]), .B1(d2[49]), .C1(GND_net), .D1(GND_net), .CIN(n12032), 
          .COUT(n12033), .S0(n5189[12]), .S1(n5189[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1074_14.INIT0 = 16'h5666;
    defparam add_1074_14.INIT1 = 16'h5666;
    defparam add_1074_14.INJECT1_0 = "NO";
    defparam add_1074_14.INJECT1_1 = "NO";
    LUT4 i11_4_lut (.A(n21), .B(n19), .C(n15), .D(n16), .Z(n31)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i9_4_lut (.A(count[9]), .B(count[3]), .C(count[4]), .D(count[0]), 
         .Z(n21)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i9_4_lut.init = 16'hfffe;
    CCU2D add_1090_19 (.A0(d5[52]), .B0(n5644), .C0(n5645[16]), .D0(d4[52]), 
          .A1(d5[53]), .B1(n5644), .C1(n5645[17]), .D1(d4[53]), .CIN(n11892), 
          .COUT(n11893), .S0(d5_71__N_706[52]), .S1(d5_71__N_706[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1090_19.INIT0 = 16'h74b8;
    defparam add_1090_19.INIT1 = 16'h74b8;
    defparam add_1090_19.INJECT1_0 = "NO";
    defparam add_1090_19.INJECT1_1 = "NO";
    CCU2D add_1090_17 (.A0(d5[50]), .B0(n5644), .C0(n5645[14]), .D0(d4[50]), 
          .A1(d5[51]), .B1(n5644), .C1(n5645[15]), .D1(d4[51]), .CIN(n11891), 
          .COUT(n11892), .S0(d5_71__N_706[50]), .S1(d5_71__N_706[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1090_17.INIT0 = 16'h74b8;
    defparam add_1090_17.INIT1 = 16'h74b8;
    defparam add_1090_17.INJECT1_0 = "NO";
    defparam add_1090_17.INJECT1_1 = "NO";
    CCU2D add_1090_15 (.A0(d5[48]), .B0(n5644), .C0(n5645[12]), .D0(d4[48]), 
          .A1(d5[49]), .B1(n5644), .C1(n5645[13]), .D1(d4[49]), .CIN(n11890), 
          .COUT(n11891), .S0(d5_71__N_706[48]), .S1(d5_71__N_706[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1090_15.INIT0 = 16'h74b8;
    defparam add_1090_15.INIT1 = 16'h74b8;
    defparam add_1090_15.INJECT1_0 = "NO";
    defparam add_1090_15.INJECT1_1 = "NO";
    CCU2D add_1090_13 (.A0(d5[46]), .B0(n5644), .C0(n5645[10]), .D0(d4[46]), 
          .A1(d5[47]), .B1(n5644), .C1(n5645[11]), .D1(d4[47]), .CIN(n11889), 
          .COUT(n11890), .S0(d5_71__N_706[46]), .S1(d5_71__N_706[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1090_13.INIT0 = 16'h74b8;
    defparam add_1090_13.INIT1 = 16'h74b8;
    defparam add_1090_13.INJECT1_0 = "NO";
    defparam add_1090_13.INJECT1_1 = "NO";
    CCU2D add_1090_11 (.A0(d5[44]), .B0(n5644), .C0(n5645[8]), .D0(d4[44]), 
          .A1(d5[45]), .B1(n5644), .C1(n5645[9]), .D1(d4[45]), .CIN(n11888), 
          .COUT(n11889), .S0(d5_71__N_706[44]), .S1(d5_71__N_706[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1090_11.INIT0 = 16'h74b8;
    defparam add_1090_11.INIT1 = 16'h74b8;
    defparam add_1090_11.INJECT1_0 = "NO";
    defparam add_1090_11.INJECT1_1 = "NO";
    CCU2D add_1090_9 (.A0(d5[42]), .B0(n5644), .C0(n5645[6]), .D0(d4[42]), 
          .A1(d5[43]), .B1(n5644), .C1(n5645[7]), .D1(d4[43]), .CIN(n11887), 
          .COUT(n11888), .S0(d5_71__N_706[42]), .S1(d5_71__N_706[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1090_9.INIT0 = 16'h74b8;
    defparam add_1090_9.INIT1 = 16'h74b8;
    defparam add_1090_9.INJECT1_0 = "NO";
    defparam add_1090_9.INJECT1_1 = "NO";
    CCU2D add_1090_7 (.A0(d5[40]), .B0(n5644), .C0(n5645[4]), .D0(d4[40]), 
          .A1(d5[41]), .B1(n5644), .C1(n5645[5]), .D1(d4[41]), .CIN(n11886), 
          .COUT(n11887), .S0(d5_71__N_706[40]), .S1(d5_71__N_706[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1090_7.INIT0 = 16'h74b8;
    defparam add_1090_7.INIT1 = 16'h74b8;
    defparam add_1090_7.INJECT1_0 = "NO";
    defparam add_1090_7.INJECT1_1 = "NO";
    LUT4 i7_4_lut (.A(count[10]), .B(count[1]), .C(count[5]), .D(count[6]), 
         .Z(n19)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i7_4_lut.init = 16'hfffe;
    CCU2D add_1090_5 (.A0(d5[38]), .B0(n5644), .C0(n5645[2]), .D0(d4[38]), 
          .A1(d5[39]), .B1(n5644), .C1(n5645[3]), .D1(d4[39]), .CIN(n11885), 
          .COUT(n11886), .S0(d5_71__N_706[38]), .S1(d5_71__N_706[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1090_5.INIT0 = 16'h74b8;
    defparam add_1090_5.INIT1 = 16'h74b8;
    defparam add_1090_5.INJECT1_0 = "NO";
    defparam add_1090_5.INJECT1_1 = "NO";
    CCU2D add_1090_3 (.A0(d5[36]), .B0(n5644), .C0(n5645[0]), .D0(d4[36]), 
          .A1(d5[37]), .B1(n5644), .C1(n5645[1]), .D1(d4[37]), .CIN(n11884), 
          .COUT(n11885), .S0(d5_71__N_706[36]), .S1(d5_71__N_706[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1090_3.INIT0 = 16'h74b8;
    defparam add_1090_3.INIT1 = 16'h74b8;
    defparam add_1090_3.INJECT1_0 = "NO";
    defparam add_1090_3.INJECT1_1 = "NO";
    CCU2D add_1090_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5644), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11884));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1090_1.INIT0 = 16'hF000;
    defparam add_1090_1.INIT1 = 16'h0555;
    defparam add_1090_1.INJECT1_0 = "NO";
    defparam add_1090_1.INJECT1_1 = "NO";
    CCU2D add_1074_12 (.A0(d1[46]), .B0(d2[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[47]), .B1(d2[47]), .C1(GND_net), .D1(GND_net), .CIN(n12031), 
          .COUT(n12032), .S0(n5189[10]), .S1(n5189[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1074_12.INIT0 = 16'h5666;
    defparam add_1074_12.INIT1 = 16'h5666;
    defparam add_1074_12.INJECT1_0 = "NO";
    defparam add_1074_12.INJECT1_1 = "NO";
    CCU2D add_1074_10 (.A0(d1[44]), .B0(d2[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[45]), .B1(d2[45]), .C1(GND_net), .D1(GND_net), .CIN(n12030), 
          .COUT(n12031), .S0(n5189[8]), .S1(n5189[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1074_10.INIT0 = 16'h5666;
    defparam add_1074_10.INIT1 = 16'h5666;
    defparam add_1074_10.INJECT1_0 = "NO";
    defparam add_1074_10.INJECT1_1 = "NO";
    CCU2D add_1074_8 (.A0(d1[42]), .B0(d2[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[43]), .B1(d2[43]), .C1(GND_net), .D1(GND_net), .CIN(n12029), 
          .COUT(n12030), .S0(n5189[6]), .S1(n5189[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1074_8.INIT0 = 16'h5666;
    defparam add_1074_8.INIT1 = 16'h5666;
    defparam add_1074_8.INJECT1_0 = "NO";
    defparam add_1074_8.INJECT1_1 = "NO";
    CCU2D add_1074_4 (.A0(d1[38]), .B0(d2[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[39]), .B1(d2[39]), .C1(GND_net), .D1(GND_net), .CIN(n12027), 
          .COUT(n12028), .S0(n5189[2]), .S1(n5189[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1074_4.INIT0 = 16'h5666;
    defparam add_1074_4.INIT1 = 16'h5666;
    defparam add_1074_4.INJECT1_0 = "NO";
    defparam add_1074_4.INJECT1_1 = "NO";
    CCU2D add_1089_2 (.A0(d4[36]), .B0(d5[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[37]), .B1(d5[37]), .C1(GND_net), .D1(GND_net), .COUT(n11904), 
          .S1(n5645[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1089_2.INIT0 = 16'h7000;
    defparam add_1089_2.INIT1 = 16'h5666;
    defparam add_1089_2.INJECT1_0 = "NO";
    defparam add_1089_2.INJECT1_1 = "NO";
    CCU2D add_1074_2 (.A0(d1[36]), .B0(d2[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[37]), .B1(d2[37]), .C1(GND_net), .D1(GND_net), .COUT(n12027), 
          .S1(n5189[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1074_2.INIT0 = 16'h7000;
    defparam add_1074_2.INIT1 = 16'h5666;
    defparam add_1074_2.INJECT1_0 = "NO";
    defparam add_1074_2.INJECT1_1 = "NO";
    CCU2D add_1075_37 (.A0(d2[70]), .B0(n5188), .C0(n5189[34]), .D0(d1[70]), 
          .A1(d2[71]), .B1(n5188), .C1(n5189[35]), .D1(d1[71]), .CIN(n12024), 
          .S0(d2_71__N_490[70]), .S1(d2_71__N_490[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1075_37.INIT0 = 16'h74b8;
    defparam add_1075_37.INIT1 = 16'h74b8;
    defparam add_1075_37.INJECT1_0 = "NO";
    defparam add_1075_37.INJECT1_1 = "NO";
    CCU2D add_1075_35 (.A0(d2[68]), .B0(n5188), .C0(n5189[32]), .D0(d1[68]), 
          .A1(d2[69]), .B1(n5188), .C1(n5189[33]), .D1(d1[69]), .CIN(n12023), 
          .COUT(n12024), .S0(d2_71__N_490[68]), .S1(d2_71__N_490[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1075_35.INIT0 = 16'h74b8;
    defparam add_1075_35.INIT1 = 16'h74b8;
    defparam add_1075_35.INJECT1_0 = "NO";
    defparam add_1075_35.INJECT1_1 = "NO";
    CCU2D add_1104_35 (.A0(d_tmp[69]), .B0(d_d_tmp[69]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[70]), .B1(d_d_tmp[70]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11622), .COUT(n11623), .S0(n6101[33]), 
          .S1(n6101[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1104_35.INIT0 = 16'h5999;
    defparam add_1104_35.INIT1 = 16'h5999;
    defparam add_1104_35.INJECT1_0 = "NO";
    defparam add_1104_35.INJECT1_1 = "NO";
    CCU2D add_1104_33 (.A0(d_tmp[67]), .B0(d_d_tmp[67]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[68]), .B1(d_d_tmp[68]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11621), .COUT(n11622), .S0(n6101[31]), 
          .S1(n6101[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1104_33.INIT0 = 16'h5999;
    defparam add_1104_33.INIT1 = 16'h5999;
    defparam add_1104_33.INJECT1_0 = "NO";
    defparam add_1104_33.INJECT1_1 = "NO";
    CCU2D add_1104_31 (.A0(d_tmp[65]), .B0(d_d_tmp[65]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[66]), .B1(d_d_tmp[66]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11620), .COUT(n11621), .S0(n6101[29]), 
          .S1(n6101[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1104_31.INIT0 = 16'h5999;
    defparam add_1104_31.INIT1 = 16'h5999;
    defparam add_1104_31.INJECT1_0 = "NO";
    defparam add_1104_31.INJECT1_1 = "NO";
    CCU2D add_1104_29 (.A0(d_tmp[63]), .B0(d_d_tmp[63]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[64]), .B1(d_d_tmp[64]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11619), .COUT(n11620), .S0(n6101[27]), 
          .S1(n6101[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1104_29.INIT0 = 16'h5999;
    defparam add_1104_29.INIT1 = 16'h5999;
    defparam add_1104_29.INJECT1_0 = "NO";
    defparam add_1104_29.INJECT1_1 = "NO";
    CCU2D add_1104_27 (.A0(d_tmp[61]), .B0(d_d_tmp[61]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[62]), .B1(d_d_tmp[62]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11618), .COUT(n11619), .S0(n6101[25]), 
          .S1(n6101[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1104_27.INIT0 = 16'h5999;
    defparam add_1104_27.INIT1 = 16'h5999;
    defparam add_1104_27.INJECT1_0 = "NO";
    defparam add_1104_27.INJECT1_1 = "NO";
    CCU2D add_1104_25 (.A0(d_tmp[59]), .B0(d_d_tmp[59]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[60]), .B1(d_d_tmp[60]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11617), .COUT(n11618), .S0(n6101[23]), 
          .S1(n6101[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1104_25.INIT0 = 16'h5999;
    defparam add_1104_25.INIT1 = 16'h5999;
    defparam add_1104_25.INJECT1_0 = "NO";
    defparam add_1104_25.INJECT1_1 = "NO";
    CCU2D add_1104_23 (.A0(d_tmp[57]), .B0(d_d_tmp[57]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[58]), .B1(d_d_tmp[58]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11616), .COUT(n11617), .S0(n6101[21]), 
          .S1(n6101[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1104_23.INIT0 = 16'h5999;
    defparam add_1104_23.INIT1 = 16'h5999;
    defparam add_1104_23.INJECT1_0 = "NO";
    defparam add_1104_23.INJECT1_1 = "NO";
    CCU2D add_1104_21 (.A0(d_tmp[55]), .B0(d_d_tmp[55]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[56]), .B1(d_d_tmp[56]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11615), .COUT(n11616), .S0(n6101[19]), 
          .S1(n6101[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1104_21.INIT0 = 16'h5999;
    defparam add_1104_21.INIT1 = 16'h5999;
    defparam add_1104_21.INJECT1_0 = "NO";
    defparam add_1104_21.INJECT1_1 = "NO";
    CCU2D add_1104_19 (.A0(d_tmp[53]), .B0(d_d_tmp[53]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[54]), .B1(d_d_tmp[54]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11614), .COUT(n11615), .S0(n6101[17]), 
          .S1(n6101[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1104_19.INIT0 = 16'h5999;
    defparam add_1104_19.INIT1 = 16'h5999;
    defparam add_1104_19.INJECT1_0 = "NO";
    defparam add_1104_19.INJECT1_1 = "NO";
    CCU2D add_1079_24 (.A0(d2[58]), .B0(d3[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[59]), .B1(d3[59]), .C1(GND_net), .D1(GND_net), .CIN(n11996), 
          .COUT(n11997), .S0(n5341[22]), .S1(n5341[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1079_24.INIT0 = 16'h5666;
    defparam add_1079_24.INIT1 = 16'h5666;
    defparam add_1079_24.INJECT1_0 = "NO";
    defparam add_1079_24.INJECT1_1 = "NO";
    CCU2D add_1104_17 (.A0(d_tmp[51]), .B0(d_d_tmp[51]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[52]), .B1(d_d_tmp[52]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11613), .COUT(n11614), .S0(n6101[15]), 
          .S1(n6101[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1104_17.INIT0 = 16'h5999;
    defparam add_1104_17.INIT1 = 16'h5999;
    defparam add_1104_17.INJECT1_0 = "NO";
    defparam add_1104_17.INJECT1_1 = "NO";
    CCU2D add_1104_15 (.A0(d_tmp[49]), .B0(d_d_tmp[49]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[50]), .B1(d_d_tmp[50]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11612), .COUT(n11613), .S0(n6101[13]), 
          .S1(n6101[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1104_15.INIT0 = 16'h5999;
    defparam add_1104_15.INIT1 = 16'h5999;
    defparam add_1104_15.INJECT1_0 = "NO";
    defparam add_1104_15.INJECT1_1 = "NO";
    CCU2D add_1104_13 (.A0(d_tmp[47]), .B0(d_d_tmp[47]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[48]), .B1(d_d_tmp[48]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11611), .COUT(n11612), .S0(n6101[11]), 
          .S1(n6101[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1104_13.INIT0 = 16'h5999;
    defparam add_1104_13.INIT1 = 16'h5999;
    defparam add_1104_13.INJECT1_0 = "NO";
    defparam add_1104_13.INJECT1_1 = "NO";
    CCU2D add_1084_36 (.A0(d3[70]), .B0(d4[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[71]), .B1(d4[71]), .C1(GND_net), .D1(GND_net), .CIN(n11961), 
          .S0(n5493[34]), .S1(n5493[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1084_36.INIT0 = 16'h5666;
    defparam add_1084_36.INIT1 = 16'h5666;
    defparam add_1084_36.INJECT1_0 = "NO";
    defparam add_1084_36.INJECT1_1 = "NO";
    CCU2D add_1079_22 (.A0(d2[56]), .B0(d3[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[57]), .B1(d3[57]), .C1(GND_net), .D1(GND_net), .CIN(n11995), 
          .COUT(n11996), .S0(n5341[20]), .S1(n5341[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1079_22.INIT0 = 16'h5666;
    defparam add_1079_22.INIT1 = 16'h5666;
    defparam add_1079_22.INJECT1_0 = "NO";
    defparam add_1079_22.INJECT1_1 = "NO";
    CCU2D add_1084_34 (.A0(d3[68]), .B0(d4[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[69]), .B1(d4[69]), .C1(GND_net), .D1(GND_net), .CIN(n11960), 
          .COUT(n11961), .S0(n5493[32]), .S1(n5493[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1084_34.INIT0 = 16'h5666;
    defparam add_1084_34.INIT1 = 16'h5666;
    defparam add_1084_34.INJECT1_0 = "NO";
    defparam add_1084_34.INJECT1_1 = "NO";
    CCU2D add_1079_34 (.A0(d2[68]), .B0(d3[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[69]), .B1(d3[69]), .C1(GND_net), .D1(GND_net), .CIN(n12001), 
          .COUT(n12002), .S0(n5341[32]), .S1(n5341[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1079_34.INIT0 = 16'h5666;
    defparam add_1079_34.INIT1 = 16'h5666;
    defparam add_1079_34.INJECT1_0 = "NO";
    defparam add_1079_34.INJECT1_1 = "NO";
    CCU2D add_1079_20 (.A0(d2[54]), .B0(d3[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[55]), .B1(d3[55]), .C1(GND_net), .D1(GND_net), .CIN(n11994), 
          .COUT(n11995), .S0(n5341[18]), .S1(n5341[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1079_20.INIT0 = 16'h5666;
    defparam add_1079_20.INIT1 = 16'h5666;
    defparam add_1079_20.INJECT1_0 = "NO";
    defparam add_1079_20.INJECT1_1 = "NO";
    CCU2D add_1079_32 (.A0(d2[66]), .B0(d3[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[67]), .B1(d3[67]), .C1(GND_net), .D1(GND_net), .CIN(n12000), 
          .COUT(n12001), .S0(n5341[30]), .S1(n5341[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1079_32.INIT0 = 16'h5666;
    defparam add_1079_32.INIT1 = 16'h5666;
    defparam add_1079_32.INJECT1_0 = "NO";
    defparam add_1079_32.INJECT1_1 = "NO";
    CCU2D add_1075_3 (.A0(d2[36]), .B0(n5188), .C0(n5189[0]), .D0(d1[36]), 
          .A1(d2[37]), .B1(n5188), .C1(n5189[1]), .D1(d1[37]), .CIN(n12007), 
          .COUT(n12008), .S0(d2_71__N_490[36]), .S1(d2_71__N_490[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1075_3.INIT0 = 16'h74b8;
    defparam add_1075_3.INIT1 = 16'h74b8;
    defparam add_1075_3.INJECT1_0 = "NO";
    defparam add_1075_3.INJECT1_1 = "NO";
    CCU2D add_1079_30 (.A0(d2[64]), .B0(d3[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[65]), .B1(d3[65]), .C1(GND_net), .D1(GND_net), .CIN(n11999), 
          .COUT(n12000), .S0(n5341[28]), .S1(n5341[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1079_30.INIT0 = 16'h5666;
    defparam add_1079_30.INIT1 = 16'h5666;
    defparam add_1079_30.INJECT1_0 = "NO";
    defparam add_1079_30.INJECT1_1 = "NO";
    CCU2D add_1079_18 (.A0(d2[52]), .B0(d3[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[53]), .B1(d3[53]), .C1(GND_net), .D1(GND_net), .CIN(n11993), 
          .COUT(n11994), .S0(n5341[16]), .S1(n5341[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1079_18.INIT0 = 16'h5666;
    defparam add_1079_18.INIT1 = 16'h5666;
    defparam add_1079_18.INJECT1_0 = "NO";
    defparam add_1079_18.INJECT1_1 = "NO";
    CCU2D add_1084_32 (.A0(d3[66]), .B0(d4[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[67]), .B1(d4[67]), .C1(GND_net), .D1(GND_net), .CIN(n11959), 
          .COUT(n11960), .S0(n5493[30]), .S1(n5493[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1084_32.INIT0 = 16'h5666;
    defparam add_1084_32.INIT1 = 16'h5666;
    defparam add_1084_32.INJECT1_0 = "NO";
    defparam add_1084_32.INJECT1_1 = "NO";
    CCU2D add_1079_28 (.A0(d2[62]), .B0(d3[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[63]), .B1(d3[63]), .C1(GND_net), .D1(GND_net), .CIN(n11998), 
          .COUT(n11999), .S0(n5341[26]), .S1(n5341[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1079_28.INIT0 = 16'h5666;
    defparam add_1079_28.INIT1 = 16'h5666;
    defparam add_1079_28.INJECT1_0 = "NO";
    defparam add_1079_28.INJECT1_1 = "NO";
    CCU2D add_1075_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5188), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n12007));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1075_1.INIT0 = 16'hF000;
    defparam add_1075_1.INIT1 = 16'h0555;
    defparam add_1075_1.INJECT1_0 = "NO";
    defparam add_1075_1.INJECT1_1 = "NO";
    CCU2D add_1070_5 (.A0(d1[38]), .B0(n5036), .C0(n5037[2]), .D0(MixerOutCos[11]), 
          .A1(d1[39]), .B1(n5036), .C1(n5037[3]), .D1(MixerOutCos[11]), 
          .CIN(n12049), .COUT(n12050), .S0(d1_71__N_418[38]), .S1(d1_71__N_418[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1070_5.INIT0 = 16'h74b8;
    defparam add_1070_5.INIT1 = 16'h74b8;
    defparam add_1070_5.INJECT1_0 = "NO";
    defparam add_1070_5.INJECT1_1 = "NO";
    CCU2D add_1070_3 (.A0(d1[36]), .B0(n5036), .C0(n5037[0]), .D0(MixerOutCos[11]), 
          .A1(d1[37]), .B1(n5036), .C1(n5037[1]), .D1(MixerOutCos[11]), 
          .CIN(n12048), .COUT(n12049), .S0(d1_71__N_418[36]), .S1(d1_71__N_418[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1070_3.INIT0 = 16'h74b8;
    defparam add_1070_3.INIT1 = 16'h74b8;
    defparam add_1070_3.INJECT1_0 = "NO";
    defparam add_1070_3.INJECT1_1 = "NO";
    CCU2D add_1075_33 (.A0(d2[66]), .B0(n5188), .C0(n5189[30]), .D0(d1[66]), 
          .A1(d2[67]), .B1(n5188), .C1(n5189[31]), .D1(d1[67]), .CIN(n12022), 
          .COUT(n12023), .S0(d2_71__N_490[66]), .S1(d2_71__N_490[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1075_33.INIT0 = 16'h74b8;
    defparam add_1075_33.INIT1 = 16'h74b8;
    defparam add_1075_33.INJECT1_0 = "NO";
    defparam add_1075_33.INJECT1_1 = "NO";
    CCU2D add_1090_35 (.A0(d5[68]), .B0(n5644), .C0(n5645[32]), .D0(d4[68]), 
          .A1(d5[69]), .B1(n5644), .C1(n5645[33]), .D1(d4[69]), .CIN(n11900), 
          .COUT(n11901), .S0(d5_71__N_706[68]), .S1(d5_71__N_706[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1090_35.INIT0 = 16'h74b8;
    defparam add_1090_35.INIT1 = 16'h74b8;
    defparam add_1090_35.INJECT1_0 = "NO";
    defparam add_1090_35.INJECT1_1 = "NO";
    CCU2D add_1075_29 (.A0(d2[62]), .B0(n5188), .C0(n5189[26]), .D0(d1[62]), 
          .A1(d2[63]), .B1(n5188), .C1(n5189[27]), .D1(d1[63]), .CIN(n12020), 
          .COUT(n12021), .S0(d2_71__N_490[62]), .S1(d2_71__N_490[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1075_29.INIT0 = 16'h74b8;
    defparam add_1075_29.INIT1 = 16'h74b8;
    defparam add_1075_29.INJECT1_0 = "NO";
    defparam add_1075_29.INJECT1_1 = "NO";
    CCU2D add_1070_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5036), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n12048));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1070_1.INIT0 = 16'hF000;
    defparam add_1070_1.INIT1 = 16'h0555;
    defparam add_1070_1.INJECT1_0 = "NO";
    defparam add_1070_1.INJECT1_1 = "NO";
    CCU2D add_1079_26 (.A0(d2[60]), .B0(d3[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[61]), .B1(d3[61]), .C1(GND_net), .D1(GND_net), .CIN(n11997), 
          .COUT(n11998), .S0(n5341[24]), .S1(n5341[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1079_26.INIT0 = 16'h5666;
    defparam add_1079_26.INIT1 = 16'h5666;
    defparam add_1079_26.INJECT1_0 = "NO";
    defparam add_1079_26.INJECT1_1 = "NO";
    LUT4 i5686_4_lut (.A(n13121), .B(n13), .C(n13123), .D(n13103), .Z(count_15__N_1458)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i5686_4_lut.init = 16'h2000;
    CCU2D add_1074_36 (.A0(d1[70]), .B0(d2[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[71]), .B1(d2[71]), .C1(GND_net), .D1(GND_net), .CIN(n12043), 
          .S0(n5189[34]), .S1(n5189[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1074_36.INIT0 = 16'h5666;
    defparam add_1074_36.INIT1 = 16'h5666;
    defparam add_1074_36.INJECT1_0 = "NO";
    defparam add_1074_36.INJECT1_1 = "NO";
    LUT4 i5653_4_lut (.A(count[1]), .B(count[9]), .C(count[8]), .D(count[7]), 
         .Z(n13121)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5653_4_lut.init = 16'h8000;
    CCU2D add_1090_33 (.A0(d5[66]), .B0(n5644), .C0(n5645[30]), .D0(d4[66]), 
          .A1(d5[67]), .B1(n5644), .C1(n5645[31]), .D1(d4[67]), .CIN(n11899), 
          .COUT(n11900), .S0(d5_71__N_706[66]), .S1(d5_71__N_706[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1090_33.INIT0 = 16'h74b8;
    defparam add_1090_33.INIT1 = 16'h74b8;
    defparam add_1090_33.INJECT1_0 = "NO";
    defparam add_1090_33.INJECT1_1 = "NO";
    LUT4 i1_2_lut (.A(n12790), .B(count[3]), .Z(n13)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut.init = 16'hbbbb;
    CCU2D add_1084_30 (.A0(d3[64]), .B0(d4[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[65]), .B1(d4[65]), .C1(GND_net), .D1(GND_net), .CIN(n11958), 
          .COUT(n11959), .S0(n5493[28]), .S1(n5493[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1084_30.INIT0 = 16'h5666;
    defparam add_1084_30.INIT1 = 16'h5666;
    defparam add_1084_30.INJECT1_0 = "NO";
    defparam add_1084_30.INJECT1_1 = "NO";
    CCU2D add_1084_28 (.A0(d3[62]), .B0(d4[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[63]), .B1(d4[63]), .C1(GND_net), .D1(GND_net), .CIN(n11957), 
          .COUT(n11958), .S0(n5493[26]), .S1(n5493[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1084_28.INIT0 = 16'h5666;
    defparam add_1084_28.INIT1 = 16'h5666;
    defparam add_1084_28.INJECT1_0 = "NO";
    defparam add_1084_28.INJECT1_1 = "NO";
    CCU2D add_1084_26 (.A0(d3[60]), .B0(d4[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[61]), .B1(d4[61]), .C1(GND_net), .D1(GND_net), .CIN(n11956), 
          .COUT(n11957), .S0(n5493[24]), .S1(n5493[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1084_26.INIT0 = 16'h5666;
    defparam add_1084_26.INIT1 = 16'h5666;
    defparam add_1084_26.INJECT1_0 = "NO";
    defparam add_1084_26.INJECT1_1 = "NO";
    CCU2D add_1084_24 (.A0(d3[58]), .B0(d4[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[59]), .B1(d4[59]), .C1(GND_net), .D1(GND_net), .CIN(n11955), 
          .COUT(n11956), .S0(n5493[22]), .S1(n5493[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1084_24.INIT0 = 16'h5666;
    defparam add_1084_24.INIT1 = 16'h5666;
    defparam add_1084_24.INJECT1_0 = "NO";
    defparam add_1084_24.INJECT1_1 = "NO";
    LUT4 i5655_4_lut (.A(count[4]), .B(count[6]), .C(count[2]), .D(count[0]), 
         .Z(n13123)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5655_4_lut.init = 16'h8000;
    CCU2D add_1084_22 (.A0(d3[56]), .B0(d4[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[57]), .B1(d4[57]), .C1(GND_net), .D1(GND_net), .CIN(n11954), 
          .COUT(n11955), .S0(n5493[20]), .S1(n5493[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1084_22.INIT0 = 16'h5666;
    defparam add_1084_22.INIT1 = 16'h5666;
    defparam add_1084_22.INJECT1_0 = "NO";
    defparam add_1084_22.INJECT1_1 = "NO";
    LUT4 i5635_2_lut (.A(count[10]), .B(count[5]), .Z(n13103)) /* synthesis lut_function=(A (B)) */ ;
    defparam i5635_2_lut.init = 16'h8888;
    CCU2D add_1084_20 (.A0(d3[54]), .B0(d4[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[55]), .B1(d4[55]), .C1(GND_net), .D1(GND_net), .CIN(n11953), 
          .COUT(n11954), .S0(n5493[18]), .S1(n5493[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1084_20.INIT0 = 16'h5666;
    defparam add_1084_20.INIT1 = 16'h5666;
    defparam add_1084_20.INJECT1_0 = "NO";
    defparam add_1084_20.INJECT1_1 = "NO";
    CCU2D add_1084_18 (.A0(d3[52]), .B0(d4[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[53]), .B1(d4[53]), .C1(GND_net), .D1(GND_net), .CIN(n11952), 
          .COUT(n11953), .S0(n5493[16]), .S1(n5493[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1084_18.INIT0 = 16'h5666;
    defparam add_1084_18.INIT1 = 16'h5666;
    defparam add_1084_18.INJECT1_0 = "NO";
    defparam add_1084_18.INJECT1_1 = "NO";
    CCU2D add_1084_16 (.A0(d3[50]), .B0(d4[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[51]), .B1(d4[51]), .C1(GND_net), .D1(GND_net), .CIN(n11951), 
          .COUT(n11952), .S0(n5493[14]), .S1(n5493[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1084_16.INIT0 = 16'h5666;
    defparam add_1084_16.INIT1 = 16'h5666;
    defparam add_1084_16.INJECT1_0 = "NO";
    defparam add_1084_16.INJECT1_1 = "NO";
    CCU2D add_1104_11 (.A0(d_tmp[45]), .B0(d_d_tmp[45]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[46]), .B1(d_d_tmp[46]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11610), .COUT(n11611), .S0(n6101[9]), 
          .S1(n6101[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1104_11.INIT0 = 16'h5999;
    defparam add_1104_11.INIT1 = 16'h5999;
    defparam add_1104_11.INJECT1_0 = "NO";
    defparam add_1104_11.INJECT1_1 = "NO";
    CCU2D add_1084_14 (.A0(d3[48]), .B0(d4[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[49]), .B1(d4[49]), .C1(GND_net), .D1(GND_net), .CIN(n11950), 
          .COUT(n11951), .S0(n5493[12]), .S1(n5493[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1084_14.INIT0 = 16'h5666;
    defparam add_1084_14.INIT1 = 16'h5666;
    defparam add_1084_14.INJECT1_0 = "NO";
    defparam add_1084_14.INJECT1_1 = "NO";
    CCU2D add_1084_12 (.A0(d3[46]), .B0(d4[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[47]), .B1(d4[47]), .C1(GND_net), .D1(GND_net), .CIN(n11949), 
          .COUT(n11950), .S0(n5493[10]), .S1(n5493[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1084_12.INIT0 = 16'h5666;
    defparam add_1084_12.INIT1 = 16'h5666;
    defparam add_1084_12.INJECT1_0 = "NO";
    defparam add_1084_12.INJECT1_1 = "NO";
    CCU2D add_1084_10 (.A0(d3[44]), .B0(d4[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[45]), .B1(d4[45]), .C1(GND_net), .D1(GND_net), .CIN(n11948), 
          .COUT(n11949), .S0(n5493[8]), .S1(n5493[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1084_10.INIT0 = 16'h5666;
    defparam add_1084_10.INIT1 = 16'h5666;
    defparam add_1084_10.INJECT1_0 = "NO";
    defparam add_1084_10.INJECT1_1 = "NO";
    CCU2D add_1084_8 (.A0(d3[42]), .B0(d4[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[43]), .B1(d4[43]), .C1(GND_net), .D1(GND_net), .CIN(n11947), 
          .COUT(n11948), .S0(n5493[6]), .S1(n5493[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1084_8.INIT0 = 16'h5666;
    defparam add_1084_8.INIT1 = 16'h5666;
    defparam add_1084_8.INJECT1_0 = "NO";
    defparam add_1084_8.INJECT1_1 = "NO";
    CCU2D add_1084_6 (.A0(d3[40]), .B0(d4[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[41]), .B1(d4[41]), .C1(GND_net), .D1(GND_net), .CIN(n11946), 
          .COUT(n11947), .S0(n5493[4]), .S1(n5493[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1084_6.INIT0 = 16'h5666;
    defparam add_1084_6.INIT1 = 16'h5666;
    defparam add_1084_6.INJECT1_0 = "NO";
    defparam add_1084_6.INJECT1_1 = "NO";
    CCU2D add_1084_4 (.A0(d3[38]), .B0(d4[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[39]), .B1(d4[39]), .C1(GND_net), .D1(GND_net), .CIN(n11945), 
          .COUT(n11946), .S0(n5493[2]), .S1(n5493[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1084_4.INIT0 = 16'h5666;
    defparam add_1084_4.INIT1 = 16'h5666;
    defparam add_1084_4.INJECT1_0 = "NO";
    defparam add_1084_4.INJECT1_1 = "NO";
    CCU2D add_1084_2 (.A0(d3[36]), .B0(d4[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[37]), .B1(d4[37]), .C1(GND_net), .D1(GND_net), .COUT(n11945), 
          .S1(n5493[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1084_2.INIT0 = 16'h7000;
    defparam add_1084_2.INIT1 = 16'h5666;
    defparam add_1084_2.INJECT1_0 = "NO";
    defparam add_1084_2.INJECT1_1 = "NO";
    CCU2D add_1085_37 (.A0(d4[70]), .B0(n5492), .C0(n5493[34]), .D0(d3[70]), 
          .A1(d4[71]), .B1(n5492), .C1(n5493[35]), .D1(d3[71]), .CIN(n11942), 
          .S0(d4_71__N_634[70]), .S1(d4_71__N_634[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1085_37.INIT0 = 16'h74b8;
    defparam add_1085_37.INIT1 = 16'h74b8;
    defparam add_1085_37.INJECT1_0 = "NO";
    defparam add_1085_37.INJECT1_1 = "NO";
    CCU2D add_1085_35 (.A0(d4[68]), .B0(n5492), .C0(n5493[32]), .D0(d3[68]), 
          .A1(d4[69]), .B1(n5492), .C1(n5493[33]), .D1(d3[69]), .CIN(n11941), 
          .COUT(n11942), .S0(d4_71__N_634[68]), .S1(d4_71__N_634[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1085_35.INIT0 = 16'h74b8;
    defparam add_1085_35.INIT1 = 16'h74b8;
    defparam add_1085_35.INJECT1_0 = "NO";
    defparam add_1085_35.INJECT1_1 = "NO";
    CCU2D add_1085_33 (.A0(d4[66]), .B0(n5492), .C0(n5493[30]), .D0(d3[66]), 
          .A1(d4[67]), .B1(n5492), .C1(n5493[31]), .D1(d3[67]), .CIN(n11940), 
          .COUT(n11941), .S0(d4_71__N_634[66]), .S1(d4_71__N_634[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1085_33.INIT0 = 16'h74b8;
    defparam add_1085_33.INIT1 = 16'h74b8;
    defparam add_1085_33.INJECT1_0 = "NO";
    defparam add_1085_33.INJECT1_1 = "NO";
    LUT4 i4_4_lut (.A(n7), .B(count[15]), .C(count[11]), .D(count[14]), 
         .Z(n12790)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i4_4_lut.init = 16'hffef;
    CCU2D add_1085_31 (.A0(d4[64]), .B0(n5492), .C0(n5493[28]), .D0(d3[64]), 
          .A1(d4[65]), .B1(n5492), .C1(n5493[29]), .D1(d3[65]), .CIN(n11939), 
          .COUT(n11940), .S0(d4_71__N_634[64]), .S1(d4_71__N_634[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1085_31.INIT0 = 16'h74b8;
    defparam add_1085_31.INIT1 = 16'h74b8;
    defparam add_1085_31.INJECT1_0 = "NO";
    defparam add_1085_31.INJECT1_1 = "NO";
    LUT4 i2_2_lut (.A(count[13]), .B(count[12]), .Z(n7)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    CCU2D add_1085_29 (.A0(d4[62]), .B0(n5492), .C0(n5493[26]), .D0(d3[62]), 
          .A1(d4[63]), .B1(n5492), .C1(n5493[27]), .D1(d3[63]), .CIN(n11938), 
          .COUT(n11939), .S0(d4_71__N_634[62]), .S1(d4_71__N_634[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1085_29.INIT0 = 16'h74b8;
    defparam add_1085_29.INIT1 = 16'h74b8;
    defparam add_1085_29.INJECT1_0 = "NO";
    defparam add_1085_29.INJECT1_1 = "NO";
    CCU2D add_1085_27 (.A0(d4[60]), .B0(n5492), .C0(n5493[24]), .D0(d3[60]), 
          .A1(d4[61]), .B1(n5492), .C1(n5493[25]), .D1(d3[61]), .CIN(n11937), 
          .COUT(n11938), .S0(d4_71__N_634[60]), .S1(d4_71__N_634[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1085_27.INIT0 = 16'h74b8;
    defparam add_1085_27.INIT1 = 16'h74b8;
    defparam add_1085_27.INJECT1_0 = "NO";
    defparam add_1085_27.INJECT1_1 = "NO";
    CCU2D add_1085_25 (.A0(d4[58]), .B0(n5492), .C0(n5493[22]), .D0(d3[58]), 
          .A1(d4[59]), .B1(n5492), .C1(n5493[23]), .D1(d3[59]), .CIN(n11936), 
          .COUT(n11937), .S0(d4_71__N_634[58]), .S1(d4_71__N_634[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1085_25.INIT0 = 16'h74b8;
    defparam add_1085_25.INIT1 = 16'h74b8;
    defparam add_1085_25.INJECT1_0 = "NO";
    defparam add_1085_25.INJECT1_1 = "NO";
    LUT4 i5686_4_lut_rep_97 (.A(n13121), .B(n13), .C(n13123), .D(n13103), 
         .Z(n13507)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i5686_4_lut_rep_97.init = 16'h2000;
    CCU2D add_1085_23 (.A0(d4[56]), .B0(n5492), .C0(n5493[20]), .D0(d3[56]), 
          .A1(d4[57]), .B1(n5492), .C1(n5493[21]), .D1(d3[57]), .CIN(n11935), 
          .COUT(n11936), .S0(d4_71__N_634[56]), .S1(d4_71__N_634[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1085_23.INIT0 = 16'h74b8;
    defparam add_1085_23.INIT1 = 16'h74b8;
    defparam add_1085_23.INJECT1_0 = "NO";
    defparam add_1085_23.INJECT1_1 = "NO";
    CCU2D add_1085_21 (.A0(d4[54]), .B0(n5492), .C0(n5493[18]), .D0(d3[54]), 
          .A1(d4[55]), .B1(n5492), .C1(n5493[19]), .D1(d3[55]), .CIN(n11934), 
          .COUT(n11935), .S0(d4_71__N_634[54]), .S1(d4_71__N_634[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1085_21.INIT0 = 16'h74b8;
    defparam add_1085_21.INIT1 = 16'h74b8;
    defparam add_1085_21.INJECT1_0 = "NO";
    defparam add_1085_21.INJECT1_1 = "NO";
    CCU2D add_1085_19 (.A0(d4[52]), .B0(n5492), .C0(n5493[16]), .D0(d3[52]), 
          .A1(d4[53]), .B1(n5492), .C1(n5493[17]), .D1(d3[53]), .CIN(n11933), 
          .COUT(n11934), .S0(d4_71__N_634[52]), .S1(d4_71__N_634[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1085_19.INIT0 = 16'h74b8;
    defparam add_1085_19.INIT1 = 16'h74b8;
    defparam add_1085_19.INJECT1_0 = "NO";
    defparam add_1085_19.INJECT1_1 = "NO";
    LUT4 i3_2_lut (.A(count[8]), .B(count[7]), .Z(n15)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i3_2_lut.init = 16'heeee;
    CCU2D add_1085_17 (.A0(d4[50]), .B0(n5492), .C0(n5493[14]), .D0(d3[50]), 
          .A1(d4[51]), .B1(n5492), .C1(n5493[15]), .D1(d3[51]), .CIN(n11932), 
          .COUT(n11933), .S0(d4_71__N_634[50]), .S1(d4_71__N_634[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1085_17.INIT0 = 16'h74b8;
    defparam add_1085_17.INIT1 = 16'h74b8;
    defparam add_1085_17.INJECT1_0 = "NO";
    defparam add_1085_17.INJECT1_1 = "NO";
    CCU2D add_1085_15 (.A0(d4[48]), .B0(n5492), .C0(n5493[12]), .D0(d3[48]), 
          .A1(d4[49]), .B1(n5492), .C1(n5493[13]), .D1(d3[49]), .CIN(n11931), 
          .COUT(n11932), .S0(d4_71__N_634[48]), .S1(d4_71__N_634[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1085_15.INIT0 = 16'h74b8;
    defparam add_1085_15.INIT1 = 16'h74b8;
    defparam add_1085_15.INJECT1_0 = "NO";
    defparam add_1085_15.INJECT1_1 = "NO";
    CCU2D add_1085_13 (.A0(d4[46]), .B0(n5492), .C0(n5493[10]), .D0(d3[46]), 
          .A1(d4[47]), .B1(n5492), .C1(n5493[11]), .D1(d3[47]), .CIN(n11930), 
          .COUT(n11931), .S0(d4_71__N_634[46]), .S1(d4_71__N_634[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1085_13.INIT0 = 16'h74b8;
    defparam add_1085_13.INIT1 = 16'h74b8;
    defparam add_1085_13.INJECT1_0 = "NO";
    defparam add_1085_13.INJECT1_1 = "NO";
    LUT4 i4_2_lut (.A(n12790), .B(count[2]), .Z(n16)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i4_2_lut.init = 16'heeee;
    CCU2D add_1085_11 (.A0(d4[44]), .B0(n5492), .C0(n5493[8]), .D0(d3[44]), 
          .A1(d4[45]), .B1(n5492), .C1(n5493[9]), .D1(d3[45]), .CIN(n11929), 
          .COUT(n11930), .S0(d4_71__N_634[44]), .S1(d4_71__N_634[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1085_11.INIT0 = 16'h74b8;
    defparam add_1085_11.INIT1 = 16'h74b8;
    defparam add_1085_11.INJECT1_0 = "NO";
    defparam add_1085_11.INJECT1_1 = "NO";
    CCU2D add_1085_9 (.A0(d4[42]), .B0(n5492), .C0(n5493[6]), .D0(d3[42]), 
          .A1(d4[43]), .B1(n5492), .C1(n5493[7]), .D1(d3[43]), .CIN(n11928), 
          .COUT(n11929), .S0(d4_71__N_634[42]), .S1(d4_71__N_634[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1085_9.INIT0 = 16'h74b8;
    defparam add_1085_9.INIT1 = 16'h74b8;
    defparam add_1085_9.INJECT1_0 = "NO";
    defparam add_1085_9.INJECT1_1 = "NO";
    CCU2D add_1085_7 (.A0(d4[40]), .B0(n5492), .C0(n5493[4]), .D0(d3[40]), 
          .A1(d4[41]), .B1(n5492), .C1(n5493[5]), .D1(d3[41]), .CIN(n11927), 
          .COUT(n11928), .S0(d4_71__N_634[40]), .S1(d4_71__N_634[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1085_7.INIT0 = 16'h74b8;
    defparam add_1085_7.INIT1 = 16'h74b8;
    defparam add_1085_7.INJECT1_0 = "NO";
    defparam add_1085_7.INJECT1_1 = "NO";
    CCU2D add_1085_5 (.A0(d4[38]), .B0(n5492), .C0(n5493[2]), .D0(d3[38]), 
          .A1(d4[39]), .B1(n5492), .C1(n5493[3]), .D1(d3[39]), .CIN(n11926), 
          .COUT(n11927), .S0(d4_71__N_634[38]), .S1(d4_71__N_634[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1085_5.INIT0 = 16'h74b8;
    defparam add_1085_5.INIT1 = 16'h74b8;
    defparam add_1085_5.INJECT1_0 = "NO";
    defparam add_1085_5.INJECT1_1 = "NO";
    CCU2D add_1085_3 (.A0(d4[36]), .B0(n5492), .C0(n5493[0]), .D0(d3[36]), 
          .A1(d4[37]), .B1(n5492), .C1(n5493[1]), .D1(d3[37]), .CIN(n11925), 
          .COUT(n11926), .S0(d4_71__N_634[36]), .S1(d4_71__N_634[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1085_3.INIT0 = 16'h74b8;
    defparam add_1085_3.INIT1 = 16'h74b8;
    defparam add_1085_3.INJECT1_0 = "NO";
    defparam add_1085_3.INJECT1_1 = "NO";
    CCU2D add_1085_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5492), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11925));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1085_1.INIT0 = 16'hF000;
    defparam add_1085_1.INIT1 = 16'h0555;
    defparam add_1085_1.INJECT1_0 = "NO";
    defparam add_1085_1.INJECT1_1 = "NO";
    CCU2D add_1089_36 (.A0(d4[70]), .B0(d5[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[71]), .B1(d5[71]), .C1(GND_net), .D1(GND_net), .CIN(n11920), 
          .S0(n5645[34]), .S1(n5645[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1089_36.INIT0 = 16'h5666;
    defparam add_1089_36.INIT1 = 16'h5666;
    defparam add_1089_36.INJECT1_0 = "NO";
    defparam add_1089_36.INJECT1_1 = "NO";
    CCU2D add_1089_34 (.A0(d4[68]), .B0(d5[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[69]), .B1(d5[69]), .C1(GND_net), .D1(GND_net), .CIN(n11919), 
          .COUT(n11920), .S0(n5645[32]), .S1(n5645[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1089_34.INIT0 = 16'h5666;
    defparam add_1089_34.INIT1 = 16'h5666;
    defparam add_1089_34.INJECT1_0 = "NO";
    defparam add_1089_34.INJECT1_1 = "NO";
    CCU2D add_1089_32 (.A0(d4[66]), .B0(d5[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[67]), .B1(d5[67]), .C1(GND_net), .D1(GND_net), .CIN(n11918), 
          .COUT(n11919), .S0(n5645[30]), .S1(n5645[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1089_32.INIT0 = 16'h5666;
    defparam add_1089_32.INIT1 = 16'h5666;
    defparam add_1089_32.INJECT1_0 = "NO";
    defparam add_1089_32.INJECT1_1 = "NO";
    CCU2D add_1089_30 (.A0(d4[64]), .B0(d5[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[65]), .B1(d5[65]), .C1(GND_net), .D1(GND_net), .CIN(n11917), 
          .COUT(n11918), .S0(n5645[28]), .S1(n5645[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1089_30.INIT0 = 16'h5666;
    defparam add_1089_30.INIT1 = 16'h5666;
    defparam add_1089_30.INJECT1_0 = "NO";
    defparam add_1089_30.INJECT1_1 = "NO";
    LUT4 i4948_2_lut (.A(d2[36]), .B(d3[36]), .Z(n5341[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4948_2_lut.init = 16'h6666;
    CCU2D add_1089_28 (.A0(d4[62]), .B0(d5[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[63]), .B1(d5[63]), .C1(GND_net), .D1(GND_net), .CIN(n11916), 
          .COUT(n11917), .S0(n5645[26]), .S1(n5645[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1089_28.INIT0 = 16'h5666;
    defparam add_1089_28.INIT1 = 16'h5666;
    defparam add_1089_28.INJECT1_0 = "NO";
    defparam add_1089_28.INJECT1_1 = "NO";
    CCU2D add_1089_26 (.A0(d4[60]), .B0(d5[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[61]), .B1(d5[61]), .C1(GND_net), .D1(GND_net), .CIN(n11915), 
          .COUT(n11916), .S0(n5645[24]), .S1(n5645[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1089_26.INIT0 = 16'h5666;
    defparam add_1089_26.INIT1 = 16'h5666;
    defparam add_1089_26.INJECT1_0 = "NO";
    defparam add_1089_26.INJECT1_1 = "NO";
    CCU2D add_1089_24 (.A0(d4[58]), .B0(d5[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[59]), .B1(d5[59]), .C1(GND_net), .D1(GND_net), .CIN(n11914), 
          .COUT(n11915), .S0(n5645[22]), .S1(n5645[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1089_24.INIT0 = 16'h5666;
    defparam add_1089_24.INIT1 = 16'h5666;
    defparam add_1089_24.INJECT1_0 = "NO";
    defparam add_1089_24.INJECT1_1 = "NO";
    CCU2D add_1089_22 (.A0(d4[56]), .B0(d5[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[57]), .B1(d5[57]), .C1(GND_net), .D1(GND_net), .CIN(n11913), 
          .COUT(n11914), .S0(n5645[20]), .S1(n5645[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1089_22.INIT0 = 16'h5666;
    defparam add_1089_22.INIT1 = 16'h5666;
    defparam add_1089_22.INJECT1_0 = "NO";
    defparam add_1089_22.INJECT1_1 = "NO";
    CCU2D add_1089_20 (.A0(d4[54]), .B0(d5[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[55]), .B1(d5[55]), .C1(GND_net), .D1(GND_net), .CIN(n11912), 
          .COUT(n11913), .S0(n5645[18]), .S1(n5645[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1089_20.INIT0 = 16'h5666;
    defparam add_1089_20.INIT1 = 16'h5666;
    defparam add_1089_20.INJECT1_0 = "NO";
    defparam add_1089_20.INJECT1_1 = "NO";
    FD1P3AX d_tmp_i0_i1 (.D(d5[1]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i2 (.D(d5[2]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i3 (.D(d5[3]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i4 (.D(d5[4]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i5 (.D(d5[5]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i6 (.D(d5[6]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i7 (.D(d5[7]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i8 (.D(d5[8]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i9 (.D(d5[9]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i10 (.D(d5[10]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i11 (.D(d5[11]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i12 (.D(d5[12]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i13 (.D(d5[13]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i14 (.D(d5[14]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i15 (.D(d5[15]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i16 (.D(d5[16]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i17 (.D(d5[17]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i18 (.D(d5[18]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i19 (.D(d5[19]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i20 (.D(d5[20]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i21 (.D(d5[21]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i22 (.D(d5[22]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i23 (.D(d5[23]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i24 (.D(d5[24]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i25 (.D(d5[25]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i26 (.D(d5[26]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i27 (.D(d5[27]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i28 (.D(d5[28]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i29 (.D(d5[29]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i30 (.D(d5[30]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i31 (.D(d5[31]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i32 (.D(d5[32]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i33 (.D(d5[33]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i34 (.D(d5[34]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i35 (.D(d5[35]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i36 (.D(d5[36]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i37 (.D(d5[37]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i38 (.D(d5[38]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i39 (.D(d5[39]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i40 (.D(d5[40]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i41 (.D(d5[41]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i42 (.D(d5[42]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i43 (.D(d5[43]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i44 (.D(d5[44]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i45 (.D(d5[45]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i46 (.D(d5[46]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i47 (.D(d5[47]), .SP(osc_clk_enable_744), .CK(osc_clk), 
            .Q(d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i48 (.D(d5[48]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i49 (.D(d5[49]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i50 (.D(d5[50]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i51 (.D(d5[51]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i52 (.D(d5[52]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i53 (.D(d5[53]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i54 (.D(d5[54]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i55 (.D(d5[55]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i56 (.D(d5[56]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i57 (.D(d5[57]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i58 (.D(d5[58]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i59 (.D(d5[59]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i60 (.D(d5[60]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i61 (.D(d5[61]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i62 (.D(d5[62]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i63 (.D(d5[63]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i64 (.D(d5[64]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i65 (.D(d5[65]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i66 (.D(d5[66]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i67 (.D(d5[67]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i68 (.D(d5[68]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i69 (.D(d5[69]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i70 (.D(d5[70]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i71 (.D(d5[71]), .SP(count_15__N_1458), .CK(osc_clk), 
            .Q(d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i1 (.D(d_tmp[1]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i2 (.D(d_tmp[2]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i3 (.D(d_tmp[3]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i4 (.D(d_tmp[4]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i5 (.D(d_tmp[5]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i6 (.D(d_tmp[6]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i7 (.D(d_tmp[7]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i8 (.D(d_tmp[8]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i9 (.D(d_tmp[9]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i10 (.D(d_tmp[10]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i11 (.D(d_tmp[11]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i12 (.D(d_tmp[12]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i13 (.D(d_tmp[13]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i14 (.D(d_tmp[14]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i15 (.D(d_tmp[15]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i16 (.D(d_tmp[16]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i17 (.D(d_tmp[17]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i18 (.D(d_tmp[18]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i19 (.D(d_tmp[19]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i20 (.D(d_tmp[20]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i21 (.D(d_tmp[21]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i22 (.D(d_tmp[22]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i23 (.D(d_tmp[23]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i24 (.D(d_tmp[24]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i25 (.D(d_tmp[25]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i26 (.D(d_tmp[26]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i27 (.D(d_tmp[27]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i28 (.D(d_tmp[28]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i29 (.D(d_tmp[29]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i30 (.D(d_tmp[30]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i31 (.D(d_tmp[31]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i32 (.D(d_tmp[32]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i33 (.D(d_tmp[33]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i34 (.D(d_tmp[34]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i35 (.D(d_tmp[35]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i36 (.D(d_tmp[36]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i37 (.D(d_tmp[37]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i38 (.D(d_tmp[38]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i39 (.D(d_tmp[39]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i40 (.D(d_tmp[40]), .SP(osc_clk_enable_784), .CK(osc_clk), 
            .Q(d_d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i41 (.D(d_tmp[41]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i42 (.D(d_tmp[42]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i43 (.D(d_tmp[43]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i44 (.D(d_tmp[44]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i45 (.D(d_tmp[45]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i46 (.D(d_tmp[46]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i47 (.D(d_tmp[47]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i48 (.D(d_tmp[48]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i49 (.D(d_tmp[49]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i50 (.D(d_tmp[50]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i51 (.D(d_tmp[51]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i52 (.D(d_tmp[52]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i53 (.D(d_tmp[53]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i54 (.D(d_tmp[54]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i55 (.D(d_tmp[55]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i56 (.D(d_tmp[56]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i57 (.D(d_tmp[57]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i58 (.D(d_tmp[58]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i59 (.D(d_tmp[59]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i60 (.D(d_tmp[60]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i61 (.D(d_tmp[61]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i62 (.D(d_tmp[62]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i63 (.D(d_tmp[63]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i64 (.D(d_tmp[64]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i65 (.D(d_tmp[65]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i66 (.D(d_tmp[66]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i67 (.D(d_tmp[67]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i68 (.D(d_tmp[68]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i69 (.D(d_tmp[69]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i70 (.D(d_tmp[70]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i71 (.D(d_tmp[71]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d_d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i71.GSR = "ENABLED";
    FD1S3AX d2_i1 (.D(d2_71__N_490[1]), .CK(osc_clk), .Q(d2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i1.GSR = "ENABLED";
    FD1S3AX d2_i2 (.D(d2_71__N_490[2]), .CK(osc_clk), .Q(d2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i2.GSR = "ENABLED";
    FD1S3AX d2_i3 (.D(d2_71__N_490[3]), .CK(osc_clk), .Q(d2[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i3.GSR = "ENABLED";
    FD1S3AX d2_i4 (.D(d2_71__N_490[4]), .CK(osc_clk), .Q(d2[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i4.GSR = "ENABLED";
    FD1S3AX d2_i5 (.D(d2_71__N_490[5]), .CK(osc_clk), .Q(d2[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i5.GSR = "ENABLED";
    FD1S3AX d2_i6 (.D(d2_71__N_490[6]), .CK(osc_clk), .Q(d2[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i6.GSR = "ENABLED";
    FD1S3AX d2_i7 (.D(d2_71__N_490[7]), .CK(osc_clk), .Q(d2[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i7.GSR = "ENABLED";
    FD1S3AX d2_i8 (.D(d2_71__N_490[8]), .CK(osc_clk), .Q(d2[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i8.GSR = "ENABLED";
    FD1S3AX d2_i9 (.D(d2_71__N_490[9]), .CK(osc_clk), .Q(d2[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i9.GSR = "ENABLED";
    FD1S3AX d2_i10 (.D(d2_71__N_490[10]), .CK(osc_clk), .Q(d2[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i10.GSR = "ENABLED";
    FD1S3AX d2_i11 (.D(d2_71__N_490[11]), .CK(osc_clk), .Q(d2[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i11.GSR = "ENABLED";
    FD1S3AX d2_i12 (.D(d2_71__N_490[12]), .CK(osc_clk), .Q(d2[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i12.GSR = "ENABLED";
    FD1S3AX d2_i13 (.D(d2_71__N_490[13]), .CK(osc_clk), .Q(d2[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i13.GSR = "ENABLED";
    FD1S3AX d2_i14 (.D(d2_71__N_490[14]), .CK(osc_clk), .Q(d2[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i14.GSR = "ENABLED";
    FD1S3AX d2_i15 (.D(d2_71__N_490[15]), .CK(osc_clk), .Q(d2[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i15.GSR = "ENABLED";
    FD1S3AX d2_i16 (.D(d2_71__N_490[16]), .CK(osc_clk), .Q(d2[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i16.GSR = "ENABLED";
    FD1S3AX d2_i17 (.D(d2_71__N_490[17]), .CK(osc_clk), .Q(d2[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i17.GSR = "ENABLED";
    FD1S3AX d2_i18 (.D(d2_71__N_490[18]), .CK(osc_clk), .Q(d2[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i18.GSR = "ENABLED";
    FD1S3AX d2_i19 (.D(d2_71__N_490[19]), .CK(osc_clk), .Q(d2[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i19.GSR = "ENABLED";
    FD1S3AX d2_i20 (.D(d2_71__N_490[20]), .CK(osc_clk), .Q(d2[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i20.GSR = "ENABLED";
    FD1S3AX d2_i21 (.D(d2_71__N_490[21]), .CK(osc_clk), .Q(d2[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i21.GSR = "ENABLED";
    FD1S3AX d2_i22 (.D(d2_71__N_490[22]), .CK(osc_clk), .Q(d2[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i22.GSR = "ENABLED";
    FD1S3AX d2_i23 (.D(d2_71__N_490[23]), .CK(osc_clk), .Q(d2[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i23.GSR = "ENABLED";
    FD1S3AX d2_i24 (.D(d2_71__N_490[24]), .CK(osc_clk), .Q(d2[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i24.GSR = "ENABLED";
    FD1S3AX d2_i25 (.D(d2_71__N_490[25]), .CK(osc_clk), .Q(d2[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i25.GSR = "ENABLED";
    FD1S3AX d2_i26 (.D(d2_71__N_490[26]), .CK(osc_clk), .Q(d2[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i26.GSR = "ENABLED";
    FD1S3AX d2_i27 (.D(d2_71__N_490[27]), .CK(osc_clk), .Q(d2[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i27.GSR = "ENABLED";
    FD1S3AX d2_i28 (.D(d2_71__N_490[28]), .CK(osc_clk), .Q(d2[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i28.GSR = "ENABLED";
    FD1S3AX d2_i29 (.D(d2_71__N_490[29]), .CK(osc_clk), .Q(d2[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i29.GSR = "ENABLED";
    FD1S3AX d2_i30 (.D(d2_71__N_490[30]), .CK(osc_clk), .Q(d2[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i30.GSR = "ENABLED";
    FD1S3AX d2_i31 (.D(d2_71__N_490[31]), .CK(osc_clk), .Q(d2[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i31.GSR = "ENABLED";
    FD1S3AX d2_i32 (.D(d2_71__N_490[32]), .CK(osc_clk), .Q(d2[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i32.GSR = "ENABLED";
    FD1S3AX d2_i33 (.D(d2_71__N_490[33]), .CK(osc_clk), .Q(d2[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i33.GSR = "ENABLED";
    FD1S3AX d2_i34 (.D(d2_71__N_490[34]), .CK(osc_clk), .Q(d2[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i34.GSR = "ENABLED";
    FD1S3AX d2_i35 (.D(d2_71__N_490[35]), .CK(osc_clk), .Q(d2[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i35.GSR = "ENABLED";
    FD1S3AX d2_i36 (.D(d2_71__N_490[36]), .CK(osc_clk), .Q(d2[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i36.GSR = "ENABLED";
    FD1S3AX d2_i37 (.D(d2_71__N_490[37]), .CK(osc_clk), .Q(d2[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i37.GSR = "ENABLED";
    FD1S3AX d2_i38 (.D(d2_71__N_490[38]), .CK(osc_clk), .Q(d2[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i38.GSR = "ENABLED";
    FD1S3AX d2_i39 (.D(d2_71__N_490[39]), .CK(osc_clk), .Q(d2[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i39.GSR = "ENABLED";
    FD1S3AX d2_i40 (.D(d2_71__N_490[40]), .CK(osc_clk), .Q(d2[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i40.GSR = "ENABLED";
    FD1S3AX d2_i41 (.D(d2_71__N_490[41]), .CK(osc_clk), .Q(d2[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i41.GSR = "ENABLED";
    FD1S3AX d2_i42 (.D(d2_71__N_490[42]), .CK(osc_clk), .Q(d2[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i42.GSR = "ENABLED";
    FD1S3AX d2_i43 (.D(d2_71__N_490[43]), .CK(osc_clk), .Q(d2[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i43.GSR = "ENABLED";
    FD1S3AX d2_i44 (.D(d2_71__N_490[44]), .CK(osc_clk), .Q(d2[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i44.GSR = "ENABLED";
    FD1S3AX d2_i45 (.D(d2_71__N_490[45]), .CK(osc_clk), .Q(d2[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i45.GSR = "ENABLED";
    FD1S3AX d2_i46 (.D(d2_71__N_490[46]), .CK(osc_clk), .Q(d2[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i46.GSR = "ENABLED";
    FD1S3AX d2_i47 (.D(d2_71__N_490[47]), .CK(osc_clk), .Q(d2[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i47.GSR = "ENABLED";
    FD1S3AX d2_i48 (.D(d2_71__N_490[48]), .CK(osc_clk), .Q(d2[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i48.GSR = "ENABLED";
    FD1S3AX d2_i49 (.D(d2_71__N_490[49]), .CK(osc_clk), .Q(d2[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i49.GSR = "ENABLED";
    FD1S3AX d2_i50 (.D(d2_71__N_490[50]), .CK(osc_clk), .Q(d2[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i50.GSR = "ENABLED";
    FD1S3AX d2_i51 (.D(d2_71__N_490[51]), .CK(osc_clk), .Q(d2[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i51.GSR = "ENABLED";
    FD1S3AX d2_i52 (.D(d2_71__N_490[52]), .CK(osc_clk), .Q(d2[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i52.GSR = "ENABLED";
    FD1S3AX d2_i53 (.D(d2_71__N_490[53]), .CK(osc_clk), .Q(d2[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i53.GSR = "ENABLED";
    FD1S3AX d2_i54 (.D(d2_71__N_490[54]), .CK(osc_clk), .Q(d2[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i54.GSR = "ENABLED";
    FD1S3AX d2_i55 (.D(d2_71__N_490[55]), .CK(osc_clk), .Q(d2[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i55.GSR = "ENABLED";
    FD1S3AX d2_i56 (.D(d2_71__N_490[56]), .CK(osc_clk), .Q(d2[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i56.GSR = "ENABLED";
    FD1S3AX d2_i57 (.D(d2_71__N_490[57]), .CK(osc_clk), .Q(d2[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i57.GSR = "ENABLED";
    FD1S3AX d2_i58 (.D(d2_71__N_490[58]), .CK(osc_clk), .Q(d2[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i58.GSR = "ENABLED";
    FD1S3AX d2_i59 (.D(d2_71__N_490[59]), .CK(osc_clk), .Q(d2[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i59.GSR = "ENABLED";
    FD1S3AX d2_i60 (.D(d2_71__N_490[60]), .CK(osc_clk), .Q(d2[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i60.GSR = "ENABLED";
    FD1S3AX d2_i61 (.D(d2_71__N_490[61]), .CK(osc_clk), .Q(d2[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i61.GSR = "ENABLED";
    FD1S3AX d2_i62 (.D(d2_71__N_490[62]), .CK(osc_clk), .Q(d2[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i62.GSR = "ENABLED";
    FD1S3AX d2_i63 (.D(d2_71__N_490[63]), .CK(osc_clk), .Q(d2[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i63.GSR = "ENABLED";
    FD1S3AX d2_i64 (.D(d2_71__N_490[64]), .CK(osc_clk), .Q(d2[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i64.GSR = "ENABLED";
    FD1S3AX d2_i65 (.D(d2_71__N_490[65]), .CK(osc_clk), .Q(d2[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i65.GSR = "ENABLED";
    FD1S3AX d2_i66 (.D(d2_71__N_490[66]), .CK(osc_clk), .Q(d2[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i66.GSR = "ENABLED";
    FD1S3AX d2_i67 (.D(d2_71__N_490[67]), .CK(osc_clk), .Q(d2[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i67.GSR = "ENABLED";
    FD1S3AX d2_i68 (.D(d2_71__N_490[68]), .CK(osc_clk), .Q(d2[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i68.GSR = "ENABLED";
    FD1S3AX d2_i69 (.D(d2_71__N_490[69]), .CK(osc_clk), .Q(d2[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i69.GSR = "ENABLED";
    FD1S3AX d2_i70 (.D(d2_71__N_490[70]), .CK(osc_clk), .Q(d2[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i70.GSR = "ENABLED";
    FD1S3AX d2_i71 (.D(d2_71__N_490[71]), .CK(osc_clk), .Q(d2[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i71.GSR = "ENABLED";
    FD1S3AX d3_i1 (.D(d3_71__N_562[1]), .CK(osc_clk), .Q(d3[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i1.GSR = "ENABLED";
    FD1S3AX d3_i2 (.D(d3_71__N_562[2]), .CK(osc_clk), .Q(d3[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i2.GSR = "ENABLED";
    FD1S3AX d3_i3 (.D(d3_71__N_562[3]), .CK(osc_clk), .Q(d3[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i3.GSR = "ENABLED";
    FD1S3AX d3_i4 (.D(d3_71__N_562[4]), .CK(osc_clk), .Q(d3[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i4.GSR = "ENABLED";
    FD1S3AX d3_i5 (.D(d3_71__N_562[5]), .CK(osc_clk), .Q(d3[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i5.GSR = "ENABLED";
    FD1S3AX d3_i6 (.D(d3_71__N_562[6]), .CK(osc_clk), .Q(d3[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i6.GSR = "ENABLED";
    FD1S3AX d3_i7 (.D(d3_71__N_562[7]), .CK(osc_clk), .Q(d3[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i7.GSR = "ENABLED";
    FD1S3AX d3_i8 (.D(d3_71__N_562[8]), .CK(osc_clk), .Q(d3[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i8.GSR = "ENABLED";
    FD1S3AX d3_i9 (.D(d3_71__N_562[9]), .CK(osc_clk), .Q(d3[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i9.GSR = "ENABLED";
    FD1S3AX d3_i10 (.D(d3_71__N_562[10]), .CK(osc_clk), .Q(d3[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i10.GSR = "ENABLED";
    FD1S3AX d3_i11 (.D(d3_71__N_562[11]), .CK(osc_clk), .Q(d3[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i11.GSR = "ENABLED";
    FD1S3AX d3_i12 (.D(d3_71__N_562[12]), .CK(osc_clk), .Q(d3[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i12.GSR = "ENABLED";
    FD1S3AX d3_i13 (.D(d3_71__N_562[13]), .CK(osc_clk), .Q(d3[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i13.GSR = "ENABLED";
    FD1S3AX d3_i14 (.D(d3_71__N_562[14]), .CK(osc_clk), .Q(d3[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i14.GSR = "ENABLED";
    FD1S3AX d3_i15 (.D(d3_71__N_562[15]), .CK(osc_clk), .Q(d3[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i15.GSR = "ENABLED";
    FD1S3AX d3_i16 (.D(d3_71__N_562[16]), .CK(osc_clk), .Q(d3[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i16.GSR = "ENABLED";
    FD1S3AX d3_i17 (.D(d3_71__N_562[17]), .CK(osc_clk), .Q(d3[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i17.GSR = "ENABLED";
    FD1S3AX d3_i18 (.D(d3_71__N_562[18]), .CK(osc_clk), .Q(d3[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i18.GSR = "ENABLED";
    FD1S3AX d3_i19 (.D(d3_71__N_562[19]), .CK(osc_clk), .Q(d3[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i19.GSR = "ENABLED";
    FD1S3AX d3_i20 (.D(d3_71__N_562[20]), .CK(osc_clk), .Q(d3[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i20.GSR = "ENABLED";
    FD1S3AX d3_i21 (.D(d3_71__N_562[21]), .CK(osc_clk), .Q(d3[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i21.GSR = "ENABLED";
    FD1S3AX d3_i22 (.D(d3_71__N_562[22]), .CK(osc_clk), .Q(d3[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i22.GSR = "ENABLED";
    FD1S3AX d3_i23 (.D(d3_71__N_562[23]), .CK(osc_clk), .Q(d3[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i23.GSR = "ENABLED";
    FD1S3AX d3_i24 (.D(d3_71__N_562[24]), .CK(osc_clk), .Q(d3[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i24.GSR = "ENABLED";
    FD1S3AX d3_i25 (.D(d3_71__N_562[25]), .CK(osc_clk), .Q(d3[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i25.GSR = "ENABLED";
    FD1S3AX d3_i26 (.D(d3_71__N_562[26]), .CK(osc_clk), .Q(d3[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i26.GSR = "ENABLED";
    FD1S3AX d3_i27 (.D(d3_71__N_562[27]), .CK(osc_clk), .Q(d3[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i27.GSR = "ENABLED";
    FD1S3AX d3_i28 (.D(d3_71__N_562[28]), .CK(osc_clk), .Q(d3[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i28.GSR = "ENABLED";
    FD1S3AX d3_i29 (.D(d3_71__N_562[29]), .CK(osc_clk), .Q(d3[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i29.GSR = "ENABLED";
    FD1S3AX d3_i30 (.D(d3_71__N_562[30]), .CK(osc_clk), .Q(d3[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i30.GSR = "ENABLED";
    FD1S3AX d3_i31 (.D(d3_71__N_562[31]), .CK(osc_clk), .Q(d3[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i31.GSR = "ENABLED";
    FD1S3AX d3_i32 (.D(d3_71__N_562[32]), .CK(osc_clk), .Q(d3[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i32.GSR = "ENABLED";
    FD1S3AX d3_i33 (.D(d3_71__N_562[33]), .CK(osc_clk), .Q(d3[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i33.GSR = "ENABLED";
    FD1S3AX d3_i34 (.D(d3_71__N_562[34]), .CK(osc_clk), .Q(d3[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i34.GSR = "ENABLED";
    FD1S3AX d3_i35 (.D(d3_71__N_562[35]), .CK(osc_clk), .Q(d3[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i35.GSR = "ENABLED";
    FD1S3AX d3_i36 (.D(d3_71__N_562[36]), .CK(osc_clk), .Q(d3[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i36.GSR = "ENABLED";
    FD1S3AX d3_i37 (.D(d3_71__N_562[37]), .CK(osc_clk), .Q(d3[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i37.GSR = "ENABLED";
    FD1S3AX d3_i38 (.D(d3_71__N_562[38]), .CK(osc_clk), .Q(d3[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i38.GSR = "ENABLED";
    FD1S3AX d3_i39 (.D(d3_71__N_562[39]), .CK(osc_clk), .Q(d3[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i39.GSR = "ENABLED";
    FD1S3AX d3_i40 (.D(d3_71__N_562[40]), .CK(osc_clk), .Q(d3[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i40.GSR = "ENABLED";
    FD1S3AX d3_i41 (.D(d3_71__N_562[41]), .CK(osc_clk), .Q(d3[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i41.GSR = "ENABLED";
    FD1S3AX d3_i42 (.D(d3_71__N_562[42]), .CK(osc_clk), .Q(d3[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i42.GSR = "ENABLED";
    FD1S3AX d3_i43 (.D(d3_71__N_562[43]), .CK(osc_clk), .Q(d3[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i43.GSR = "ENABLED";
    FD1S3AX d3_i44 (.D(d3_71__N_562[44]), .CK(osc_clk), .Q(d3[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i44.GSR = "ENABLED";
    FD1S3AX d3_i45 (.D(d3_71__N_562[45]), .CK(osc_clk), .Q(d3[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i45.GSR = "ENABLED";
    FD1S3AX d3_i46 (.D(d3_71__N_562[46]), .CK(osc_clk), .Q(d3[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i46.GSR = "ENABLED";
    FD1S3AX d3_i47 (.D(d3_71__N_562[47]), .CK(osc_clk), .Q(d3[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i47.GSR = "ENABLED";
    FD1S3AX d3_i48 (.D(d3_71__N_562[48]), .CK(osc_clk), .Q(d3[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i48.GSR = "ENABLED";
    FD1S3AX d3_i49 (.D(d3_71__N_562[49]), .CK(osc_clk), .Q(d3[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i49.GSR = "ENABLED";
    FD1S3AX d3_i50 (.D(d3_71__N_562[50]), .CK(osc_clk), .Q(d3[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i50.GSR = "ENABLED";
    FD1S3AX d3_i51 (.D(d3_71__N_562[51]), .CK(osc_clk), .Q(d3[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i51.GSR = "ENABLED";
    FD1S3AX d3_i52 (.D(d3_71__N_562[52]), .CK(osc_clk), .Q(d3[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i52.GSR = "ENABLED";
    FD1S3AX d3_i53 (.D(d3_71__N_562[53]), .CK(osc_clk), .Q(d3[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i53.GSR = "ENABLED";
    FD1S3AX d3_i54 (.D(d3_71__N_562[54]), .CK(osc_clk), .Q(d3[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i54.GSR = "ENABLED";
    FD1S3AX d3_i55 (.D(d3_71__N_562[55]), .CK(osc_clk), .Q(d3[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i55.GSR = "ENABLED";
    FD1S3AX d3_i56 (.D(d3_71__N_562[56]), .CK(osc_clk), .Q(d3[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i56.GSR = "ENABLED";
    FD1S3AX d3_i57 (.D(d3_71__N_562[57]), .CK(osc_clk), .Q(d3[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i57.GSR = "ENABLED";
    FD1S3AX d3_i58 (.D(d3_71__N_562[58]), .CK(osc_clk), .Q(d3[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i58.GSR = "ENABLED";
    FD1S3AX d3_i59 (.D(d3_71__N_562[59]), .CK(osc_clk), .Q(d3[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i59.GSR = "ENABLED";
    FD1S3AX d3_i60 (.D(d3_71__N_562[60]), .CK(osc_clk), .Q(d3[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i60.GSR = "ENABLED";
    FD1S3AX d3_i61 (.D(d3_71__N_562[61]), .CK(osc_clk), .Q(d3[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i61.GSR = "ENABLED";
    FD1S3AX d3_i62 (.D(d3_71__N_562[62]), .CK(osc_clk), .Q(d3[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i62.GSR = "ENABLED";
    FD1S3AX d3_i63 (.D(d3_71__N_562[63]), .CK(osc_clk), .Q(d3[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i63.GSR = "ENABLED";
    FD1S3AX d3_i64 (.D(d3_71__N_562[64]), .CK(osc_clk), .Q(d3[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i64.GSR = "ENABLED";
    FD1S3AX d3_i65 (.D(d3_71__N_562[65]), .CK(osc_clk), .Q(d3[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i65.GSR = "ENABLED";
    FD1S3AX d3_i66 (.D(d3_71__N_562[66]), .CK(osc_clk), .Q(d3[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i66.GSR = "ENABLED";
    FD1S3AX d3_i67 (.D(d3_71__N_562[67]), .CK(osc_clk), .Q(d3[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i67.GSR = "ENABLED";
    FD1S3AX d3_i68 (.D(d3_71__N_562[68]), .CK(osc_clk), .Q(d3[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i68.GSR = "ENABLED";
    FD1S3AX d3_i69 (.D(d3_71__N_562[69]), .CK(osc_clk), .Q(d3[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i69.GSR = "ENABLED";
    FD1S3AX d3_i70 (.D(d3_71__N_562[70]), .CK(osc_clk), .Q(d3[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i70.GSR = "ENABLED";
    FD1S3AX d3_i71 (.D(d3_71__N_562[71]), .CK(osc_clk), .Q(d3[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i71.GSR = "ENABLED";
    FD1S3AX d4_i1 (.D(d4_71__N_634[1]), .CK(osc_clk), .Q(d4[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i1.GSR = "ENABLED";
    FD1S3AX d4_i2 (.D(d4_71__N_634[2]), .CK(osc_clk), .Q(d4[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i2.GSR = "ENABLED";
    FD1S3AX d4_i3 (.D(d4_71__N_634[3]), .CK(osc_clk), .Q(d4[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i3.GSR = "ENABLED";
    FD1S3AX d4_i4 (.D(d4_71__N_634[4]), .CK(osc_clk), .Q(d4[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i4.GSR = "ENABLED";
    FD1S3AX d4_i5 (.D(d4_71__N_634[5]), .CK(osc_clk), .Q(d4[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i5.GSR = "ENABLED";
    FD1S3AX d4_i6 (.D(d4_71__N_634[6]), .CK(osc_clk), .Q(d4[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i6.GSR = "ENABLED";
    FD1S3AX d4_i7 (.D(d4_71__N_634[7]), .CK(osc_clk), .Q(d4[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i7.GSR = "ENABLED";
    FD1S3AX d4_i8 (.D(d4_71__N_634[8]), .CK(osc_clk), .Q(d4[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i8.GSR = "ENABLED";
    FD1S3AX d4_i9 (.D(d4_71__N_634[9]), .CK(osc_clk), .Q(d4[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i9.GSR = "ENABLED";
    FD1S3AX d4_i10 (.D(d4_71__N_634[10]), .CK(osc_clk), .Q(d4[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i10.GSR = "ENABLED";
    FD1S3AX d4_i11 (.D(d4_71__N_634[11]), .CK(osc_clk), .Q(d4[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i11.GSR = "ENABLED";
    FD1S3AX d4_i12 (.D(d4_71__N_634[12]), .CK(osc_clk), .Q(d4[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i12.GSR = "ENABLED";
    FD1S3AX d4_i13 (.D(d4_71__N_634[13]), .CK(osc_clk), .Q(d4[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i13.GSR = "ENABLED";
    FD1S3AX d4_i14 (.D(d4_71__N_634[14]), .CK(osc_clk), .Q(d4[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i14.GSR = "ENABLED";
    FD1S3AX d4_i15 (.D(d4_71__N_634[15]), .CK(osc_clk), .Q(d4[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i15.GSR = "ENABLED";
    FD1S3AX d4_i16 (.D(d4_71__N_634[16]), .CK(osc_clk), .Q(d4[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i16.GSR = "ENABLED";
    FD1S3AX d4_i17 (.D(d4_71__N_634[17]), .CK(osc_clk), .Q(d4[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i17.GSR = "ENABLED";
    FD1S3AX d4_i18 (.D(d4_71__N_634[18]), .CK(osc_clk), .Q(d4[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i18.GSR = "ENABLED";
    FD1S3AX d4_i19 (.D(d4_71__N_634[19]), .CK(osc_clk), .Q(d4[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i19.GSR = "ENABLED";
    FD1S3AX d4_i20 (.D(d4_71__N_634[20]), .CK(osc_clk), .Q(d4[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i20.GSR = "ENABLED";
    FD1S3AX d4_i21 (.D(d4_71__N_634[21]), .CK(osc_clk), .Q(d4[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i21.GSR = "ENABLED";
    FD1S3AX d4_i22 (.D(d4_71__N_634[22]), .CK(osc_clk), .Q(d4[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i22.GSR = "ENABLED";
    FD1S3AX d4_i23 (.D(d4_71__N_634[23]), .CK(osc_clk), .Q(d4[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i23.GSR = "ENABLED";
    FD1S3AX d4_i24 (.D(d4_71__N_634[24]), .CK(osc_clk), .Q(d4[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i24.GSR = "ENABLED";
    FD1S3AX d4_i25 (.D(d4_71__N_634[25]), .CK(osc_clk), .Q(d4[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i25.GSR = "ENABLED";
    FD1S3AX d4_i26 (.D(d4_71__N_634[26]), .CK(osc_clk), .Q(d4[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i26.GSR = "ENABLED";
    FD1S3AX d4_i27 (.D(d4_71__N_634[27]), .CK(osc_clk), .Q(d4[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i27.GSR = "ENABLED";
    FD1S3AX d4_i28 (.D(d4_71__N_634[28]), .CK(osc_clk), .Q(d4[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i28.GSR = "ENABLED";
    FD1S3AX d4_i29 (.D(d4_71__N_634[29]), .CK(osc_clk), .Q(d4[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i29.GSR = "ENABLED";
    FD1S3AX d4_i30 (.D(d4_71__N_634[30]), .CK(osc_clk), .Q(d4[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i30.GSR = "ENABLED";
    FD1S3AX d4_i31 (.D(d4_71__N_634[31]), .CK(osc_clk), .Q(d4[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i31.GSR = "ENABLED";
    FD1S3AX d4_i32 (.D(d4_71__N_634[32]), .CK(osc_clk), .Q(d4[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i32.GSR = "ENABLED";
    FD1S3AX d4_i33 (.D(d4_71__N_634[33]), .CK(osc_clk), .Q(d4[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i33.GSR = "ENABLED";
    FD1S3AX d4_i34 (.D(d4_71__N_634[34]), .CK(osc_clk), .Q(d4[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i34.GSR = "ENABLED";
    FD1S3AX d4_i35 (.D(d4_71__N_634[35]), .CK(osc_clk), .Q(d4[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i35.GSR = "ENABLED";
    FD1S3AX d4_i36 (.D(d4_71__N_634[36]), .CK(osc_clk), .Q(d4[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i36.GSR = "ENABLED";
    FD1S3AX d4_i37 (.D(d4_71__N_634[37]), .CK(osc_clk), .Q(d4[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i37.GSR = "ENABLED";
    FD1S3AX d4_i38 (.D(d4_71__N_634[38]), .CK(osc_clk), .Q(d4[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i38.GSR = "ENABLED";
    FD1S3AX d4_i39 (.D(d4_71__N_634[39]), .CK(osc_clk), .Q(d4[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i39.GSR = "ENABLED";
    FD1S3AX d4_i40 (.D(d4_71__N_634[40]), .CK(osc_clk), .Q(d4[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i40.GSR = "ENABLED";
    FD1S3AX d4_i41 (.D(d4_71__N_634[41]), .CK(osc_clk), .Q(d4[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i41.GSR = "ENABLED";
    FD1S3AX d4_i42 (.D(d4_71__N_634[42]), .CK(osc_clk), .Q(d4[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i42.GSR = "ENABLED";
    FD1S3AX d4_i43 (.D(d4_71__N_634[43]), .CK(osc_clk), .Q(d4[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i43.GSR = "ENABLED";
    FD1S3AX d4_i44 (.D(d4_71__N_634[44]), .CK(osc_clk), .Q(d4[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i44.GSR = "ENABLED";
    FD1S3AX d4_i45 (.D(d4_71__N_634[45]), .CK(osc_clk), .Q(d4[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i45.GSR = "ENABLED";
    FD1S3AX d4_i46 (.D(d4_71__N_634[46]), .CK(osc_clk), .Q(d4[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i46.GSR = "ENABLED";
    FD1S3AX d4_i47 (.D(d4_71__N_634[47]), .CK(osc_clk), .Q(d4[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i47.GSR = "ENABLED";
    FD1S3AX d4_i48 (.D(d4_71__N_634[48]), .CK(osc_clk), .Q(d4[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i48.GSR = "ENABLED";
    FD1S3AX d4_i49 (.D(d4_71__N_634[49]), .CK(osc_clk), .Q(d4[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i49.GSR = "ENABLED";
    FD1S3AX d4_i50 (.D(d4_71__N_634[50]), .CK(osc_clk), .Q(d4[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i50.GSR = "ENABLED";
    FD1S3AX d4_i51 (.D(d4_71__N_634[51]), .CK(osc_clk), .Q(d4[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i51.GSR = "ENABLED";
    FD1S3AX d4_i52 (.D(d4_71__N_634[52]), .CK(osc_clk), .Q(d4[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i52.GSR = "ENABLED";
    FD1S3AX d4_i53 (.D(d4_71__N_634[53]), .CK(osc_clk), .Q(d4[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i53.GSR = "ENABLED";
    FD1S3AX d4_i54 (.D(d4_71__N_634[54]), .CK(osc_clk), .Q(d4[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i54.GSR = "ENABLED";
    FD1S3AX d4_i55 (.D(d4_71__N_634[55]), .CK(osc_clk), .Q(d4[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i55.GSR = "ENABLED";
    FD1S3AX d4_i56 (.D(d4_71__N_634[56]), .CK(osc_clk), .Q(d4[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i56.GSR = "ENABLED";
    FD1S3AX d4_i57 (.D(d4_71__N_634[57]), .CK(osc_clk), .Q(d4[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i57.GSR = "ENABLED";
    FD1S3AX d4_i58 (.D(d4_71__N_634[58]), .CK(osc_clk), .Q(d4[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i58.GSR = "ENABLED";
    FD1S3AX d4_i59 (.D(d4_71__N_634[59]), .CK(osc_clk), .Q(d4[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i59.GSR = "ENABLED";
    FD1S3AX d4_i60 (.D(d4_71__N_634[60]), .CK(osc_clk), .Q(d4[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i60.GSR = "ENABLED";
    FD1S3AX d4_i61 (.D(d4_71__N_634[61]), .CK(osc_clk), .Q(d4[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i61.GSR = "ENABLED";
    FD1S3AX d4_i62 (.D(d4_71__N_634[62]), .CK(osc_clk), .Q(d4[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i62.GSR = "ENABLED";
    FD1S3AX d4_i63 (.D(d4_71__N_634[63]), .CK(osc_clk), .Q(d4[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i63.GSR = "ENABLED";
    FD1S3AX d4_i64 (.D(d4_71__N_634[64]), .CK(osc_clk), .Q(d4[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i64.GSR = "ENABLED";
    FD1S3AX d4_i65 (.D(d4_71__N_634[65]), .CK(osc_clk), .Q(d4[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i65.GSR = "ENABLED";
    FD1S3AX d4_i66 (.D(d4_71__N_634[66]), .CK(osc_clk), .Q(d4[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i66.GSR = "ENABLED";
    FD1S3AX d4_i67 (.D(d4_71__N_634[67]), .CK(osc_clk), .Q(d4[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i67.GSR = "ENABLED";
    FD1S3AX d4_i68 (.D(d4_71__N_634[68]), .CK(osc_clk), .Q(d4[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i68.GSR = "ENABLED";
    FD1S3AX d4_i69 (.D(d4_71__N_634[69]), .CK(osc_clk), .Q(d4[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i69.GSR = "ENABLED";
    FD1S3AX d4_i70 (.D(d4_71__N_634[70]), .CK(osc_clk), .Q(d4[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i70.GSR = "ENABLED";
    FD1S3AX d4_i71 (.D(d4_71__N_634[71]), .CK(osc_clk), .Q(d4[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i71.GSR = "ENABLED";
    FD1S3AX d5_i1 (.D(d5_71__N_706[1]), .CK(osc_clk), .Q(d5[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i1.GSR = "ENABLED";
    FD1S3AX d5_i2 (.D(d5_71__N_706[2]), .CK(osc_clk), .Q(d5[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i2.GSR = "ENABLED";
    FD1S3AX d5_i3 (.D(d5_71__N_706[3]), .CK(osc_clk), .Q(d5[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i3.GSR = "ENABLED";
    FD1S3AX d5_i4 (.D(d5_71__N_706[4]), .CK(osc_clk), .Q(d5[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i4.GSR = "ENABLED";
    FD1S3AX d5_i5 (.D(d5_71__N_706[5]), .CK(osc_clk), .Q(d5[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i5.GSR = "ENABLED";
    FD1S3AX d5_i6 (.D(d5_71__N_706[6]), .CK(osc_clk), .Q(d5[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i6.GSR = "ENABLED";
    FD1S3AX d5_i7 (.D(d5_71__N_706[7]), .CK(osc_clk), .Q(d5[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i7.GSR = "ENABLED";
    FD1S3AX d5_i8 (.D(d5_71__N_706[8]), .CK(osc_clk), .Q(d5[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i8.GSR = "ENABLED";
    FD1S3AX d5_i9 (.D(d5_71__N_706[9]), .CK(osc_clk), .Q(d5[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i9.GSR = "ENABLED";
    FD1S3AX d5_i10 (.D(d5_71__N_706[10]), .CK(osc_clk), .Q(d5[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i10.GSR = "ENABLED";
    FD1S3AX d5_i11 (.D(d5_71__N_706[11]), .CK(osc_clk), .Q(d5[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i11.GSR = "ENABLED";
    FD1S3AX d5_i12 (.D(d5_71__N_706[12]), .CK(osc_clk), .Q(d5[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i12.GSR = "ENABLED";
    FD1S3AX d5_i13 (.D(d5_71__N_706[13]), .CK(osc_clk), .Q(d5[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i13.GSR = "ENABLED";
    FD1S3AX d5_i14 (.D(d5_71__N_706[14]), .CK(osc_clk), .Q(d5[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i14.GSR = "ENABLED";
    FD1S3AX d5_i15 (.D(d5_71__N_706[15]), .CK(osc_clk), .Q(d5[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i15.GSR = "ENABLED";
    FD1S3AX d5_i16 (.D(d5_71__N_706[16]), .CK(osc_clk), .Q(d5[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i16.GSR = "ENABLED";
    FD1S3AX d5_i17 (.D(d5_71__N_706[17]), .CK(osc_clk), .Q(d5[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i17.GSR = "ENABLED";
    FD1S3AX d5_i18 (.D(d5_71__N_706[18]), .CK(osc_clk), .Q(d5[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i18.GSR = "ENABLED";
    FD1S3AX d5_i19 (.D(d5_71__N_706[19]), .CK(osc_clk), .Q(d5[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i19.GSR = "ENABLED";
    FD1S3AX d5_i20 (.D(d5_71__N_706[20]), .CK(osc_clk), .Q(d5[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i20.GSR = "ENABLED";
    FD1S3AX d5_i21 (.D(d5_71__N_706[21]), .CK(osc_clk), .Q(d5[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i21.GSR = "ENABLED";
    FD1S3AX d5_i22 (.D(d5_71__N_706[22]), .CK(osc_clk), .Q(d5[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i22.GSR = "ENABLED";
    FD1S3AX d5_i23 (.D(d5_71__N_706[23]), .CK(osc_clk), .Q(d5[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i23.GSR = "ENABLED";
    FD1S3AX d5_i24 (.D(d5_71__N_706[24]), .CK(osc_clk), .Q(d5[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i24.GSR = "ENABLED";
    FD1S3AX d5_i25 (.D(d5_71__N_706[25]), .CK(osc_clk), .Q(d5[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i25.GSR = "ENABLED";
    FD1S3AX d5_i26 (.D(d5_71__N_706[26]), .CK(osc_clk), .Q(d5[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i26.GSR = "ENABLED";
    FD1S3AX d5_i27 (.D(d5_71__N_706[27]), .CK(osc_clk), .Q(d5[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i27.GSR = "ENABLED";
    FD1S3AX d5_i28 (.D(d5_71__N_706[28]), .CK(osc_clk), .Q(d5[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i28.GSR = "ENABLED";
    FD1S3AX d5_i29 (.D(d5_71__N_706[29]), .CK(osc_clk), .Q(d5[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i29.GSR = "ENABLED";
    FD1S3AX d5_i30 (.D(d5_71__N_706[30]), .CK(osc_clk), .Q(d5[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i30.GSR = "ENABLED";
    FD1S3AX d5_i31 (.D(d5_71__N_706[31]), .CK(osc_clk), .Q(d5[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i31.GSR = "ENABLED";
    FD1S3AX d5_i32 (.D(d5_71__N_706[32]), .CK(osc_clk), .Q(d5[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i32.GSR = "ENABLED";
    FD1S3AX d5_i33 (.D(d5_71__N_706[33]), .CK(osc_clk), .Q(d5[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i33.GSR = "ENABLED";
    FD1S3AX d5_i34 (.D(d5_71__N_706[34]), .CK(osc_clk), .Q(d5[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i34.GSR = "ENABLED";
    FD1S3AX d5_i35 (.D(d5_71__N_706[35]), .CK(osc_clk), .Q(d5[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i35.GSR = "ENABLED";
    FD1S3AX d5_i36 (.D(d5_71__N_706[36]), .CK(osc_clk), .Q(d5[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i36.GSR = "ENABLED";
    FD1S3AX d5_i37 (.D(d5_71__N_706[37]), .CK(osc_clk), .Q(d5[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i37.GSR = "ENABLED";
    FD1S3AX d5_i38 (.D(d5_71__N_706[38]), .CK(osc_clk), .Q(d5[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i38.GSR = "ENABLED";
    FD1S3AX d5_i39 (.D(d5_71__N_706[39]), .CK(osc_clk), .Q(d5[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i39.GSR = "ENABLED";
    FD1S3AX d5_i40 (.D(d5_71__N_706[40]), .CK(osc_clk), .Q(d5[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i40.GSR = "ENABLED";
    FD1S3AX d5_i41 (.D(d5_71__N_706[41]), .CK(osc_clk), .Q(d5[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i41.GSR = "ENABLED";
    FD1S3AX d5_i42 (.D(d5_71__N_706[42]), .CK(osc_clk), .Q(d5[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i42.GSR = "ENABLED";
    FD1S3AX d5_i43 (.D(d5_71__N_706[43]), .CK(osc_clk), .Q(d5[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i43.GSR = "ENABLED";
    FD1S3AX d5_i44 (.D(d5_71__N_706[44]), .CK(osc_clk), .Q(d5[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i44.GSR = "ENABLED";
    FD1S3AX d5_i45 (.D(d5_71__N_706[45]), .CK(osc_clk), .Q(d5[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i45.GSR = "ENABLED";
    FD1S3AX d5_i46 (.D(d5_71__N_706[46]), .CK(osc_clk), .Q(d5[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i46.GSR = "ENABLED";
    FD1S3AX d5_i47 (.D(d5_71__N_706[47]), .CK(osc_clk), .Q(d5[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i47.GSR = "ENABLED";
    FD1S3AX d5_i48 (.D(d5_71__N_706[48]), .CK(osc_clk), .Q(d5[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i48.GSR = "ENABLED";
    FD1S3AX d5_i49 (.D(d5_71__N_706[49]), .CK(osc_clk), .Q(d5[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i49.GSR = "ENABLED";
    FD1S3AX d5_i50 (.D(d5_71__N_706[50]), .CK(osc_clk), .Q(d5[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i50.GSR = "ENABLED";
    FD1S3AX d5_i51 (.D(d5_71__N_706[51]), .CK(osc_clk), .Q(d5[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i51.GSR = "ENABLED";
    FD1S3AX d5_i52 (.D(d5_71__N_706[52]), .CK(osc_clk), .Q(d5[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i52.GSR = "ENABLED";
    FD1S3AX d5_i53 (.D(d5_71__N_706[53]), .CK(osc_clk), .Q(d5[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i53.GSR = "ENABLED";
    FD1S3AX d5_i54 (.D(d5_71__N_706[54]), .CK(osc_clk), .Q(d5[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i54.GSR = "ENABLED";
    FD1S3AX d5_i55 (.D(d5_71__N_706[55]), .CK(osc_clk), .Q(d5[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i55.GSR = "ENABLED";
    FD1S3AX d5_i56 (.D(d5_71__N_706[56]), .CK(osc_clk), .Q(d5[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i56.GSR = "ENABLED";
    FD1S3AX d5_i57 (.D(d5_71__N_706[57]), .CK(osc_clk), .Q(d5[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i57.GSR = "ENABLED";
    FD1S3AX d5_i58 (.D(d5_71__N_706[58]), .CK(osc_clk), .Q(d5[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i58.GSR = "ENABLED";
    FD1S3AX d5_i59 (.D(d5_71__N_706[59]), .CK(osc_clk), .Q(d5[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i59.GSR = "ENABLED";
    FD1S3AX d5_i60 (.D(d5_71__N_706[60]), .CK(osc_clk), .Q(d5[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i60.GSR = "ENABLED";
    FD1S3AX d5_i61 (.D(d5_71__N_706[61]), .CK(osc_clk), .Q(d5[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i61.GSR = "ENABLED";
    FD1S3AX d5_i62 (.D(d5_71__N_706[62]), .CK(osc_clk), .Q(d5[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i62.GSR = "ENABLED";
    FD1S3AX d5_i63 (.D(d5_71__N_706[63]), .CK(osc_clk), .Q(d5[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i63.GSR = "ENABLED";
    FD1S3AX d5_i64 (.D(d5_71__N_706[64]), .CK(osc_clk), .Q(d5[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i64.GSR = "ENABLED";
    FD1S3AX d5_i65 (.D(d5_71__N_706[65]), .CK(osc_clk), .Q(d5[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i65.GSR = "ENABLED";
    FD1S3AX d5_i66 (.D(d5_71__N_706[66]), .CK(osc_clk), .Q(d5[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i66.GSR = "ENABLED";
    FD1S3AX d5_i67 (.D(d5_71__N_706[67]), .CK(osc_clk), .Q(d5[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i67.GSR = "ENABLED";
    FD1S3AX d5_i68 (.D(d5_71__N_706[68]), .CK(osc_clk), .Q(d5[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i68.GSR = "ENABLED";
    FD1S3AX d5_i69 (.D(d5_71__N_706[69]), .CK(osc_clk), .Q(d5[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i69.GSR = "ENABLED";
    FD1S3AX d5_i70 (.D(d5_71__N_706[70]), .CK(osc_clk), .Q(d5[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i70.GSR = "ENABLED";
    FD1S3AX d5_i71 (.D(d5_71__N_706[71]), .CK(osc_clk), .Q(d5[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i71.GSR = "ENABLED";
    FD1P3AX d6_i0_i1 (.D(d6_71__N_1459[1]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d6_i0_i2 (.D(d6_71__N_1459[2]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d6_i0_i3 (.D(d6_71__N_1459[3]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d6_i0_i4 (.D(d6_71__N_1459[4]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d6_i0_i5 (.D(d6_71__N_1459[5]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d6_i0_i6 (.D(d6_71__N_1459[6]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d6_i0_i7 (.D(d6_71__N_1459[7]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d6_i0_i8 (.D(d6_71__N_1459[8]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d6_i0_i9 (.D(d6_71__N_1459[9]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d6_i0_i10 (.D(d6_71__N_1459[10]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d6_i0_i11 (.D(d6_71__N_1459[11]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d6_i0_i12 (.D(d6_71__N_1459[12]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d6_i0_i13 (.D(d6_71__N_1459[13]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d6_i0_i14 (.D(d6_71__N_1459[14]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d6_i0_i15 (.D(d6_71__N_1459[15]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d6_i0_i16 (.D(d6_71__N_1459[16]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d6_i0_i17 (.D(d6_71__N_1459[17]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d6_i0_i18 (.D(d6_71__N_1459[18]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d6_i0_i19 (.D(d6_71__N_1459[19]), .SP(osc_clk_enable_834), .CK(osc_clk), 
            .Q(d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d6_i0_i20 (.D(d6_71__N_1459[20]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d6_i0_i21 (.D(d6_71__N_1459[21]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d6_i0_i22 (.D(d6_71__N_1459[22]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d6_i0_i23 (.D(d6_71__N_1459[23]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d6_i0_i24 (.D(d6_71__N_1459[24]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d6_i0_i25 (.D(d6_71__N_1459[25]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d6_i0_i26 (.D(d6_71__N_1459[26]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d6_i0_i27 (.D(d6_71__N_1459[27]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d6_i0_i28 (.D(d6_71__N_1459[28]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d6_i0_i29 (.D(d6_71__N_1459[29]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d6_i0_i30 (.D(d6_71__N_1459[30]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d6_i0_i31 (.D(d6_71__N_1459[31]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d6_i0_i32 (.D(d6_71__N_1459[32]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d6_i0_i33 (.D(d6_71__N_1459[33]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d6_i0_i34 (.D(d6_71__N_1459[34]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d6_i0_i35 (.D(d6_71__N_1459[35]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d6_i0_i36 (.D(d6_71__N_1459[36]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d6_i0_i37 (.D(d6_71__N_1459[37]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d6_i0_i38 (.D(d6_71__N_1459[38]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d6_i0_i39 (.D(d6_71__N_1459[39]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d6_i0_i40 (.D(d6_71__N_1459[40]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d6_i0_i41 (.D(d6_71__N_1459[41]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d6_i0_i42 (.D(d6_71__N_1459[42]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d6_i0_i43 (.D(d6_71__N_1459[43]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d6_i0_i44 (.D(d6_71__N_1459[44]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d6_i0_i45 (.D(d6_71__N_1459[45]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d6_i0_i46 (.D(d6_71__N_1459[46]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d6_i0_i47 (.D(d6_71__N_1459[47]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d6_i0_i48 (.D(d6_71__N_1459[48]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d6_i0_i49 (.D(d6_71__N_1459[49]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d6_i0_i50 (.D(d6_71__N_1459[50]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d6_i0_i51 (.D(d6_71__N_1459[51]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d6_i0_i52 (.D(d6_71__N_1459[52]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d6_i0_i53 (.D(d6_71__N_1459[53]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d6_i0_i54 (.D(d6_71__N_1459[54]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d6_i0_i55 (.D(d6_71__N_1459[55]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d6_i0_i56 (.D(d6_71__N_1459[56]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d6_i0_i57 (.D(d6_71__N_1459[57]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d6_i0_i58 (.D(d6_71__N_1459[58]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d6_i0_i59 (.D(d6_71__N_1459[59]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d6_i0_i60 (.D(d6_71__N_1459[60]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d6_i0_i61 (.D(d6_71__N_1459[61]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d6_i0_i62 (.D(d6_71__N_1459[62]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d6_i0_i63 (.D(d6_71__N_1459[63]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d6_i0_i64 (.D(d6_71__N_1459[64]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d6_i0_i65 (.D(d6_71__N_1459[65]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d6_i0_i66 (.D(d6_71__N_1459[66]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d6_i0_i67 (.D(d6_71__N_1459[67]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d6_i0_i68 (.D(d6_71__N_1459[68]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d6_i0_i69 (.D(d6_71__N_1459[69]), .SP(osc_clk_enable_884), .CK(osc_clk), 
            .Q(d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d6_i0_i70 (.D(d6_71__N_1459[70]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d6_i0_i71 (.D(d6_71__N_1459[71]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i1 (.D(d6[1]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i2 (.D(d6[2]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i3 (.D(d6[3]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i4 (.D(d6[4]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i5 (.D(d6[5]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i6 (.D(d6[6]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i7 (.D(d6[7]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i8 (.D(d6[8]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i9 (.D(d6[9]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i10 (.D(d6[10]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i11 (.D(d6[11]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i12 (.D(d6[12]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i13 (.D(d6[13]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i14 (.D(d6[14]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i15 (.D(d6[15]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i16 (.D(d6[16]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i17 (.D(d6[17]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i18 (.D(d6[18]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i19 (.D(d6[19]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i20 (.D(d6[20]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i21 (.D(d6[21]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i22 (.D(d6[22]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i23 (.D(d6[23]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i24 (.D(d6[24]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i25 (.D(d6[25]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i26 (.D(d6[26]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i27 (.D(d6[27]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i28 (.D(d6[28]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i29 (.D(d6[29]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i30 (.D(d6[30]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i31 (.D(d6[31]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i32 (.D(d6[32]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i33 (.D(d6[33]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i34 (.D(d6[34]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i35 (.D(d6[35]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i36 (.D(d6[36]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i37 (.D(d6[37]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i38 (.D(d6[38]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i39 (.D(d6[39]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i40 (.D(d6[40]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i41 (.D(d6[41]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i42 (.D(d6[42]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i43 (.D(d6[43]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i44 (.D(d6[44]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i45 (.D(d6[45]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i46 (.D(d6[46]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i47 (.D(d6[47]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i48 (.D(d6[48]), .SP(osc_clk_enable_934), .CK(osc_clk), 
            .Q(d_d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i49 (.D(d6[49]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d_d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i50 (.D(d6[50]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d_d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i51 (.D(d6[51]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d_d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i52 (.D(d6[52]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d_d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i53 (.D(d6[53]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d_d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i54 (.D(d6[54]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d_d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i55 (.D(d6[55]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d_d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i56 (.D(d6[56]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d_d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i57 (.D(d6[57]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d_d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i58 (.D(d6[58]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d_d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i59 (.D(d6[59]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d_d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i60 (.D(d6[60]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d_d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i61 (.D(d6[61]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d_d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i62 (.D(d6[62]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d_d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i63 (.D(d6[63]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d_d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i64 (.D(d6[64]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d_d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i65 (.D(d6[65]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d_d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i66 (.D(d6[66]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d_d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i67 (.D(d6[67]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d_d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i68 (.D(d6[68]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d_d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i69 (.D(d6[69]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d_d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i70 (.D(d6[70]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d_d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i71 (.D(d6[71]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d_d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d7_i0_i1 (.D(d7_71__N_1531[1]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d7_i0_i2 (.D(d7_71__N_1531[2]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d7_i0_i3 (.D(d7_71__N_1531[3]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d7_i0_i4 (.D(d7_71__N_1531[4]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d7_i0_i5 (.D(d7_71__N_1531[5]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d7_i0_i6 (.D(d7_71__N_1531[6]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d7_i0_i7 (.D(d7_71__N_1531[7]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d7_i0_i8 (.D(d7_71__N_1531[8]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d7_i0_i9 (.D(d7_71__N_1531[9]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d7_i0_i10 (.D(d7_71__N_1531[10]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d7_i0_i11 (.D(d7_71__N_1531[11]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d7_i0_i12 (.D(d7_71__N_1531[12]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d7_i0_i13 (.D(d7_71__N_1531[13]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d7_i0_i14 (.D(d7_71__N_1531[14]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d7_i0_i15 (.D(d7_71__N_1531[15]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d7_i0_i16 (.D(d7_71__N_1531[16]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d7_i0_i17 (.D(d7_71__N_1531[17]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d7_i0_i18 (.D(d7_71__N_1531[18]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d7_i0_i19 (.D(d7_71__N_1531[19]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d7_i0_i20 (.D(d7_71__N_1531[20]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d7_i0_i21 (.D(d7_71__N_1531[21]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d7_i0_i22 (.D(d7_71__N_1531[22]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d7_i0_i23 (.D(d7_71__N_1531[23]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d7_i0_i24 (.D(d7_71__N_1531[24]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d7_i0_i25 (.D(d7_71__N_1531[25]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d7_i0_i26 (.D(d7_71__N_1531[26]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d7_i0_i27 (.D(d7_71__N_1531[27]), .SP(osc_clk_enable_984), .CK(osc_clk), 
            .Q(d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d7_i0_i28 (.D(d7_71__N_1531[28]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d7_i0_i29 (.D(d7_71__N_1531[29]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d7_i0_i30 (.D(d7_71__N_1531[30]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d7_i0_i31 (.D(d7_71__N_1531[31]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d7_i0_i32 (.D(d7_71__N_1531[32]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d7_i0_i33 (.D(d7_71__N_1531[33]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d7_i0_i34 (.D(d7_71__N_1531[34]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d7_i0_i35 (.D(d7_71__N_1531[35]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d7_i0_i36 (.D(d7_71__N_1531[36]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d7_i0_i37 (.D(d7_71__N_1531[37]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d7_i0_i38 (.D(d7_71__N_1531[38]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d7_i0_i39 (.D(d7_71__N_1531[39]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d7_i0_i40 (.D(d7_71__N_1531[40]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d7_i0_i41 (.D(d7_71__N_1531[41]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d7_i0_i42 (.D(d7_71__N_1531[42]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d7_i0_i43 (.D(d7_71__N_1531[43]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d7_i0_i44 (.D(d7_71__N_1531[44]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d7_i0_i45 (.D(d7_71__N_1531[45]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d7_i0_i46 (.D(d7_71__N_1531[46]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d7_i0_i47 (.D(d7_71__N_1531[47]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d7_i0_i48 (.D(d7_71__N_1531[48]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d7_i0_i49 (.D(d7_71__N_1531[49]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d7_i0_i50 (.D(d7_71__N_1531[50]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d7_i0_i51 (.D(d7_71__N_1531[51]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d7_i0_i52 (.D(d7_71__N_1531[52]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d7_i0_i53 (.D(d7_71__N_1531[53]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d7_i0_i54 (.D(d7_71__N_1531[54]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d7_i0_i55 (.D(d7_71__N_1531[55]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d7_i0_i56 (.D(d7_71__N_1531[56]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d7_i0_i57 (.D(d7_71__N_1531[57]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d7_i0_i58 (.D(d7_71__N_1531[58]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d7_i0_i59 (.D(d7_71__N_1531[59]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d7_i0_i60 (.D(d7_71__N_1531[60]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d7_i0_i61 (.D(d7_71__N_1531[61]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d7_i0_i62 (.D(d7_71__N_1531[62]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d7_i0_i63 (.D(d7_71__N_1531[63]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d7_i0_i64 (.D(d7_71__N_1531[64]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d7_i0_i65 (.D(d7_71__N_1531[65]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d7_i0_i66 (.D(d7_71__N_1531[66]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d7_i0_i67 (.D(d7_71__N_1531[67]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d7_i0_i68 (.D(d7_71__N_1531[68]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d7_i0_i69 (.D(d7_71__N_1531[69]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d7_i0_i70 (.D(d7_71__N_1531[70]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d7_i0_i71 (.D(d7_71__N_1531[71]), .SP(osc_clk_enable_1034), 
            .CK(osc_clk), .Q(d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i1 (.D(d7[1]), .SP(osc_clk_enable_1034), .CK(osc_clk), 
            .Q(d_d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i2 (.D(d7[2]), .SP(osc_clk_enable_1034), .CK(osc_clk), 
            .Q(d_d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i3 (.D(d7[3]), .SP(osc_clk_enable_1034), .CK(osc_clk), 
            .Q(d_d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i4 (.D(d7[4]), .SP(osc_clk_enable_1034), .CK(osc_clk), 
            .Q(d_d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i5 (.D(d7[5]), .SP(osc_clk_enable_1034), .CK(osc_clk), 
            .Q(d_d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i6 (.D(d7[6]), .SP(osc_clk_enable_1034), .CK(osc_clk), 
            .Q(d_d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i7 (.D(d7[7]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i8 (.D(d7[8]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i9 (.D(d7[9]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i10 (.D(d7[10]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i11 (.D(d7[11]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i12 (.D(d7[12]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i13 (.D(d7[13]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i14 (.D(d7[14]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i15 (.D(d7[15]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i16 (.D(d7[16]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i17 (.D(d7[17]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i18 (.D(d7[18]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i19 (.D(d7[19]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i20 (.D(d7[20]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i21 (.D(d7[21]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i22 (.D(d7[22]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i23 (.D(d7[23]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i24 (.D(d7[24]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i25 (.D(d7[25]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i26 (.D(d7[26]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i27 (.D(d7[27]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i28 (.D(d7[28]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i29 (.D(d7[29]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i30 (.D(d7[30]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i31 (.D(d7[31]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i32 (.D(d7[32]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i33 (.D(d7[33]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i34 (.D(d7[34]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i35 (.D(d7[35]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i36 (.D(d7[36]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i37 (.D(d7[37]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i38 (.D(d7[38]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i39 (.D(d7[39]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i40 (.D(d7[40]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i41 (.D(d7[41]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i42 (.D(d7[42]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i43 (.D(d7[43]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i44 (.D(d7[44]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i45 (.D(d7[45]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i46 (.D(d7[46]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i47 (.D(d7[47]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i48 (.D(d7[48]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i49 (.D(d7[49]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i50 (.D(d7[50]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i51 (.D(d7[51]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i52 (.D(d7[52]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i53 (.D(d7[53]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i54 (.D(d7[54]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i55 (.D(d7[55]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i56 (.D(d7[56]), .SP(osc_clk_enable_1084), .CK(osc_clk), 
            .Q(d_d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i57 (.D(d7[57]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d_d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i58 (.D(d7[58]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d_d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i59 (.D(d7[59]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d_d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i60 (.D(d7[60]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d_d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i61 (.D(d7[61]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d_d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i62 (.D(d7[62]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d_d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i63 (.D(d7[63]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d_d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i64 (.D(d7[64]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d_d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i65 (.D(d7[65]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d_d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i66 (.D(d7[66]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d_d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i67 (.D(d7[67]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d_d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i68 (.D(d7[68]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d_d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i69 (.D(d7[69]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d_d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i70 (.D(d7[70]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d_d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i71 (.D(d7[71]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d_d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d8_i0_i1 (.D(d8_71__N_1603[1]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d8_i0_i2 (.D(d8_71__N_1603[2]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d8_i0_i3 (.D(d8_71__N_1603[3]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d8_i0_i4 (.D(d8_71__N_1603[4]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d8_i0_i5 (.D(d8_71__N_1603[5]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d8_i0_i6 (.D(d8_71__N_1603[6]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d8_i0_i7 (.D(d8_71__N_1603[7]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d8_i0_i8 (.D(d8_71__N_1603[8]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d8_i0_i9 (.D(d8_71__N_1603[9]), .SP(osc_clk_enable_1134), .CK(osc_clk), 
            .Q(d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d8_i0_i10 (.D(d8_71__N_1603[10]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d8_i0_i11 (.D(d8_71__N_1603[11]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d8_i0_i12 (.D(d8_71__N_1603[12]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d8_i0_i13 (.D(d8_71__N_1603[13]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d8_i0_i14 (.D(d8_71__N_1603[14]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d8_i0_i15 (.D(d8_71__N_1603[15]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d8_i0_i16 (.D(d8_71__N_1603[16]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d8_i0_i17 (.D(d8_71__N_1603[17]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d8_i0_i18 (.D(d8_71__N_1603[18]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d8_i0_i19 (.D(d8_71__N_1603[19]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d8_i0_i20 (.D(d8_71__N_1603[20]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d8_i0_i21 (.D(d8_71__N_1603[21]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d8_i0_i22 (.D(d8_71__N_1603[22]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d8_i0_i23 (.D(d8_71__N_1603[23]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d8_i0_i24 (.D(d8_71__N_1603[24]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d8_i0_i25 (.D(d8_71__N_1603[25]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d8_i0_i26 (.D(d8_71__N_1603[26]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d8_i0_i27 (.D(d8_71__N_1603[27]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d8_i0_i28 (.D(d8_71__N_1603[28]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d8_i0_i29 (.D(d8_71__N_1603[29]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d8_i0_i30 (.D(d8_71__N_1603[30]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d8_i0_i31 (.D(d8_71__N_1603[31]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d8_i0_i32 (.D(d8_71__N_1603[32]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d8_i0_i33 (.D(d8_71__N_1603[33]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d8_i0_i34 (.D(d8_71__N_1603[34]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d8_i0_i35 (.D(d8_71__N_1603[35]), .SP(osc_clk_enable_1134), 
            .CK(osc_clk), .Q(d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d8_i0_i36 (.D(d8_71__N_1603[36]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d8_i0_i37 (.D(d8_71__N_1603[37]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d8_i0_i38 (.D(d8_71__N_1603[38]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d8_i0_i39 (.D(d8_71__N_1603[39]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d8_i0_i40 (.D(d8_71__N_1603[40]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d8_i0_i41 (.D(d8_71__N_1603[41]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d8_i0_i42 (.D(d8_71__N_1603[42]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d8_i0_i43 (.D(d8_71__N_1603[43]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d8_i0_i44 (.D(d8_71__N_1603[44]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d8_i0_i45 (.D(d8_71__N_1603[45]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d8_i0_i46 (.D(d8_71__N_1603[46]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d8_i0_i47 (.D(d8_71__N_1603[47]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d8_i0_i48 (.D(d8_71__N_1603[48]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d8_i0_i49 (.D(d8_71__N_1603[49]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d8_i0_i50 (.D(d8_71__N_1603[50]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d8_i0_i51 (.D(d8_71__N_1603[51]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d8_i0_i52 (.D(d8_71__N_1603[52]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d8_i0_i53 (.D(d8_71__N_1603[53]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d8_i0_i54 (.D(d8_71__N_1603[54]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d8_i0_i55 (.D(d8_71__N_1603[55]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d8_i0_i56 (.D(d8_71__N_1603[56]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d8_i0_i57 (.D(d8_71__N_1603[57]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d8_i0_i58 (.D(d8_71__N_1603[58]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d8_i0_i59 (.D(d8_71__N_1603[59]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d8_i0_i60 (.D(d8_71__N_1603[60]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d8_i0_i61 (.D(d8_71__N_1603[61]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d8_i0_i62 (.D(d8_71__N_1603[62]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d8_i0_i63 (.D(d8_71__N_1603[63]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d8_i0_i64 (.D(d8_71__N_1603[64]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d8_i0_i65 (.D(d8_71__N_1603[65]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d8_i0_i66 (.D(d8_71__N_1603[66]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d8_i0_i67 (.D(d8_71__N_1603[67]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d8_i0_i68 (.D(d8_71__N_1603[68]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d8_i0_i69 (.D(d8_71__N_1603[69]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d8_i0_i70 (.D(d8_71__N_1603[70]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d8_i0_i71 (.D(d8_71__N_1603[71]), .SP(osc_clk_enable_1184), 
            .CK(osc_clk), .Q(d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i1 (.D(d8[1]), .SP(osc_clk_enable_1184), .CK(osc_clk), 
            .Q(d_d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i2 (.D(d8[2]), .SP(osc_clk_enable_1184), .CK(osc_clk), 
            .Q(d_d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i3 (.D(d8[3]), .SP(osc_clk_enable_1184), .CK(osc_clk), 
            .Q(d_d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i4 (.D(d8[4]), .SP(osc_clk_enable_1184), .CK(osc_clk), 
            .Q(d_d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i5 (.D(d8[5]), .SP(osc_clk_enable_1184), .CK(osc_clk), 
            .Q(d_d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i6 (.D(d8[6]), .SP(osc_clk_enable_1184), .CK(osc_clk), 
            .Q(d_d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i7 (.D(d8[7]), .SP(osc_clk_enable_1184), .CK(osc_clk), 
            .Q(d_d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i8 (.D(d8[8]), .SP(osc_clk_enable_1184), .CK(osc_clk), 
            .Q(d_d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i9 (.D(d8[9]), .SP(osc_clk_enable_1184), .CK(osc_clk), 
            .Q(d_d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i10 (.D(d8[10]), .SP(osc_clk_enable_1184), .CK(osc_clk), 
            .Q(d_d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i11 (.D(d8[11]), .SP(osc_clk_enable_1184), .CK(osc_clk), 
            .Q(d_d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i12 (.D(d8[12]), .SP(osc_clk_enable_1184), .CK(osc_clk), 
            .Q(d_d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i13 (.D(d8[13]), .SP(osc_clk_enable_1184), .CK(osc_clk), 
            .Q(d_d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i14 (.D(d8[14]), .SP(osc_clk_enable_1184), .CK(osc_clk), 
            .Q(d_d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i15 (.D(d8[15]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i16 (.D(d8[16]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i17 (.D(d8[17]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i18 (.D(d8[18]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i19 (.D(d8[19]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i20 (.D(d8[20]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i21 (.D(d8[21]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i22 (.D(d8[22]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i23 (.D(d8[23]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i24 (.D(d8[24]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i25 (.D(d8[25]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i26 (.D(d8[26]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i27 (.D(d8[27]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i28 (.D(d8[28]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i29 (.D(d8[29]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i30 (.D(d8[30]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i31 (.D(d8[31]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i32 (.D(d8[32]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i33 (.D(d8[33]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i34 (.D(d8[34]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i35 (.D(d8[35]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i36 (.D(d8[36]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i37 (.D(d8[37]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i38 (.D(d8[38]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i39 (.D(d8[39]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i40 (.D(d8[40]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i41 (.D(d8[41]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i42 (.D(d8[42]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i43 (.D(d8[43]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i44 (.D(d8[44]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i45 (.D(d8[45]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i46 (.D(d8[46]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i47 (.D(d8[47]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i48 (.D(d8[48]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i49 (.D(d8[49]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i50 (.D(d8[50]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i51 (.D(d8[51]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i52 (.D(d8[52]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i53 (.D(d8[53]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i54 (.D(d8[54]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i55 (.D(d8[55]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i56 (.D(d8[56]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i57 (.D(d8[57]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i58 (.D(d8[58]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i59 (.D(d8[59]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i60 (.D(d8[60]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i61 (.D(d8[61]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i62 (.D(d8[62]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i63 (.D(d8[63]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i64 (.D(d8[64]), .SP(osc_clk_enable_1234), .CK(osc_clk), 
            .Q(d_d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i65 (.D(d8[65]), .SP(osc_clk_enable_1284), .CK(osc_clk), 
            .Q(d_d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i66 (.D(d8[66]), .SP(osc_clk_enable_1284), .CK(osc_clk), 
            .Q(d_d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i67 (.D(d8[67]), .SP(osc_clk_enable_1284), .CK(osc_clk), 
            .Q(d_d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i68 (.D(d8[68]), .SP(osc_clk_enable_1284), .CK(osc_clk), 
            .Q(d_d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i69 (.D(d8[69]), .SP(osc_clk_enable_1284), .CK(osc_clk), 
            .Q(d_d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i70 (.D(d8[70]), .SP(osc_clk_enable_1284), .CK(osc_clk), 
            .Q(d_d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i71 (.D(d8[71]), .SP(osc_clk_enable_1284), .CK(osc_clk), 
            .Q(d_d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d9_i0_i1 (.D(d9_71__N_1675[1]), .SP(osc_clk_enable_1284), .CK(osc_clk), 
            .Q(d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d9_i0_i2 (.D(d9_71__N_1675[2]), .SP(osc_clk_enable_1284), .CK(osc_clk), 
            .Q(d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d9_i0_i3 (.D(d9_71__N_1675[3]), .SP(osc_clk_enable_1284), .CK(osc_clk), 
            .Q(d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d9_i0_i4 (.D(d9_71__N_1675[4]), .SP(osc_clk_enable_1284), .CK(osc_clk), 
            .Q(d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d9_i0_i5 (.D(d9_71__N_1675[5]), .SP(osc_clk_enable_1284), .CK(osc_clk), 
            .Q(d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d9_i0_i6 (.D(d9_71__N_1675[6]), .SP(osc_clk_enable_1284), .CK(osc_clk), 
            .Q(d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d9_i0_i7 (.D(d9_71__N_1675[7]), .SP(osc_clk_enable_1284), .CK(osc_clk), 
            .Q(d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d9_i0_i8 (.D(d9_71__N_1675[8]), .SP(osc_clk_enable_1284), .CK(osc_clk), 
            .Q(d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d9_i0_i9 (.D(d9_71__N_1675[9]), .SP(osc_clk_enable_1284), .CK(osc_clk), 
            .Q(d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d9_i0_i10 (.D(d9_71__N_1675[10]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d9_i0_i11 (.D(d9_71__N_1675[11]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d9_i0_i12 (.D(d9_71__N_1675[12]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d9_i0_i13 (.D(d9_71__N_1675[13]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d9_i0_i14 (.D(d9_71__N_1675[14]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d9_i0_i15 (.D(d9_71__N_1675[15]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d9_i0_i16 (.D(d9_71__N_1675[16]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d9_i0_i17 (.D(d9_71__N_1675[17]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d9_i0_i18 (.D(d9_71__N_1675[18]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d9_i0_i19 (.D(d9_71__N_1675[19]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d9_i0_i20 (.D(d9_71__N_1675[20]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d9_i0_i21 (.D(d9_71__N_1675[21]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d9_i0_i22 (.D(d9_71__N_1675[22]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d9_i0_i23 (.D(d9_71__N_1675[23]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d9_i0_i24 (.D(d9_71__N_1675[24]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d9_i0_i25 (.D(d9_71__N_1675[25]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d9_i0_i26 (.D(d9_71__N_1675[26]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d9_i0_i27 (.D(d9_71__N_1675[27]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d9_i0_i28 (.D(d9_71__N_1675[28]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d9_i0_i29 (.D(d9_71__N_1675[29]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d9_i0_i30 (.D(d9_71__N_1675[30]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d9_i0_i31 (.D(d9_71__N_1675[31]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d9_i0_i32 (.D(d9_71__N_1675[32]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d9_i0_i33 (.D(d9_71__N_1675[33]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d9_i0_i34 (.D(d9_71__N_1675[34]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d9_i0_i35 (.D(d9_71__N_1675[35]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d9_i0_i36 (.D(d9_71__N_1675[36]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d9_i0_i37 (.D(d9_71__N_1675[37]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d9_i0_i38 (.D(d9_71__N_1675[38]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d9_i0_i39 (.D(d9_71__N_1675[39]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d9_i0_i40 (.D(d9_71__N_1675[40]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d9_i0_i41 (.D(d9_71__N_1675[41]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d9_i0_i42 (.D(d9_71__N_1675[42]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d9_i0_i43 (.D(d9_71__N_1675[43]), .SP(osc_clk_enable_1284), 
            .CK(osc_clk), .Q(d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d9_i0_i44 (.D(d9_71__N_1675[44]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d9_i0_i45 (.D(d9_71__N_1675[45]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d9_i0_i46 (.D(d9_71__N_1675[46]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d9_i0_i47 (.D(d9_71__N_1675[47]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d9_i0_i48 (.D(d9_71__N_1675[48]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d9_i0_i49 (.D(d9_71__N_1675[49]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d9_i0_i50 (.D(d9_71__N_1675[50]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d9_i0_i51 (.D(d9_71__N_1675[51]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d9_i0_i52 (.D(d9_71__N_1675[52]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d9_i0_i53 (.D(d9_71__N_1675[53]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d9_i0_i54 (.D(d9_71__N_1675[54]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d9_i0_i55 (.D(d9_71__N_1675[55]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d9_i0_i56 (.D(d9_71__N_1675[56]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d9_i0_i57 (.D(d9_71__N_1675[57]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d9_i0_i58 (.D(d9_71__N_1675[58]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d9_i0_i59 (.D(d9_71__N_1675[59]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d9_i0_i60 (.D(d9_71__N_1675[60]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d9_i0_i61 (.D(d9_71__N_1675[61]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d9_i0_i62 (.D(d9_71__N_1675[62]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d9_i0_i63 (.D(d9_71__N_1675[63]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d9_i0_i64 (.D(d9_71__N_1675[64]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d9_i0_i65 (.D(d9_71__N_1675[65]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d9_i0_i66 (.D(d9_71__N_1675[66]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d9_i0_i67 (.D(d9_71__N_1675[67]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d9_i0_i68 (.D(d9_71__N_1675[68]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d9_i0_i69 (.D(d9_71__N_1675[69]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d9_i0_i70 (.D(d9_71__N_1675[70]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d9_i0_i71 (.D(d9_71__N_1675[71]), .SP(osc_clk_enable_1334), 
            .CK(osc_clk), .Q(d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i1 (.D(d9[1]), .SP(osc_clk_enable_1334), .CK(osc_clk), 
            .Q(d_d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i2 (.D(d9[2]), .SP(osc_clk_enable_1334), .CK(osc_clk), 
            .Q(d_d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i3 (.D(d9[3]), .SP(osc_clk_enable_1334), .CK(osc_clk), 
            .Q(d_d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i4 (.D(d9[4]), .SP(osc_clk_enable_1334), .CK(osc_clk), 
            .Q(d_d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i5 (.D(d9[5]), .SP(osc_clk_enable_1334), .CK(osc_clk), 
            .Q(d_d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i6 (.D(d9[6]), .SP(osc_clk_enable_1334), .CK(osc_clk), 
            .Q(d_d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i7 (.D(d9[7]), .SP(osc_clk_enable_1334), .CK(osc_clk), 
            .Q(d_d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i8 (.D(d9[8]), .SP(osc_clk_enable_1334), .CK(osc_clk), 
            .Q(d_d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i9 (.D(d9[9]), .SP(osc_clk_enable_1334), .CK(osc_clk), 
            .Q(d_d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i10 (.D(d9[10]), .SP(osc_clk_enable_1334), .CK(osc_clk), 
            .Q(d_d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i11 (.D(d9[11]), .SP(osc_clk_enable_1334), .CK(osc_clk), 
            .Q(d_d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i12 (.D(d9[12]), .SP(osc_clk_enable_1334), .CK(osc_clk), 
            .Q(d_d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i13 (.D(d9[13]), .SP(osc_clk_enable_1334), .CK(osc_clk), 
            .Q(d_d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i14 (.D(d9[14]), .SP(osc_clk_enable_1334), .CK(osc_clk), 
            .Q(d_d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i15 (.D(d9[15]), .SP(osc_clk_enable_1334), .CK(osc_clk), 
            .Q(d_d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i16 (.D(d9[16]), .SP(osc_clk_enable_1334), .CK(osc_clk), 
            .Q(d_d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i17 (.D(d9[17]), .SP(osc_clk_enable_1334), .CK(osc_clk), 
            .Q(d_d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i18 (.D(d9[18]), .SP(osc_clk_enable_1334), .CK(osc_clk), 
            .Q(d_d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i19 (.D(d9[19]), .SP(osc_clk_enable_1334), .CK(osc_clk), 
            .Q(d_d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i20 (.D(d9[20]), .SP(osc_clk_enable_1334), .CK(osc_clk), 
            .Q(d_d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i21 (.D(d9[21]), .SP(osc_clk_enable_1334), .CK(osc_clk), 
            .Q(d_d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i22 (.D(d9[22]), .SP(osc_clk_enable_1334), .CK(osc_clk), 
            .Q(d_d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i23 (.D(d9[23]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i24 (.D(d9[24]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i25 (.D(d9[25]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i26 (.D(d9[26]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i27 (.D(d9[27]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i28 (.D(d9[28]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i29 (.D(d9[29]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i30 (.D(d9[30]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i31 (.D(d9[31]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i32 (.D(d9[32]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i33 (.D(d9[33]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i34 (.D(d9[34]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i35 (.D(d9[35]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i36 (.D(d9[36]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i37 (.D(d9[37]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i38 (.D(d9[38]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i39 (.D(d9[39]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i40 (.D(d9[40]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i41 (.D(d9[41]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i42 (.D(d9[42]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i43 (.D(d9[43]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i44 (.D(d9[44]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i45 (.D(d9[45]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i46 (.D(d9[46]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i47 (.D(d9[47]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i48 (.D(d9[48]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i49 (.D(d9[49]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i50 (.D(d9[50]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i51 (.D(d9[51]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i52 (.D(d9[52]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i53 (.D(d9[53]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i54 (.D(d9[54]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i55 (.D(d9[55]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i56 (.D(d9[56]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i57 (.D(d9[57]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i58 (.D(d9[58]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i59 (.D(d9[59]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i60 (.D(d9[60]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i61 (.D(d9[61]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i62 (.D(d9[62]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i63 (.D(d9[63]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i64 (.D(d9[64]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i65 (.D(d9[65]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i66 (.D(d9[66]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i67 (.D(d9[67]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i68 (.D(d9[68]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i69 (.D(d9[69]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i70 (.D(d9[70]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i71 (.D(d9[71]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d_d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d10__i2 (.D(d10_71__N_1747[57]), .SP(osc_clk_enable_1384), .CK(osc_clk), 
            .Q(d10[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i2.GSR = "ENABLED";
    FD1P3AX d10__i3 (.D(d10_71__N_1747[58]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i3.GSR = "ENABLED";
    FD1P3AX d10__i4 (.D(d10_71__N_1747[59]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[59] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i4.GSR = "ENABLED";
    FD1P3AX d10__i5 (.D(d10_71__N_1747[60]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[60] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i5.GSR = "ENABLED";
    FD1P3AX d10__i6 (.D(d10_71__N_1747[61]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[61] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i6.GSR = "ENABLED";
    FD1P3AX d10__i7 (.D(d10_71__N_1747[62]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[62] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i7.GSR = "ENABLED";
    FD1P3AX d10__i8 (.D(d10_71__N_1747[63]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[63] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i8.GSR = "ENABLED";
    FD1P3AX d10__i9 (.D(d10_71__N_1747[64]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[64] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i9.GSR = "ENABLED";
    FD1P3AX d10__i10 (.D(d10_71__N_1747[65]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[65] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i10.GSR = "ENABLED";
    FD1P3AX d10__i11 (.D(d10_71__N_1747[66]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[66] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i11.GSR = "ENABLED";
    FD1P3AX d10__i12 (.D(d10_71__N_1747[67]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[67] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i12.GSR = "ENABLED";
    FD1P3AX d10__i13 (.D(d10_71__N_1747[68]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[68] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i13.GSR = "ENABLED";
    FD1P3AX d10__i14 (.D(d10_71__N_1747[69]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[69] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i14.GSR = "ENABLED";
    FD1P3AX d10__i15 (.D(d10_71__N_1747[70]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[70] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i15.GSR = "ENABLED";
    FD1P3AX d10__i16 (.D(d10_71__N_1747[71]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[71] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i16.GSR = "ENABLED";
    FD1P3AX d_out_i0_i1 (.D(d_out_11__N_1819[1]), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i1.GSR = "ENABLED";
    FD1P3AX d_out_i0_i2 (.D(\d_out_11__N_1819[2] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i2.GSR = "ENABLED";
    FD1P3AX d_out_i0_i3 (.D(\d_out_11__N_1819[3] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i3.GSR = "ENABLED";
    FD1P3AX d_out_i0_i4 (.D(\d_out_11__N_1819[4] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i4.GSR = "ENABLED";
    FD1P3AX d_out_i0_i5 (.D(\d_out_11__N_1819[5] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i5.GSR = "ENABLED";
    FD1P3AX d_out_i0_i6 (.D(\d_out_11__N_1819[6] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i6.GSR = "ENABLED";
    FD1P3AX d_out_i0_i7 (.D(\d_out_11__N_1819[7] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i7.GSR = "ENABLED";
    FD1P3AX d_out_i0_i8 (.D(\d_out_11__N_1819[8] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i8.GSR = "ENABLED";
    FD1P3AX d_out_i0_i9 (.D(\d_out_11__N_1819[9] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i9.GSR = "ENABLED";
    FD1P3AX d_out_i0_i10 (.D(\d_out_11__N_1819[10] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i10.GSR = "ENABLED";
    FD1P3AX d_out_i0_i11 (.D(\d_out_11__N_1819[11] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i11.GSR = "ENABLED";
    FD1S3AX d1_i1 (.D(d1_71__N_418[1]), .CK(osc_clk), .Q(d1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i1.GSR = "ENABLED";
    FD1S3AX d1_i2 (.D(d1_71__N_418[2]), .CK(osc_clk), .Q(d1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i2.GSR = "ENABLED";
    FD1S3AX d1_i3 (.D(d1_71__N_418[3]), .CK(osc_clk), .Q(d1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i3.GSR = "ENABLED";
    FD1S3AX d1_i4 (.D(d1_71__N_418[4]), .CK(osc_clk), .Q(d1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i4.GSR = "ENABLED";
    FD1S3AX d1_i5 (.D(d1_71__N_418[5]), .CK(osc_clk), .Q(d1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i5.GSR = "ENABLED";
    FD1S3AX d1_i6 (.D(d1_71__N_418[6]), .CK(osc_clk), .Q(d1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i6.GSR = "ENABLED";
    FD1S3AX d1_i7 (.D(d1_71__N_418[7]), .CK(osc_clk), .Q(d1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i7.GSR = "ENABLED";
    FD1S3AX d1_i8 (.D(d1_71__N_418[8]), .CK(osc_clk), .Q(d1[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i8.GSR = "ENABLED";
    FD1S3AX d1_i9 (.D(d1_71__N_418[9]), .CK(osc_clk), .Q(d1[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i9.GSR = "ENABLED";
    FD1S3AX d1_i10 (.D(d1_71__N_418[10]), .CK(osc_clk), .Q(d1[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i10.GSR = "ENABLED";
    FD1S3AX d1_i11 (.D(d1_71__N_418[11]), .CK(osc_clk), .Q(d1[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i11.GSR = "ENABLED";
    FD1S3AX d1_i12 (.D(d1_71__N_418[12]), .CK(osc_clk), .Q(d1[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i12.GSR = "ENABLED";
    FD1S3AX d1_i13 (.D(d1_71__N_418[13]), .CK(osc_clk), .Q(d1[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i13.GSR = "ENABLED";
    FD1S3AX d1_i14 (.D(d1_71__N_418[14]), .CK(osc_clk), .Q(d1[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i14.GSR = "ENABLED";
    FD1S3AX d1_i15 (.D(d1_71__N_418[15]), .CK(osc_clk), .Q(d1[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i15.GSR = "ENABLED";
    FD1S3AX d1_i16 (.D(d1_71__N_418[16]), .CK(osc_clk), .Q(d1[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i16.GSR = "ENABLED";
    FD1S3AX d1_i17 (.D(d1_71__N_418[17]), .CK(osc_clk), .Q(d1[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i17.GSR = "ENABLED";
    FD1S3AX d1_i18 (.D(d1_71__N_418[18]), .CK(osc_clk), .Q(d1[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i18.GSR = "ENABLED";
    FD1S3AX d1_i19 (.D(d1_71__N_418[19]), .CK(osc_clk), .Q(d1[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i19.GSR = "ENABLED";
    FD1S3AX d1_i20 (.D(d1_71__N_418[20]), .CK(osc_clk), .Q(d1[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i20.GSR = "ENABLED";
    FD1S3AX d1_i21 (.D(d1_71__N_418[21]), .CK(osc_clk), .Q(d1[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i21.GSR = "ENABLED";
    FD1S3AX d1_i22 (.D(d1_71__N_418[22]), .CK(osc_clk), .Q(d1[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i22.GSR = "ENABLED";
    FD1S3AX d1_i23 (.D(d1_71__N_418[23]), .CK(osc_clk), .Q(d1[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i23.GSR = "ENABLED";
    FD1S3AX d1_i24 (.D(d1_71__N_418[24]), .CK(osc_clk), .Q(d1[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i24.GSR = "ENABLED";
    FD1S3AX d1_i25 (.D(d1_71__N_418[25]), .CK(osc_clk), .Q(d1[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i25.GSR = "ENABLED";
    FD1S3AX d1_i26 (.D(d1_71__N_418[26]), .CK(osc_clk), .Q(d1[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i26.GSR = "ENABLED";
    FD1S3AX d1_i27 (.D(d1_71__N_418[27]), .CK(osc_clk), .Q(d1[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i27.GSR = "ENABLED";
    FD1S3AX d1_i28 (.D(d1_71__N_418[28]), .CK(osc_clk), .Q(d1[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i28.GSR = "ENABLED";
    FD1S3AX d1_i29 (.D(d1_71__N_418[29]), .CK(osc_clk), .Q(d1[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i29.GSR = "ENABLED";
    FD1S3AX d1_i30 (.D(d1_71__N_418[30]), .CK(osc_clk), .Q(d1[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i30.GSR = "ENABLED";
    FD1S3AX d1_i31 (.D(d1_71__N_418[31]), .CK(osc_clk), .Q(d1[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i31.GSR = "ENABLED";
    FD1S3AX d1_i32 (.D(d1_71__N_418[32]), .CK(osc_clk), .Q(d1[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i32.GSR = "ENABLED";
    FD1S3AX d1_i33 (.D(d1_71__N_418[33]), .CK(osc_clk), .Q(d1[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i33.GSR = "ENABLED";
    FD1S3AX d1_i34 (.D(d1_71__N_418[34]), .CK(osc_clk), .Q(d1[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i34.GSR = "ENABLED";
    FD1S3AX d1_i35 (.D(d1_71__N_418[35]), .CK(osc_clk), .Q(d1[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i35.GSR = "ENABLED";
    FD1S3AX d1_i36 (.D(d1_71__N_418[36]), .CK(osc_clk), .Q(d1[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i36.GSR = "ENABLED";
    FD1S3AX d1_i37 (.D(d1_71__N_418[37]), .CK(osc_clk), .Q(d1[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i37.GSR = "ENABLED";
    FD1S3AX d1_i38 (.D(d1_71__N_418[38]), .CK(osc_clk), .Q(d1[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i38.GSR = "ENABLED";
    FD1S3AX d1_i39 (.D(d1_71__N_418[39]), .CK(osc_clk), .Q(d1[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i39.GSR = "ENABLED";
    FD1S3AX d1_i40 (.D(d1_71__N_418[40]), .CK(osc_clk), .Q(d1[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i40.GSR = "ENABLED";
    FD1S3AX d1_i41 (.D(d1_71__N_418[41]), .CK(osc_clk), .Q(d1[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i41.GSR = "ENABLED";
    FD1S3AX d1_i42 (.D(d1_71__N_418[42]), .CK(osc_clk), .Q(d1[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i42.GSR = "ENABLED";
    FD1S3AX d1_i43 (.D(d1_71__N_418[43]), .CK(osc_clk), .Q(d1[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i43.GSR = "ENABLED";
    FD1S3AX d1_i44 (.D(d1_71__N_418[44]), .CK(osc_clk), .Q(d1[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i44.GSR = "ENABLED";
    FD1S3AX d1_i45 (.D(d1_71__N_418[45]), .CK(osc_clk), .Q(d1[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i45.GSR = "ENABLED";
    FD1S3AX d1_i46 (.D(d1_71__N_418[46]), .CK(osc_clk), .Q(d1[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i46.GSR = "ENABLED";
    FD1S3AX d1_i47 (.D(d1_71__N_418[47]), .CK(osc_clk), .Q(d1[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i47.GSR = "ENABLED";
    FD1S3AX d1_i48 (.D(d1_71__N_418[48]), .CK(osc_clk), .Q(d1[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i48.GSR = "ENABLED";
    FD1S3AX d1_i49 (.D(d1_71__N_418[49]), .CK(osc_clk), .Q(d1[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i49.GSR = "ENABLED";
    FD1S3AX d1_i50 (.D(d1_71__N_418[50]), .CK(osc_clk), .Q(d1[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i50.GSR = "ENABLED";
    FD1S3AX d1_i51 (.D(d1_71__N_418[51]), .CK(osc_clk), .Q(d1[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i51.GSR = "ENABLED";
    FD1S3AX d1_i52 (.D(d1_71__N_418[52]), .CK(osc_clk), .Q(d1[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i52.GSR = "ENABLED";
    FD1S3AX d1_i53 (.D(d1_71__N_418[53]), .CK(osc_clk), .Q(d1[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i53.GSR = "ENABLED";
    FD1S3AX d1_i54 (.D(d1_71__N_418[54]), .CK(osc_clk), .Q(d1[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i54.GSR = "ENABLED";
    FD1S3AX d1_i55 (.D(d1_71__N_418[55]), .CK(osc_clk), .Q(d1[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i55.GSR = "ENABLED";
    FD1S3AX d1_i56 (.D(d1_71__N_418[56]), .CK(osc_clk), .Q(d1[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i56.GSR = "ENABLED";
    FD1S3AX d1_i57 (.D(d1_71__N_418[57]), .CK(osc_clk), .Q(d1[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i57.GSR = "ENABLED";
    FD1S3AX d1_i58 (.D(d1_71__N_418[58]), .CK(osc_clk), .Q(d1[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i58.GSR = "ENABLED";
    FD1S3AX d1_i59 (.D(d1_71__N_418[59]), .CK(osc_clk), .Q(d1[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i59.GSR = "ENABLED";
    FD1S3AX d1_i60 (.D(d1_71__N_418[60]), .CK(osc_clk), .Q(d1[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i60.GSR = "ENABLED";
    FD1S3AX d1_i61 (.D(d1_71__N_418[61]), .CK(osc_clk), .Q(d1[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i61.GSR = "ENABLED";
    FD1S3AX d1_i62 (.D(d1_71__N_418[62]), .CK(osc_clk), .Q(d1[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i62.GSR = "ENABLED";
    FD1S3AX d1_i63 (.D(d1_71__N_418[63]), .CK(osc_clk), .Q(d1[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i63.GSR = "ENABLED";
    FD1S3AX d1_i64 (.D(d1_71__N_418[64]), .CK(osc_clk), .Q(d1[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i64.GSR = "ENABLED";
    FD1S3AX d1_i65 (.D(d1_71__N_418[65]), .CK(osc_clk), .Q(d1[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i65.GSR = "ENABLED";
    FD1S3AX d1_i66 (.D(d1_71__N_418[66]), .CK(osc_clk), .Q(d1[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i66.GSR = "ENABLED";
    FD1S3AX d1_i67 (.D(d1_71__N_418[67]), .CK(osc_clk), .Q(d1[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i67.GSR = "ENABLED";
    FD1S3AX d1_i68 (.D(d1_71__N_418[68]), .CK(osc_clk), .Q(d1[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i68.GSR = "ENABLED";
    FD1S3AX d1_i69 (.D(d1_71__N_418[69]), .CK(osc_clk), .Q(d1[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i69.GSR = "ENABLED";
    FD1S3AX d1_i70 (.D(d1_71__N_418[70]), .CK(osc_clk), .Q(d1[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i70.GSR = "ENABLED";
    FD1S3AX d1_i71 (.D(d1_71__N_418[71]), .CK(osc_clk), .Q(d1[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i71.GSR = "ENABLED";
    CCU2D add_1104_9 (.A0(d_tmp[43]), .B0(d_d_tmp[43]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[44]), .B1(d_d_tmp[44]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11609), .COUT(n11610), .S0(n6101[7]), 
          .S1(n6101[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1104_9.INIT0 = 16'h5999;
    defparam add_1104_9.INIT1 = 16'h5999;
    defparam add_1104_9.INJECT1_0 = "NO";
    defparam add_1104_9.INJECT1_1 = "NO";
    CCU2D add_1104_7 (.A0(d_tmp[41]), .B0(d_d_tmp[41]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[42]), .B1(d_d_tmp[42]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11608), .COUT(n11609), .S0(n6101[5]), 
          .S1(n6101[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1104_7.INIT0 = 16'h5999;
    defparam add_1104_7.INIT1 = 16'h5999;
    defparam add_1104_7.INJECT1_0 = "NO";
    defparam add_1104_7.INJECT1_1 = "NO";
    CCU2D add_1104_5 (.A0(d_tmp[39]), .B0(d_d_tmp[39]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[40]), .B1(d_d_tmp[40]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11607), .COUT(n11608), .S0(n6101[3]), 
          .S1(n6101[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1104_5.INIT0 = 16'h5999;
    defparam add_1104_5.INIT1 = 16'h5999;
    defparam add_1104_5.INJECT1_0 = "NO";
    defparam add_1104_5.INJECT1_1 = "NO";
    CCU2D add_1104_3 (.A0(d_tmp[37]), .B0(d_d_tmp[37]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[38]), .B1(d_d_tmp[38]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11606), .COUT(n11607), .S0(n6101[1]), 
          .S1(n6101[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1104_3.INIT0 = 16'h5999;
    defparam add_1104_3.INIT1 = 16'h5999;
    defparam add_1104_3.INJECT1_0 = "NO";
    defparam add_1104_3.INJECT1_1 = "NO";
    CCU2D add_1104_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[36]), .B1(d_d_tmp[36]), .C1(GND_net), .D1(GND_net), 
          .COUT(n11606), .S1(n6101[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1104_1.INIT0 = 16'hF000;
    defparam add_1104_1.INIT1 = 16'h5999;
    defparam add_1104_1.INJECT1_0 = "NO";
    defparam add_1104_1.INJECT1_1 = "NO";
    CCU2D add_1105_37 (.A0(d_d_tmp[70]), .B0(n6100), .C0(n6101[34]), .D0(d_tmp[70]), 
          .A1(d_d_tmp[71]), .B1(n6100), .C1(n6101[35]), .D1(d_tmp[71]), 
          .CIN(n11604), .S0(d6_71__N_1459[70]), .S1(d6_71__N_1459[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1105_37.INIT0 = 16'hb874;
    defparam add_1105_37.INIT1 = 16'hb874;
    defparam add_1105_37.INJECT1_0 = "NO";
    defparam add_1105_37.INJECT1_1 = "NO";
    CCU2D add_1105_35 (.A0(d_d_tmp[68]), .B0(n6100), .C0(n6101[32]), .D0(d_tmp[68]), 
          .A1(d_d_tmp[69]), .B1(n6100), .C1(n6101[33]), .D1(d_tmp[69]), 
          .CIN(n11603), .COUT(n11604), .S0(d6_71__N_1459[68]), .S1(d6_71__N_1459[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1105_35.INIT0 = 16'hb874;
    defparam add_1105_35.INIT1 = 16'hb874;
    defparam add_1105_35.INJECT1_0 = "NO";
    defparam add_1105_35.INJECT1_1 = "NO";
    CCU2D add_1105_33 (.A0(d_d_tmp[66]), .B0(n6100), .C0(n6101[30]), .D0(d_tmp[66]), 
          .A1(d_d_tmp[67]), .B1(n6100), .C1(n6101[31]), .D1(d_tmp[67]), 
          .CIN(n11602), .COUT(n11603), .S0(d6_71__N_1459[66]), .S1(d6_71__N_1459[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1105_33.INIT0 = 16'hb874;
    defparam add_1105_33.INIT1 = 16'hb874;
    defparam add_1105_33.INJECT1_0 = "NO";
    defparam add_1105_33.INJECT1_1 = "NO";
    CCU2D add_1105_31 (.A0(d_d_tmp[64]), .B0(n6100), .C0(n6101[28]), .D0(d_tmp[64]), 
          .A1(d_d_tmp[65]), .B1(n6100), .C1(n6101[29]), .D1(d_tmp[65]), 
          .CIN(n11601), .COUT(n11602), .S0(d6_71__N_1459[64]), .S1(d6_71__N_1459[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1105_31.INIT0 = 16'hb874;
    defparam add_1105_31.INIT1 = 16'hb874;
    defparam add_1105_31.INJECT1_0 = "NO";
    defparam add_1105_31.INJECT1_1 = "NO";
    CCU2D add_1105_29 (.A0(d_d_tmp[62]), .B0(n6100), .C0(n6101[26]), .D0(d_tmp[62]), 
          .A1(d_d_tmp[63]), .B1(n6100), .C1(n6101[27]), .D1(d_tmp[63]), 
          .CIN(n11600), .COUT(n11601), .S0(d6_71__N_1459[62]), .S1(d6_71__N_1459[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1105_29.INIT0 = 16'hb874;
    defparam add_1105_29.INIT1 = 16'hb874;
    defparam add_1105_29.INJECT1_0 = "NO";
    defparam add_1105_29.INJECT1_1 = "NO";
    CCU2D add_1105_27 (.A0(d_d_tmp[60]), .B0(n6100), .C0(n6101[24]), .D0(d_tmp[60]), 
          .A1(d_d_tmp[61]), .B1(n6100), .C1(n6101[25]), .D1(d_tmp[61]), 
          .CIN(n11599), .COUT(n11600), .S0(d6_71__N_1459[60]), .S1(d6_71__N_1459[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1105_27.INIT0 = 16'hb874;
    defparam add_1105_27.INIT1 = 16'hb874;
    defparam add_1105_27.INJECT1_0 = "NO";
    defparam add_1105_27.INJECT1_1 = "NO";
    CCU2D add_1105_25 (.A0(d_d_tmp[58]), .B0(n6100), .C0(n6101[22]), .D0(d_tmp[58]), 
          .A1(d_d_tmp[59]), .B1(n6100), .C1(n6101[23]), .D1(d_tmp[59]), 
          .CIN(n11598), .COUT(n11599), .S0(d6_71__N_1459[58]), .S1(d6_71__N_1459[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1105_25.INIT0 = 16'hb874;
    defparam add_1105_25.INIT1 = 16'hb874;
    defparam add_1105_25.INJECT1_0 = "NO";
    defparam add_1105_25.INJECT1_1 = "NO";
    CCU2D add_1105_23 (.A0(d_d_tmp[56]), .B0(n6100), .C0(n6101[20]), .D0(d_tmp[56]), 
          .A1(d_d_tmp[57]), .B1(n6100), .C1(n6101[21]), .D1(d_tmp[57]), 
          .CIN(n11597), .COUT(n11598), .S0(d6_71__N_1459[56]), .S1(d6_71__N_1459[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1105_23.INIT0 = 16'hb874;
    defparam add_1105_23.INIT1 = 16'hb874;
    defparam add_1105_23.INJECT1_0 = "NO";
    defparam add_1105_23.INJECT1_1 = "NO";
    CCU2D add_1105_21 (.A0(d_d_tmp[54]), .B0(n6100), .C0(n6101[18]), .D0(d_tmp[54]), 
          .A1(d_d_tmp[55]), .B1(n6100), .C1(n6101[19]), .D1(d_tmp[55]), 
          .CIN(n11596), .COUT(n11597), .S0(d6_71__N_1459[54]), .S1(d6_71__N_1459[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1105_21.INIT0 = 16'hb874;
    defparam add_1105_21.INIT1 = 16'hb874;
    defparam add_1105_21.INJECT1_0 = "NO";
    defparam add_1105_21.INJECT1_1 = "NO";
    CCU2D add_1105_19 (.A0(d_d_tmp[52]), .B0(n6100), .C0(n6101[16]), .D0(d_tmp[52]), 
          .A1(d_d_tmp[53]), .B1(n6100), .C1(n6101[17]), .D1(d_tmp[53]), 
          .CIN(n11595), .COUT(n11596), .S0(d6_71__N_1459[52]), .S1(d6_71__N_1459[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1105_19.INIT0 = 16'hb874;
    defparam add_1105_19.INIT1 = 16'hb874;
    defparam add_1105_19.INJECT1_0 = "NO";
    defparam add_1105_19.INJECT1_1 = "NO";
    CCU2D add_1105_17 (.A0(d_d_tmp[50]), .B0(n6100), .C0(n6101[14]), .D0(d_tmp[50]), 
          .A1(d_d_tmp[51]), .B1(n6100), .C1(n6101[15]), .D1(d_tmp[51]), 
          .CIN(n11594), .COUT(n11595), .S0(d6_71__N_1459[50]), .S1(d6_71__N_1459[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1105_17.INIT0 = 16'hb874;
    defparam add_1105_17.INIT1 = 16'hb874;
    defparam add_1105_17.INJECT1_0 = "NO";
    defparam add_1105_17.INJECT1_1 = "NO";
    CCU2D add_1105_15 (.A0(d_d_tmp[48]), .B0(n6100), .C0(n6101[12]), .D0(d_tmp[48]), 
          .A1(d_d_tmp[49]), .B1(n6100), .C1(n6101[13]), .D1(d_tmp[49]), 
          .CIN(n11593), .COUT(n11594), .S0(d6_71__N_1459[48]), .S1(d6_71__N_1459[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1105_15.INIT0 = 16'hb874;
    defparam add_1105_15.INIT1 = 16'hb874;
    defparam add_1105_15.INJECT1_0 = "NO";
    defparam add_1105_15.INJECT1_1 = "NO";
    CCU2D add_1105_13 (.A0(d_d_tmp[46]), .B0(n6100), .C0(n6101[10]), .D0(d_tmp[46]), 
          .A1(d_d_tmp[47]), .B1(n6100), .C1(n6101[11]), .D1(d_tmp[47]), 
          .CIN(n11592), .COUT(n11593), .S0(d6_71__N_1459[46]), .S1(d6_71__N_1459[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1105_13.INIT0 = 16'hb874;
    defparam add_1105_13.INIT1 = 16'hb874;
    defparam add_1105_13.INJECT1_0 = "NO";
    defparam add_1105_13.INJECT1_1 = "NO";
    CCU2D add_1105_11 (.A0(d_d_tmp[44]), .B0(n6100), .C0(n6101[8]), .D0(d_tmp[44]), 
          .A1(d_d_tmp[45]), .B1(n6100), .C1(n6101[9]), .D1(d_tmp[45]), 
          .CIN(n11591), .COUT(n11592), .S0(d6_71__N_1459[44]), .S1(d6_71__N_1459[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1105_11.INIT0 = 16'hb874;
    defparam add_1105_11.INIT1 = 16'hb874;
    defparam add_1105_11.INJECT1_0 = "NO";
    defparam add_1105_11.INJECT1_1 = "NO";
    CCU2D add_1105_9 (.A0(d_d_tmp[42]), .B0(n6100), .C0(n6101[6]), .D0(d_tmp[42]), 
          .A1(d_d_tmp[43]), .B1(n6100), .C1(n6101[7]), .D1(d_tmp[43]), 
          .CIN(n11590), .COUT(n11591), .S0(d6_71__N_1459[42]), .S1(d6_71__N_1459[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1105_9.INIT0 = 16'hb874;
    defparam add_1105_9.INIT1 = 16'hb874;
    defparam add_1105_9.INJECT1_0 = "NO";
    defparam add_1105_9.INJECT1_1 = "NO";
    CCU2D add_1105_7 (.A0(d_d_tmp[40]), .B0(n6100), .C0(n6101[4]), .D0(d_tmp[40]), 
          .A1(d_d_tmp[41]), .B1(n6100), .C1(n6101[5]), .D1(d_tmp[41]), 
          .CIN(n11589), .COUT(n11590), .S0(d6_71__N_1459[40]), .S1(d6_71__N_1459[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1105_7.INIT0 = 16'hb874;
    defparam add_1105_7.INIT1 = 16'hb874;
    defparam add_1105_7.INJECT1_0 = "NO";
    defparam add_1105_7.INJECT1_1 = "NO";
    CCU2D add_1105_5 (.A0(d_d_tmp[38]), .B0(n6100), .C0(n6101[2]), .D0(d_tmp[38]), 
          .A1(d_d_tmp[39]), .B1(n6100), .C1(n6101[3]), .D1(d_tmp[39]), 
          .CIN(n11588), .COUT(n11589), .S0(d6_71__N_1459[38]), .S1(d6_71__N_1459[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1105_5.INIT0 = 16'hb874;
    defparam add_1105_5.INIT1 = 16'hb874;
    defparam add_1105_5.INJECT1_0 = "NO";
    defparam add_1105_5.INJECT1_1 = "NO";
    CCU2D add_1105_3 (.A0(d_d_tmp[36]), .B0(n6100), .C0(n6101[0]), .D0(d_tmp[36]), 
          .A1(d_d_tmp[37]), .B1(n6100), .C1(n6101[1]), .D1(d_tmp[37]), 
          .CIN(n11587), .COUT(n11588), .S0(d6_71__N_1459[36]), .S1(d6_71__N_1459[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1105_3.INIT0 = 16'hb874;
    defparam add_1105_3.INIT1 = 16'hb874;
    defparam add_1105_3.INJECT1_0 = "NO";
    defparam add_1105_3.INJECT1_1 = "NO";
    CCU2D add_1105_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n6100), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11587));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1105_1.INIT0 = 16'hF000;
    defparam add_1105_1.INIT1 = 16'h0555;
    defparam add_1105_1.INJECT1_0 = "NO";
    defparam add_1105_1.INJECT1_1 = "NO";
    CCU2D add_1109_37 (.A0(d6[71]), .B0(d_d6[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11583), 
          .S0(n6253[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1109_37.INIT0 = 16'h5999;
    defparam add_1109_37.INIT1 = 16'h0000;
    defparam add_1109_37.INJECT1_0 = "NO";
    defparam add_1109_37.INJECT1_1 = "NO";
    CCU2D add_1109_35 (.A0(d6[69]), .B0(d_d6[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[70]), .B1(d_d6[70]), .C1(GND_net), .D1(GND_net), .CIN(n11582), 
          .COUT(n11583), .S0(n6253[33]), .S1(n6253[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1109_35.INIT0 = 16'h5999;
    defparam add_1109_35.INIT1 = 16'h5999;
    defparam add_1109_35.INJECT1_0 = "NO";
    defparam add_1109_35.INJECT1_1 = "NO";
    CCU2D add_1109_33 (.A0(d6[67]), .B0(d_d6[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[68]), .B1(d_d6[68]), .C1(GND_net), .D1(GND_net), .CIN(n11581), 
          .COUT(n11582), .S0(n6253[31]), .S1(n6253[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1109_33.INIT0 = 16'h5999;
    defparam add_1109_33.INIT1 = 16'h5999;
    defparam add_1109_33.INJECT1_0 = "NO";
    defparam add_1109_33.INJECT1_1 = "NO";
    CCU2D add_1109_31 (.A0(d6[65]), .B0(d_d6[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[66]), .B1(d_d6[66]), .C1(GND_net), .D1(GND_net), .CIN(n11580), 
          .COUT(n11581), .S0(n6253[29]), .S1(n6253[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1109_31.INIT0 = 16'h5999;
    defparam add_1109_31.INIT1 = 16'h5999;
    defparam add_1109_31.INJECT1_0 = "NO";
    defparam add_1109_31.INJECT1_1 = "NO";
    CCU2D add_1109_29 (.A0(d6[63]), .B0(d_d6[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[64]), .B1(d_d6[64]), .C1(GND_net), .D1(GND_net), .CIN(n11579), 
          .COUT(n11580), .S0(n6253[27]), .S1(n6253[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1109_29.INIT0 = 16'h5999;
    defparam add_1109_29.INIT1 = 16'h5999;
    defparam add_1109_29.INJECT1_0 = "NO";
    defparam add_1109_29.INJECT1_1 = "NO";
    CCU2D add_1109_27 (.A0(d6[61]), .B0(d_d6[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[62]), .B1(d_d6[62]), .C1(GND_net), .D1(GND_net), .CIN(n11578), 
          .COUT(n11579), .S0(n6253[25]), .S1(n6253[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1109_27.INIT0 = 16'h5999;
    defparam add_1109_27.INIT1 = 16'h5999;
    defparam add_1109_27.INJECT1_0 = "NO";
    defparam add_1109_27.INJECT1_1 = "NO";
    CCU2D add_1109_25 (.A0(d6[59]), .B0(d_d6[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[60]), .B1(d_d6[60]), .C1(GND_net), .D1(GND_net), .CIN(n11577), 
          .COUT(n11578), .S0(n6253[23]), .S1(n6253[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1109_25.INIT0 = 16'h5999;
    defparam add_1109_25.INIT1 = 16'h5999;
    defparam add_1109_25.INJECT1_0 = "NO";
    defparam add_1109_25.INJECT1_1 = "NO";
    CCU2D add_1109_23 (.A0(d6[57]), .B0(d_d6[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[58]), .B1(d_d6[58]), .C1(GND_net), .D1(GND_net), .CIN(n11576), 
          .COUT(n11577), .S0(n6253[21]), .S1(n6253[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1109_23.INIT0 = 16'h5999;
    defparam add_1109_23.INIT1 = 16'h5999;
    defparam add_1109_23.INJECT1_0 = "NO";
    defparam add_1109_23.INJECT1_1 = "NO";
    CCU2D add_1109_21 (.A0(d6[55]), .B0(d_d6[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[56]), .B1(d_d6[56]), .C1(GND_net), .D1(GND_net), .CIN(n11575), 
          .COUT(n11576), .S0(n6253[19]), .S1(n6253[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1109_21.INIT0 = 16'h5999;
    defparam add_1109_21.INIT1 = 16'h5999;
    defparam add_1109_21.INJECT1_0 = "NO";
    defparam add_1109_21.INJECT1_1 = "NO";
    CCU2D add_1109_19 (.A0(d6[53]), .B0(d_d6[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[54]), .B1(d_d6[54]), .C1(GND_net), .D1(GND_net), .CIN(n11574), 
          .COUT(n11575), .S0(n6253[17]), .S1(n6253[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1109_19.INIT0 = 16'h5999;
    defparam add_1109_19.INIT1 = 16'h5999;
    defparam add_1109_19.INJECT1_0 = "NO";
    defparam add_1109_19.INJECT1_1 = "NO";
    CCU2D add_1109_17 (.A0(d6[51]), .B0(d_d6[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[52]), .B1(d_d6[52]), .C1(GND_net), .D1(GND_net), .CIN(n11573), 
          .COUT(n11574), .S0(n6253[15]), .S1(n6253[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1109_17.INIT0 = 16'h5999;
    defparam add_1109_17.INIT1 = 16'h5999;
    defparam add_1109_17.INJECT1_0 = "NO";
    defparam add_1109_17.INJECT1_1 = "NO";
    CCU2D add_1109_15 (.A0(d6[49]), .B0(d_d6[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[50]), .B1(d_d6[50]), .C1(GND_net), .D1(GND_net), .CIN(n11572), 
          .COUT(n11573), .S0(n6253[13]), .S1(n6253[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1109_15.INIT0 = 16'h5999;
    defparam add_1109_15.INIT1 = 16'h5999;
    defparam add_1109_15.INJECT1_0 = "NO";
    defparam add_1109_15.INJECT1_1 = "NO";
    CCU2D add_1109_13 (.A0(d6[47]), .B0(d_d6[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[48]), .B1(d_d6[48]), .C1(GND_net), .D1(GND_net), .CIN(n11571), 
          .COUT(n11572), .S0(n6253[11]), .S1(n6253[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1109_13.INIT0 = 16'h5999;
    defparam add_1109_13.INIT1 = 16'h5999;
    defparam add_1109_13.INJECT1_0 = "NO";
    defparam add_1109_13.INJECT1_1 = "NO";
    CCU2D add_1109_11 (.A0(d6[45]), .B0(d_d6[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[46]), .B1(d_d6[46]), .C1(GND_net), .D1(GND_net), .CIN(n11570), 
          .COUT(n11571), .S0(n6253[9]), .S1(n6253[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1109_11.INIT0 = 16'h5999;
    defparam add_1109_11.INIT1 = 16'h5999;
    defparam add_1109_11.INJECT1_0 = "NO";
    defparam add_1109_11.INJECT1_1 = "NO";
    CCU2D add_1109_9 (.A0(d6[43]), .B0(d_d6[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[44]), .B1(d_d6[44]), .C1(GND_net), .D1(GND_net), .CIN(n11569), 
          .COUT(n11570), .S0(n6253[7]), .S1(n6253[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1109_9.INIT0 = 16'h5999;
    defparam add_1109_9.INIT1 = 16'h5999;
    defparam add_1109_9.INJECT1_0 = "NO";
    defparam add_1109_9.INJECT1_1 = "NO";
    CCU2D add_1109_7 (.A0(d6[41]), .B0(d_d6[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[42]), .B1(d_d6[42]), .C1(GND_net), .D1(GND_net), .CIN(n11568), 
          .COUT(n11569), .S0(n6253[5]), .S1(n6253[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1109_7.INIT0 = 16'h5999;
    defparam add_1109_7.INIT1 = 16'h5999;
    defparam add_1109_7.INJECT1_0 = "NO";
    defparam add_1109_7.INJECT1_1 = "NO";
    CCU2D add_1109_5 (.A0(d6[39]), .B0(d_d6[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[40]), .B1(d_d6[40]), .C1(GND_net), .D1(GND_net), .CIN(n11567), 
          .COUT(n11568), .S0(n6253[3]), .S1(n6253[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1109_5.INIT0 = 16'h5999;
    defparam add_1109_5.INIT1 = 16'h5999;
    defparam add_1109_5.INJECT1_0 = "NO";
    defparam add_1109_5.INJECT1_1 = "NO";
    CCU2D add_1109_3 (.A0(d6[37]), .B0(d_d6[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[38]), .B1(d_d6[38]), .C1(GND_net), .D1(GND_net), .CIN(n11566), 
          .COUT(n11567), .S0(n6253[1]), .S1(n6253[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1109_3.INIT0 = 16'h5999;
    defparam add_1109_3.INIT1 = 16'h5999;
    defparam add_1109_3.INJECT1_0 = "NO";
    defparam add_1109_3.INJECT1_1 = "NO";
    CCU2D add_1109_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d6[36]), .B1(d_d6[36]), .C1(GND_net), .D1(GND_net), .COUT(n11566), 
          .S1(n6253[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1109_1.INIT0 = 16'hF000;
    defparam add_1109_1.INIT1 = 16'h5999;
    defparam add_1109_1.INJECT1_0 = "NO";
    defparam add_1109_1.INJECT1_1 = "NO";
    CCU2D add_1110_37 (.A0(d_d6[70]), .B0(n6252), .C0(n6253[34]), .D0(d6[70]), 
          .A1(d_d6[71]), .B1(n6252), .C1(n6253[35]), .D1(d6[71]), .CIN(n11564), 
          .S0(d7_71__N_1531[70]), .S1(d7_71__N_1531[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1110_37.INIT0 = 16'hb874;
    defparam add_1110_37.INIT1 = 16'hb874;
    defparam add_1110_37.INJECT1_0 = "NO";
    defparam add_1110_37.INJECT1_1 = "NO";
    CCU2D add_1110_35 (.A0(d_d6[68]), .B0(n6252), .C0(n6253[32]), .D0(d6[68]), 
          .A1(d_d6[69]), .B1(n6252), .C1(n6253[33]), .D1(d6[69]), .CIN(n11563), 
          .COUT(n11564), .S0(d7_71__N_1531[68]), .S1(d7_71__N_1531[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1110_35.INIT0 = 16'hb874;
    defparam add_1110_35.INIT1 = 16'hb874;
    defparam add_1110_35.INJECT1_0 = "NO";
    defparam add_1110_35.INJECT1_1 = "NO";
    CCU2D add_1110_33 (.A0(d_d6[66]), .B0(n6252), .C0(n6253[30]), .D0(d6[66]), 
          .A1(d_d6[67]), .B1(n6252), .C1(n6253[31]), .D1(d6[67]), .CIN(n11562), 
          .COUT(n11563), .S0(d7_71__N_1531[66]), .S1(d7_71__N_1531[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1110_33.INIT0 = 16'hb874;
    defparam add_1110_33.INIT1 = 16'hb874;
    defparam add_1110_33.INJECT1_0 = "NO";
    defparam add_1110_33.INJECT1_1 = "NO";
    CCU2D add_1110_31 (.A0(d_d6[64]), .B0(n6252), .C0(n6253[28]), .D0(d6[64]), 
          .A1(d_d6[65]), .B1(n6252), .C1(n6253[29]), .D1(d6[65]), .CIN(n11561), 
          .COUT(n11562), .S0(d7_71__N_1531[64]), .S1(d7_71__N_1531[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1110_31.INIT0 = 16'hb874;
    defparam add_1110_31.INIT1 = 16'hb874;
    defparam add_1110_31.INJECT1_0 = "NO";
    defparam add_1110_31.INJECT1_1 = "NO";
    CCU2D add_1110_29 (.A0(d_d6[62]), .B0(n6252), .C0(n6253[26]), .D0(d6[62]), 
          .A1(d_d6[63]), .B1(n6252), .C1(n6253[27]), .D1(d6[63]), .CIN(n11560), 
          .COUT(n11561), .S0(d7_71__N_1531[62]), .S1(d7_71__N_1531[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1110_29.INIT0 = 16'hb874;
    defparam add_1110_29.INIT1 = 16'hb874;
    defparam add_1110_29.INJECT1_0 = "NO";
    defparam add_1110_29.INJECT1_1 = "NO";
    CCU2D add_1110_27 (.A0(d_d6[60]), .B0(n6252), .C0(n6253[24]), .D0(d6[60]), 
          .A1(d_d6[61]), .B1(n6252), .C1(n6253[25]), .D1(d6[61]), .CIN(n11559), 
          .COUT(n11560), .S0(d7_71__N_1531[60]), .S1(d7_71__N_1531[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1110_27.INIT0 = 16'hb874;
    defparam add_1110_27.INIT1 = 16'hb874;
    defparam add_1110_27.INJECT1_0 = "NO";
    defparam add_1110_27.INJECT1_1 = "NO";
    CCU2D add_1110_25 (.A0(d_d6[58]), .B0(n6252), .C0(n6253[22]), .D0(d6[58]), 
          .A1(d_d6[59]), .B1(n6252), .C1(n6253[23]), .D1(d6[59]), .CIN(n11558), 
          .COUT(n11559), .S0(d7_71__N_1531[58]), .S1(d7_71__N_1531[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1110_25.INIT0 = 16'hb874;
    defparam add_1110_25.INIT1 = 16'hb874;
    defparam add_1110_25.INJECT1_0 = "NO";
    defparam add_1110_25.INJECT1_1 = "NO";
    CCU2D add_1110_23 (.A0(d_d6[56]), .B0(n6252), .C0(n6253[20]), .D0(d6[56]), 
          .A1(d_d6[57]), .B1(n6252), .C1(n6253[21]), .D1(d6[57]), .CIN(n11557), 
          .COUT(n11558), .S0(d7_71__N_1531[56]), .S1(d7_71__N_1531[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1110_23.INIT0 = 16'hb874;
    defparam add_1110_23.INIT1 = 16'hb874;
    defparam add_1110_23.INJECT1_0 = "NO";
    defparam add_1110_23.INJECT1_1 = "NO";
    CCU2D add_1110_21 (.A0(d_d6[54]), .B0(n6252), .C0(n6253[18]), .D0(d6[54]), 
          .A1(d_d6[55]), .B1(n6252), .C1(n6253[19]), .D1(d6[55]), .CIN(n11556), 
          .COUT(n11557), .S0(d7_71__N_1531[54]), .S1(d7_71__N_1531[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1110_21.INIT0 = 16'hb874;
    defparam add_1110_21.INIT1 = 16'hb874;
    defparam add_1110_21.INJECT1_0 = "NO";
    defparam add_1110_21.INJECT1_1 = "NO";
    CCU2D add_1110_19 (.A0(d_d6[52]), .B0(n6252), .C0(n6253[16]), .D0(d6[52]), 
          .A1(d_d6[53]), .B1(n6252), .C1(n6253[17]), .D1(d6[53]), .CIN(n11555), 
          .COUT(n11556), .S0(d7_71__N_1531[52]), .S1(d7_71__N_1531[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1110_19.INIT0 = 16'hb874;
    defparam add_1110_19.INIT1 = 16'hb874;
    defparam add_1110_19.INJECT1_0 = "NO";
    defparam add_1110_19.INJECT1_1 = "NO";
    CCU2D add_1110_17 (.A0(d_d6[50]), .B0(n6252), .C0(n6253[14]), .D0(d6[50]), 
          .A1(d_d6[51]), .B1(n6252), .C1(n6253[15]), .D1(d6[51]), .CIN(n11554), 
          .COUT(n11555), .S0(d7_71__N_1531[50]), .S1(d7_71__N_1531[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1110_17.INIT0 = 16'hb874;
    defparam add_1110_17.INIT1 = 16'hb874;
    defparam add_1110_17.INJECT1_0 = "NO";
    defparam add_1110_17.INJECT1_1 = "NO";
    CCU2D add_1110_15 (.A0(d_d6[48]), .B0(n6252), .C0(n6253[12]), .D0(d6[48]), 
          .A1(d_d6[49]), .B1(n6252), .C1(n6253[13]), .D1(d6[49]), .CIN(n11553), 
          .COUT(n11554), .S0(d7_71__N_1531[48]), .S1(d7_71__N_1531[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1110_15.INIT0 = 16'hb874;
    defparam add_1110_15.INIT1 = 16'hb874;
    defparam add_1110_15.INJECT1_0 = "NO";
    defparam add_1110_15.INJECT1_1 = "NO";
    CCU2D add_1110_13 (.A0(d_d6[46]), .B0(n6252), .C0(n6253[10]), .D0(d6[46]), 
          .A1(d_d6[47]), .B1(n6252), .C1(n6253[11]), .D1(d6[47]), .CIN(n11552), 
          .COUT(n11553), .S0(d7_71__N_1531[46]), .S1(d7_71__N_1531[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1110_13.INIT0 = 16'hb874;
    defparam add_1110_13.INIT1 = 16'hb874;
    defparam add_1110_13.INJECT1_0 = "NO";
    defparam add_1110_13.INJECT1_1 = "NO";
    CCU2D add_1110_11 (.A0(d_d6[44]), .B0(n6252), .C0(n6253[8]), .D0(d6[44]), 
          .A1(d_d6[45]), .B1(n6252), .C1(n6253[9]), .D1(d6[45]), .CIN(n11551), 
          .COUT(n11552), .S0(d7_71__N_1531[44]), .S1(d7_71__N_1531[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1110_11.INIT0 = 16'hb874;
    defparam add_1110_11.INIT1 = 16'hb874;
    defparam add_1110_11.INJECT1_0 = "NO";
    defparam add_1110_11.INJECT1_1 = "NO";
    CCU2D add_1110_9 (.A0(d_d6[42]), .B0(n6252), .C0(n6253[6]), .D0(d6[42]), 
          .A1(d_d6[43]), .B1(n6252), .C1(n6253[7]), .D1(d6[43]), .CIN(n11550), 
          .COUT(n11551), .S0(d7_71__N_1531[42]), .S1(d7_71__N_1531[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1110_9.INIT0 = 16'hb874;
    defparam add_1110_9.INIT1 = 16'hb874;
    defparam add_1110_9.INJECT1_0 = "NO";
    defparam add_1110_9.INJECT1_1 = "NO";
    CCU2D add_1110_7 (.A0(d_d6[40]), .B0(n6252), .C0(n6253[4]), .D0(d6[40]), 
          .A1(d_d6[41]), .B1(n6252), .C1(n6253[5]), .D1(d6[41]), .CIN(n11549), 
          .COUT(n11550), .S0(d7_71__N_1531[40]), .S1(d7_71__N_1531[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1110_7.INIT0 = 16'hb874;
    defparam add_1110_7.INIT1 = 16'hb874;
    defparam add_1110_7.INJECT1_0 = "NO";
    defparam add_1110_7.INJECT1_1 = "NO";
    CCU2D add_1110_5 (.A0(d_d6[38]), .B0(n6252), .C0(n6253[2]), .D0(d6[38]), 
          .A1(d_d6[39]), .B1(n6252), .C1(n6253[3]), .D1(d6[39]), .CIN(n11548), 
          .COUT(n11549), .S0(d7_71__N_1531[38]), .S1(d7_71__N_1531[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1110_5.INIT0 = 16'hb874;
    defparam add_1110_5.INIT1 = 16'hb874;
    defparam add_1110_5.INJECT1_0 = "NO";
    defparam add_1110_5.INJECT1_1 = "NO";
    LUT4 i4942_2_lut (.A(d4[36]), .B(d5[36]), .Z(n5645[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4942_2_lut.init = 16'h6666;
    LUT4 i4913_2_lut (.A(d1[0]), .B(d2[0]), .Z(d2_71__N_490[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4913_2_lut.init = 16'h6666;
    CCU2D add_1110_3 (.A0(d_d6[36]), .B0(n6252), .C0(n6253[0]), .D0(d6[36]), 
          .A1(d_d6[37]), .B1(n6252), .C1(n6253[1]), .D1(d6[37]), .CIN(n11547), 
          .COUT(n11548), .S0(d7_71__N_1531[36]), .S1(d7_71__N_1531[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1110_3.INIT0 = 16'hb874;
    defparam add_1110_3.INIT1 = 16'hb874;
    defparam add_1110_3.INJECT1_0 = "NO";
    defparam add_1110_3.INJECT1_1 = "NO";
    CCU2D add_1110_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n6252), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11547));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1110_1.INIT0 = 16'hF000;
    defparam add_1110_1.INIT1 = 16'h0555;
    defparam add_1110_1.INJECT1_0 = "NO";
    defparam add_1110_1.INJECT1_1 = "NO";
    CCU2D add_1114_37 (.A0(d7[71]), .B0(d_d7[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11543), 
          .S0(n6405[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1114_37.INIT0 = 16'h5999;
    defparam add_1114_37.INIT1 = 16'h0000;
    defparam add_1114_37.INJECT1_0 = "NO";
    defparam add_1114_37.INJECT1_1 = "NO";
    CCU2D add_1114_35 (.A0(d7[69]), .B0(d_d7[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[70]), .B1(d_d7[70]), .C1(GND_net), .D1(GND_net), .CIN(n11542), 
          .COUT(n11543), .S0(n6405[33]), .S1(n6405[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1114_35.INIT0 = 16'h5999;
    defparam add_1114_35.INIT1 = 16'h5999;
    defparam add_1114_35.INJECT1_0 = "NO";
    defparam add_1114_35.INJECT1_1 = "NO";
    CCU2D add_1114_33 (.A0(d7[67]), .B0(d_d7[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[68]), .B1(d_d7[68]), .C1(GND_net), .D1(GND_net), .CIN(n11541), 
          .COUT(n11542), .S0(n6405[31]), .S1(n6405[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1114_33.INIT0 = 16'h5999;
    defparam add_1114_33.INIT1 = 16'h5999;
    defparam add_1114_33.INJECT1_0 = "NO";
    defparam add_1114_33.INJECT1_1 = "NO";
    CCU2D add_1114_31 (.A0(d7[65]), .B0(d_d7[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[66]), .B1(d_d7[66]), .C1(GND_net), .D1(GND_net), .CIN(n11540), 
          .COUT(n11541), .S0(n6405[29]), .S1(n6405[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1114_31.INIT0 = 16'h5999;
    defparam add_1114_31.INIT1 = 16'h5999;
    defparam add_1114_31.INJECT1_0 = "NO";
    defparam add_1114_31.INJECT1_1 = "NO";
    CCU2D add_1114_29 (.A0(d7[63]), .B0(d_d7[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[64]), .B1(d_d7[64]), .C1(GND_net), .D1(GND_net), .CIN(n11539), 
          .COUT(n11540), .S0(n6405[27]), .S1(n6405[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1114_29.INIT0 = 16'h5999;
    defparam add_1114_29.INIT1 = 16'h5999;
    defparam add_1114_29.INJECT1_0 = "NO";
    defparam add_1114_29.INJECT1_1 = "NO";
    CCU2D add_1114_27 (.A0(d7[61]), .B0(d_d7[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[62]), .B1(d_d7[62]), .C1(GND_net), .D1(GND_net), .CIN(n11538), 
          .COUT(n11539), .S0(n6405[25]), .S1(n6405[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1114_27.INIT0 = 16'h5999;
    defparam add_1114_27.INIT1 = 16'h5999;
    defparam add_1114_27.INJECT1_0 = "NO";
    defparam add_1114_27.INJECT1_1 = "NO";
    CCU2D add_1114_25 (.A0(d7[59]), .B0(d_d7[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[60]), .B1(d_d7[60]), .C1(GND_net), .D1(GND_net), .CIN(n11537), 
          .COUT(n11538), .S0(n6405[23]), .S1(n6405[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1114_25.INIT0 = 16'h5999;
    defparam add_1114_25.INIT1 = 16'h5999;
    defparam add_1114_25.INJECT1_0 = "NO";
    defparam add_1114_25.INJECT1_1 = "NO";
    CCU2D add_1114_23 (.A0(d7[57]), .B0(d_d7[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[58]), .B1(d_d7[58]), .C1(GND_net), .D1(GND_net), .CIN(n11536), 
          .COUT(n11537), .S0(n6405[21]), .S1(n6405[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1114_23.INIT0 = 16'h5999;
    defparam add_1114_23.INIT1 = 16'h5999;
    defparam add_1114_23.INJECT1_0 = "NO";
    defparam add_1114_23.INJECT1_1 = "NO";
    CCU2D add_1114_21 (.A0(d7[55]), .B0(d_d7[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[56]), .B1(d_d7[56]), .C1(GND_net), .D1(GND_net), .CIN(n11535), 
          .COUT(n11536), .S0(n6405[19]), .S1(n6405[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1114_21.INIT0 = 16'h5999;
    defparam add_1114_21.INIT1 = 16'h5999;
    defparam add_1114_21.INJECT1_0 = "NO";
    defparam add_1114_21.INJECT1_1 = "NO";
    CCU2D add_1114_19 (.A0(d7[53]), .B0(d_d7[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[54]), .B1(d_d7[54]), .C1(GND_net), .D1(GND_net), .CIN(n11534), 
          .COUT(n11535), .S0(n6405[17]), .S1(n6405[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1114_19.INIT0 = 16'h5999;
    defparam add_1114_19.INIT1 = 16'h5999;
    defparam add_1114_19.INJECT1_0 = "NO";
    defparam add_1114_19.INJECT1_1 = "NO";
    CCU2D add_1114_17 (.A0(d7[51]), .B0(d_d7[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[52]), .B1(d_d7[52]), .C1(GND_net), .D1(GND_net), .CIN(n11533), 
          .COUT(n11534), .S0(n6405[15]), .S1(n6405[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1114_17.INIT0 = 16'h5999;
    defparam add_1114_17.INIT1 = 16'h5999;
    defparam add_1114_17.INJECT1_0 = "NO";
    defparam add_1114_17.INJECT1_1 = "NO";
    CCU2D add_1114_15 (.A0(d7[49]), .B0(d_d7[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[50]), .B1(d_d7[50]), .C1(GND_net), .D1(GND_net), .CIN(n11532), 
          .COUT(n11533), .S0(n6405[13]), .S1(n6405[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1114_15.INIT0 = 16'h5999;
    defparam add_1114_15.INIT1 = 16'h5999;
    defparam add_1114_15.INJECT1_0 = "NO";
    defparam add_1114_15.INJECT1_1 = "NO";
    CCU2D add_1114_13 (.A0(d7[47]), .B0(d_d7[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[48]), .B1(d_d7[48]), .C1(GND_net), .D1(GND_net), .CIN(n11531), 
          .COUT(n11532), .S0(n6405[11]), .S1(n6405[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1114_13.INIT0 = 16'h5999;
    defparam add_1114_13.INIT1 = 16'h5999;
    defparam add_1114_13.INJECT1_0 = "NO";
    defparam add_1114_13.INJECT1_1 = "NO";
    CCU2D add_1114_11 (.A0(d7[45]), .B0(d_d7[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[46]), .B1(d_d7[46]), .C1(GND_net), .D1(GND_net), .CIN(n11530), 
          .COUT(n11531), .S0(n6405[9]), .S1(n6405[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1114_11.INIT0 = 16'h5999;
    defparam add_1114_11.INIT1 = 16'h5999;
    defparam add_1114_11.INJECT1_0 = "NO";
    defparam add_1114_11.INJECT1_1 = "NO";
    CCU2D add_1114_9 (.A0(d7[43]), .B0(d_d7[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[44]), .B1(d_d7[44]), .C1(GND_net), .D1(GND_net), .CIN(n11529), 
          .COUT(n11530), .S0(n6405[7]), .S1(n6405[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1114_9.INIT0 = 16'h5999;
    defparam add_1114_9.INIT1 = 16'h5999;
    defparam add_1114_9.INJECT1_0 = "NO";
    defparam add_1114_9.INJECT1_1 = "NO";
    CCU2D add_1114_7 (.A0(d7[41]), .B0(d_d7[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[42]), .B1(d_d7[42]), .C1(GND_net), .D1(GND_net), .CIN(n11528), 
          .COUT(n11529), .S0(n6405[5]), .S1(n6405[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1114_7.INIT0 = 16'h5999;
    defparam add_1114_7.INIT1 = 16'h5999;
    defparam add_1114_7.INJECT1_0 = "NO";
    defparam add_1114_7.INJECT1_1 = "NO";
    CCU2D add_1114_5 (.A0(d7[39]), .B0(d_d7[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[40]), .B1(d_d7[40]), .C1(GND_net), .D1(GND_net), .CIN(n11527), 
          .COUT(n11528), .S0(n6405[3]), .S1(n6405[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1114_5.INIT0 = 16'h5999;
    defparam add_1114_5.INIT1 = 16'h5999;
    defparam add_1114_5.INJECT1_0 = "NO";
    defparam add_1114_5.INJECT1_1 = "NO";
    CCU2D add_1114_3 (.A0(d7[37]), .B0(d_d7[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[38]), .B1(d_d7[38]), .C1(GND_net), .D1(GND_net), .CIN(n11526), 
          .COUT(n11527), .S0(n6405[1]), .S1(n6405[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1114_3.INIT0 = 16'h5999;
    defparam add_1114_3.INIT1 = 16'h5999;
    defparam add_1114_3.INJECT1_0 = "NO";
    defparam add_1114_3.INJECT1_1 = "NO";
    CCU2D add_1114_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d7[36]), .B1(d_d7[36]), .C1(GND_net), .D1(GND_net), .COUT(n11526), 
          .S1(n6405[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1114_1.INIT0 = 16'hF000;
    defparam add_1114_1.INIT1 = 16'h5999;
    defparam add_1114_1.INJECT1_0 = "NO";
    defparam add_1114_1.INJECT1_1 = "NO";
    CCU2D add_1115_37 (.A0(d_d7[70]), .B0(n6404), .C0(n6405[34]), .D0(d7[70]), 
          .A1(d_d7[71]), .B1(n6404), .C1(n6405[35]), .D1(d7[71]), .CIN(n11524), 
          .S0(d8_71__N_1603[70]), .S1(d8_71__N_1603[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1115_37.INIT0 = 16'hb874;
    defparam add_1115_37.INIT1 = 16'hb874;
    defparam add_1115_37.INJECT1_0 = "NO";
    defparam add_1115_37.INJECT1_1 = "NO";
    CCU2D add_1115_35 (.A0(d_d7[68]), .B0(n6404), .C0(n6405[32]), .D0(d7[68]), 
          .A1(d_d7[69]), .B1(n6404), .C1(n6405[33]), .D1(d7[69]), .CIN(n11523), 
          .COUT(n11524), .S0(d8_71__N_1603[68]), .S1(d8_71__N_1603[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1115_35.INIT0 = 16'hb874;
    defparam add_1115_35.INIT1 = 16'hb874;
    defparam add_1115_35.INJECT1_0 = "NO";
    defparam add_1115_35.INJECT1_1 = "NO";
    CCU2D add_1115_33 (.A0(d_d7[66]), .B0(n6404), .C0(n6405[30]), .D0(d7[66]), 
          .A1(d_d7[67]), .B1(n6404), .C1(n6405[31]), .D1(d7[67]), .CIN(n11522), 
          .COUT(n11523), .S0(d8_71__N_1603[66]), .S1(d8_71__N_1603[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1115_33.INIT0 = 16'hb874;
    defparam add_1115_33.INIT1 = 16'hb874;
    defparam add_1115_33.INJECT1_0 = "NO";
    defparam add_1115_33.INJECT1_1 = "NO";
    CCU2D add_1115_31 (.A0(d_d7[64]), .B0(n6404), .C0(n6405[28]), .D0(d7[64]), 
          .A1(d_d7[65]), .B1(n6404), .C1(n6405[29]), .D1(d7[65]), .CIN(n11521), 
          .COUT(n11522), .S0(d8_71__N_1603[64]), .S1(d8_71__N_1603[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1115_31.INIT0 = 16'hb874;
    defparam add_1115_31.INIT1 = 16'hb874;
    defparam add_1115_31.INJECT1_0 = "NO";
    defparam add_1115_31.INJECT1_1 = "NO";
    CCU2D add_1115_29 (.A0(d_d7[62]), .B0(n6404), .C0(n6405[26]), .D0(d7[62]), 
          .A1(d_d7[63]), .B1(n6404), .C1(n6405[27]), .D1(d7[63]), .CIN(n11520), 
          .COUT(n11521), .S0(d8_71__N_1603[62]), .S1(d8_71__N_1603[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1115_29.INIT0 = 16'hb874;
    defparam add_1115_29.INIT1 = 16'hb874;
    defparam add_1115_29.INJECT1_0 = "NO";
    defparam add_1115_29.INJECT1_1 = "NO";
    CCU2D add_1115_27 (.A0(d_d7[60]), .B0(n6404), .C0(n6405[24]), .D0(d7[60]), 
          .A1(d_d7[61]), .B1(n6404), .C1(n6405[25]), .D1(d7[61]), .CIN(n11519), 
          .COUT(n11520), .S0(d8_71__N_1603[60]), .S1(d8_71__N_1603[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1115_27.INIT0 = 16'hb874;
    defparam add_1115_27.INIT1 = 16'hb874;
    defparam add_1115_27.INJECT1_0 = "NO";
    defparam add_1115_27.INJECT1_1 = "NO";
    CCU2D add_1115_25 (.A0(d_d7[58]), .B0(n6404), .C0(n6405[22]), .D0(d7[58]), 
          .A1(d_d7[59]), .B1(n6404), .C1(n6405[23]), .D1(d7[59]), .CIN(n11518), 
          .COUT(n11519), .S0(d8_71__N_1603[58]), .S1(d8_71__N_1603[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1115_25.INIT0 = 16'hb874;
    defparam add_1115_25.INIT1 = 16'hb874;
    defparam add_1115_25.INJECT1_0 = "NO";
    defparam add_1115_25.INJECT1_1 = "NO";
    CCU2D add_1115_23 (.A0(d_d7[56]), .B0(n6404), .C0(n6405[20]), .D0(d7[56]), 
          .A1(d_d7[57]), .B1(n6404), .C1(n6405[21]), .D1(d7[57]), .CIN(n11517), 
          .COUT(n11518), .S0(d8_71__N_1603[56]), .S1(d8_71__N_1603[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1115_23.INIT0 = 16'hb874;
    defparam add_1115_23.INIT1 = 16'hb874;
    defparam add_1115_23.INJECT1_0 = "NO";
    defparam add_1115_23.INJECT1_1 = "NO";
    CCU2D add_1115_21 (.A0(d_d7[54]), .B0(n6404), .C0(n6405[18]), .D0(d7[54]), 
          .A1(d_d7[55]), .B1(n6404), .C1(n6405[19]), .D1(d7[55]), .CIN(n11516), 
          .COUT(n11517), .S0(d8_71__N_1603[54]), .S1(d8_71__N_1603[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1115_21.INIT0 = 16'hb874;
    defparam add_1115_21.INIT1 = 16'hb874;
    defparam add_1115_21.INJECT1_0 = "NO";
    defparam add_1115_21.INJECT1_1 = "NO";
    CCU2D add_1115_19 (.A0(d_d7[52]), .B0(n6404), .C0(n6405[16]), .D0(d7[52]), 
          .A1(d_d7[53]), .B1(n6404), .C1(n6405[17]), .D1(d7[53]), .CIN(n11515), 
          .COUT(n11516), .S0(d8_71__N_1603[52]), .S1(d8_71__N_1603[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1115_19.INIT0 = 16'hb874;
    defparam add_1115_19.INIT1 = 16'hb874;
    defparam add_1115_19.INJECT1_0 = "NO";
    defparam add_1115_19.INJECT1_1 = "NO";
    CCU2D add_1115_17 (.A0(d_d7[50]), .B0(n6404), .C0(n6405[14]), .D0(d7[50]), 
          .A1(d_d7[51]), .B1(n6404), .C1(n6405[15]), .D1(d7[51]), .CIN(n11514), 
          .COUT(n11515), .S0(d8_71__N_1603[50]), .S1(d8_71__N_1603[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1115_17.INIT0 = 16'hb874;
    defparam add_1115_17.INIT1 = 16'hb874;
    defparam add_1115_17.INJECT1_0 = "NO";
    defparam add_1115_17.INJECT1_1 = "NO";
    CCU2D add_1115_15 (.A0(d_d7[48]), .B0(n6404), .C0(n6405[12]), .D0(d7[48]), 
          .A1(d_d7[49]), .B1(n6404), .C1(n6405[13]), .D1(d7[49]), .CIN(n11513), 
          .COUT(n11514), .S0(d8_71__N_1603[48]), .S1(d8_71__N_1603[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1115_15.INIT0 = 16'hb874;
    defparam add_1115_15.INIT1 = 16'hb874;
    defparam add_1115_15.INJECT1_0 = "NO";
    defparam add_1115_15.INJECT1_1 = "NO";
    CCU2D add_1115_13 (.A0(d_d7[46]), .B0(n6404), .C0(n6405[10]), .D0(d7[46]), 
          .A1(d_d7[47]), .B1(n6404), .C1(n6405[11]), .D1(d7[47]), .CIN(n11512), 
          .COUT(n11513), .S0(d8_71__N_1603[46]), .S1(d8_71__N_1603[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1115_13.INIT0 = 16'hb874;
    defparam add_1115_13.INIT1 = 16'hb874;
    defparam add_1115_13.INJECT1_0 = "NO";
    defparam add_1115_13.INJECT1_1 = "NO";
    CCU2D add_1115_11 (.A0(d_d7[44]), .B0(n6404), .C0(n6405[8]), .D0(d7[44]), 
          .A1(d_d7[45]), .B1(n6404), .C1(n6405[9]), .D1(d7[45]), .CIN(n11511), 
          .COUT(n11512), .S0(d8_71__N_1603[44]), .S1(d8_71__N_1603[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1115_11.INIT0 = 16'hb874;
    defparam add_1115_11.INIT1 = 16'hb874;
    defparam add_1115_11.INJECT1_0 = "NO";
    defparam add_1115_11.INJECT1_1 = "NO";
    CCU2D add_1115_9 (.A0(d_d7[42]), .B0(n6404), .C0(n6405[6]), .D0(d7[42]), 
          .A1(d_d7[43]), .B1(n6404), .C1(n6405[7]), .D1(d7[43]), .CIN(n11510), 
          .COUT(n11511), .S0(d8_71__N_1603[42]), .S1(d8_71__N_1603[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1115_9.INIT0 = 16'hb874;
    defparam add_1115_9.INIT1 = 16'hb874;
    defparam add_1115_9.INJECT1_0 = "NO";
    defparam add_1115_9.INJECT1_1 = "NO";
    CCU2D add_1115_7 (.A0(d_d7[40]), .B0(n6404), .C0(n6405[4]), .D0(d7[40]), 
          .A1(d_d7[41]), .B1(n6404), .C1(n6405[5]), .D1(d7[41]), .CIN(n11509), 
          .COUT(n11510), .S0(d8_71__N_1603[40]), .S1(d8_71__N_1603[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1115_7.INIT0 = 16'hb874;
    defparam add_1115_7.INIT1 = 16'hb874;
    defparam add_1115_7.INJECT1_0 = "NO";
    defparam add_1115_7.INJECT1_1 = "NO";
    CCU2D add_1115_5 (.A0(d_d7[38]), .B0(n6404), .C0(n6405[2]), .D0(d7[38]), 
          .A1(d_d7[39]), .B1(n6404), .C1(n6405[3]), .D1(d7[39]), .CIN(n11508), 
          .COUT(n11509), .S0(d8_71__N_1603[38]), .S1(d8_71__N_1603[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1115_5.INIT0 = 16'hb874;
    defparam add_1115_5.INIT1 = 16'hb874;
    defparam add_1115_5.INJECT1_0 = "NO";
    defparam add_1115_5.INJECT1_1 = "NO";
    CCU2D add_1115_3 (.A0(d_d7[36]), .B0(n6404), .C0(n6405[0]), .D0(d7[36]), 
          .A1(d_d7[37]), .B1(n6404), .C1(n6405[1]), .D1(d7[37]), .CIN(n11507), 
          .COUT(n11508), .S0(d8_71__N_1603[36]), .S1(d8_71__N_1603[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1115_3.INIT0 = 16'hb874;
    defparam add_1115_3.INIT1 = 16'hb874;
    defparam add_1115_3.INJECT1_0 = "NO";
    defparam add_1115_3.INJECT1_1 = "NO";
    CCU2D add_1115_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n6404), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11507));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1115_1.INIT0 = 16'hF000;
    defparam add_1115_1.INIT1 = 16'h0555;
    defparam add_1115_1.INJECT1_0 = "NO";
    defparam add_1115_1.INJECT1_1 = "NO";
    CCU2D add_1119_37 (.A0(d8[71]), .B0(d_d8[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11503), 
          .S0(n6557[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1119_37.INIT0 = 16'h5999;
    defparam add_1119_37.INIT1 = 16'h0000;
    defparam add_1119_37.INJECT1_0 = "NO";
    defparam add_1119_37.INJECT1_1 = "NO";
    CCU2D add_1119_35 (.A0(d8[69]), .B0(d_d8[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[70]), .B1(d_d8[70]), .C1(GND_net), .D1(GND_net), .CIN(n11502), 
          .COUT(n11503), .S0(n6557[33]), .S1(n6557[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1119_35.INIT0 = 16'h5999;
    defparam add_1119_35.INIT1 = 16'h5999;
    defparam add_1119_35.INJECT1_0 = "NO";
    defparam add_1119_35.INJECT1_1 = "NO";
    CCU2D add_1119_33 (.A0(d8[67]), .B0(d_d8[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[68]), .B1(d_d8[68]), .C1(GND_net), .D1(GND_net), .CIN(n11501), 
          .COUT(n11502), .S0(n6557[31]), .S1(n6557[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1119_33.INIT0 = 16'h5999;
    defparam add_1119_33.INIT1 = 16'h5999;
    defparam add_1119_33.INJECT1_0 = "NO";
    defparam add_1119_33.INJECT1_1 = "NO";
    CCU2D add_1119_31 (.A0(d8[65]), .B0(d_d8[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[66]), .B1(d_d8[66]), .C1(GND_net), .D1(GND_net), .CIN(n11500), 
          .COUT(n11501), .S0(n6557[29]), .S1(n6557[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1119_31.INIT0 = 16'h5999;
    defparam add_1119_31.INIT1 = 16'h5999;
    defparam add_1119_31.INJECT1_0 = "NO";
    defparam add_1119_31.INJECT1_1 = "NO";
    CCU2D add_1119_29 (.A0(d8[63]), .B0(d_d8[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[64]), .B1(d_d8[64]), .C1(GND_net), .D1(GND_net), .CIN(n11499), 
          .COUT(n11500), .S0(n6557[27]), .S1(n6557[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1119_29.INIT0 = 16'h5999;
    defparam add_1119_29.INIT1 = 16'h5999;
    defparam add_1119_29.INJECT1_0 = "NO";
    defparam add_1119_29.INJECT1_1 = "NO";
    CCU2D add_1119_27 (.A0(d8[61]), .B0(d_d8[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[62]), .B1(d_d8[62]), .C1(GND_net), .D1(GND_net), .CIN(n11498), 
          .COUT(n11499), .S0(n6557[25]), .S1(n6557[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1119_27.INIT0 = 16'h5999;
    defparam add_1119_27.INIT1 = 16'h5999;
    defparam add_1119_27.INJECT1_0 = "NO";
    defparam add_1119_27.INJECT1_1 = "NO";
    CCU2D add_1119_25 (.A0(d8[59]), .B0(d_d8[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[60]), .B1(d_d8[60]), .C1(GND_net), .D1(GND_net), .CIN(n11497), 
          .COUT(n11498), .S0(n6557[23]), .S1(n6557[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1119_25.INIT0 = 16'h5999;
    defparam add_1119_25.INIT1 = 16'h5999;
    defparam add_1119_25.INJECT1_0 = "NO";
    defparam add_1119_25.INJECT1_1 = "NO";
    CCU2D add_1119_23 (.A0(d8[57]), .B0(d_d8[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[58]), .B1(d_d8[58]), .C1(GND_net), .D1(GND_net), .CIN(n11496), 
          .COUT(n11497), .S0(n6557[21]), .S1(n6557[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1119_23.INIT0 = 16'h5999;
    defparam add_1119_23.INIT1 = 16'h5999;
    defparam add_1119_23.INJECT1_0 = "NO";
    defparam add_1119_23.INJECT1_1 = "NO";
    CCU2D add_1119_21 (.A0(d8[55]), .B0(d_d8[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[56]), .B1(d_d8[56]), .C1(GND_net), .D1(GND_net), .CIN(n11495), 
          .COUT(n11496), .S0(n6557[19]), .S1(n6557[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1119_21.INIT0 = 16'h5999;
    defparam add_1119_21.INIT1 = 16'h5999;
    defparam add_1119_21.INJECT1_0 = "NO";
    defparam add_1119_21.INJECT1_1 = "NO";
    CCU2D add_1119_19 (.A0(d8[53]), .B0(d_d8[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[54]), .B1(d_d8[54]), .C1(GND_net), .D1(GND_net), .CIN(n11494), 
          .COUT(n11495), .S0(n6557[17]), .S1(n6557[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1119_19.INIT0 = 16'h5999;
    defparam add_1119_19.INIT1 = 16'h5999;
    defparam add_1119_19.INJECT1_0 = "NO";
    defparam add_1119_19.INJECT1_1 = "NO";
    CCU2D add_1119_17 (.A0(d8[51]), .B0(d_d8[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[52]), .B1(d_d8[52]), .C1(GND_net), .D1(GND_net), .CIN(n11493), 
          .COUT(n11494), .S0(n6557[15]), .S1(n6557[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1119_17.INIT0 = 16'h5999;
    defparam add_1119_17.INIT1 = 16'h5999;
    defparam add_1119_17.INJECT1_0 = "NO";
    defparam add_1119_17.INJECT1_1 = "NO";
    CCU2D add_1119_15 (.A0(d8[49]), .B0(d_d8[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[50]), .B1(d_d8[50]), .C1(GND_net), .D1(GND_net), .CIN(n11492), 
          .COUT(n11493), .S0(n6557[13]), .S1(n6557[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1119_15.INIT0 = 16'h5999;
    defparam add_1119_15.INIT1 = 16'h5999;
    defparam add_1119_15.INJECT1_0 = "NO";
    defparam add_1119_15.INJECT1_1 = "NO";
    CCU2D add_1119_13 (.A0(d8[47]), .B0(d_d8[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[48]), .B1(d_d8[48]), .C1(GND_net), .D1(GND_net), .CIN(n11491), 
          .COUT(n11492), .S0(n6557[11]), .S1(n6557[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1119_13.INIT0 = 16'h5999;
    defparam add_1119_13.INIT1 = 16'h5999;
    defparam add_1119_13.INJECT1_0 = "NO";
    defparam add_1119_13.INJECT1_1 = "NO";
    CCU2D add_1119_11 (.A0(d8[45]), .B0(d_d8[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[46]), .B1(d_d8[46]), .C1(GND_net), .D1(GND_net), .CIN(n11490), 
          .COUT(n11491), .S0(n6557[9]), .S1(n6557[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1119_11.INIT0 = 16'h5999;
    defparam add_1119_11.INIT1 = 16'h5999;
    defparam add_1119_11.INJECT1_0 = "NO";
    defparam add_1119_11.INJECT1_1 = "NO";
    CCU2D add_1119_9 (.A0(d8[43]), .B0(d_d8[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[44]), .B1(d_d8[44]), .C1(GND_net), .D1(GND_net), .CIN(n11489), 
          .COUT(n11490), .S0(n6557[7]), .S1(n6557[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1119_9.INIT0 = 16'h5999;
    defparam add_1119_9.INIT1 = 16'h5999;
    defparam add_1119_9.INJECT1_0 = "NO";
    defparam add_1119_9.INJECT1_1 = "NO";
    CCU2D add_1119_7 (.A0(d8[41]), .B0(d_d8[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[42]), .B1(d_d8[42]), .C1(GND_net), .D1(GND_net), .CIN(n11488), 
          .COUT(n11489), .S0(n6557[5]), .S1(n6557[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1119_7.INIT0 = 16'h5999;
    defparam add_1119_7.INIT1 = 16'h5999;
    defparam add_1119_7.INJECT1_0 = "NO";
    defparam add_1119_7.INJECT1_1 = "NO";
    CCU2D add_1119_5 (.A0(d8[39]), .B0(d_d8[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[40]), .B1(d_d8[40]), .C1(GND_net), .D1(GND_net), .CIN(n11487), 
          .COUT(n11488), .S0(n6557[3]), .S1(n6557[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1119_5.INIT0 = 16'h5999;
    defparam add_1119_5.INIT1 = 16'h5999;
    defparam add_1119_5.INJECT1_0 = "NO";
    defparam add_1119_5.INJECT1_1 = "NO";
    CCU2D add_1119_3 (.A0(d8[37]), .B0(d_d8[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[38]), .B1(d_d8[38]), .C1(GND_net), .D1(GND_net), .CIN(n11486), 
          .COUT(n11487), .S0(n6557[1]), .S1(n6557[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1119_3.INIT0 = 16'h5999;
    defparam add_1119_3.INIT1 = 16'h5999;
    defparam add_1119_3.INJECT1_0 = "NO";
    defparam add_1119_3.INJECT1_1 = "NO";
    CCU2D add_1119_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d8[36]), .B1(d_d8[36]), .C1(GND_net), .D1(GND_net), .COUT(n11486), 
          .S1(n6557[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1119_1.INIT0 = 16'hF000;
    defparam add_1119_1.INIT1 = 16'h5999;
    defparam add_1119_1.INJECT1_0 = "NO";
    defparam add_1119_1.INJECT1_1 = "NO";
    CCU2D add_1120_37 (.A0(d_d8[70]), .B0(n6556), .C0(n6557[34]), .D0(d8[70]), 
          .A1(d_d8[71]), .B1(n6556), .C1(n6557[35]), .D1(d8[71]), .CIN(n11484), 
          .S0(d9_71__N_1675[70]), .S1(d9_71__N_1675[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1120_37.INIT0 = 16'hb874;
    defparam add_1120_37.INIT1 = 16'hb874;
    defparam add_1120_37.INJECT1_0 = "NO";
    defparam add_1120_37.INJECT1_1 = "NO";
    CCU2D add_1120_35 (.A0(d_d8[68]), .B0(n6556), .C0(n6557[32]), .D0(d8[68]), 
          .A1(d_d8[69]), .B1(n6556), .C1(n6557[33]), .D1(d8[69]), .CIN(n11483), 
          .COUT(n11484), .S0(d9_71__N_1675[68]), .S1(d9_71__N_1675[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1120_35.INIT0 = 16'hb874;
    defparam add_1120_35.INIT1 = 16'hb874;
    defparam add_1120_35.INJECT1_0 = "NO";
    defparam add_1120_35.INJECT1_1 = "NO";
    CCU2D add_1120_33 (.A0(d_d8[66]), .B0(n6556), .C0(n6557[30]), .D0(d8[66]), 
          .A1(d_d8[67]), .B1(n6556), .C1(n6557[31]), .D1(d8[67]), .CIN(n11482), 
          .COUT(n11483), .S0(d9_71__N_1675[66]), .S1(d9_71__N_1675[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1120_33.INIT0 = 16'hb874;
    defparam add_1120_33.INIT1 = 16'hb874;
    defparam add_1120_33.INJECT1_0 = "NO";
    defparam add_1120_33.INJECT1_1 = "NO";
    CCU2D add_1120_31 (.A0(d_d8[64]), .B0(n6556), .C0(n6557[28]), .D0(d8[64]), 
          .A1(d_d8[65]), .B1(n6556), .C1(n6557[29]), .D1(d8[65]), .CIN(n11481), 
          .COUT(n11482), .S0(d9_71__N_1675[64]), .S1(d9_71__N_1675[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1120_31.INIT0 = 16'hb874;
    defparam add_1120_31.INIT1 = 16'hb874;
    defparam add_1120_31.INJECT1_0 = "NO";
    defparam add_1120_31.INJECT1_1 = "NO";
    CCU2D add_1120_29 (.A0(d_d8[62]), .B0(n6556), .C0(n6557[26]), .D0(d8[62]), 
          .A1(d_d8[63]), .B1(n6556), .C1(n6557[27]), .D1(d8[63]), .CIN(n11480), 
          .COUT(n11481), .S0(d9_71__N_1675[62]), .S1(d9_71__N_1675[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1120_29.INIT0 = 16'hb874;
    defparam add_1120_29.INIT1 = 16'hb874;
    defparam add_1120_29.INJECT1_0 = "NO";
    defparam add_1120_29.INJECT1_1 = "NO";
    CCU2D add_1120_27 (.A0(d_d8[60]), .B0(n6556), .C0(n6557[24]), .D0(d8[60]), 
          .A1(d_d8[61]), .B1(n6556), .C1(n6557[25]), .D1(d8[61]), .CIN(n11479), 
          .COUT(n11480), .S0(d9_71__N_1675[60]), .S1(d9_71__N_1675[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1120_27.INIT0 = 16'hb874;
    defparam add_1120_27.INIT1 = 16'hb874;
    defparam add_1120_27.INJECT1_0 = "NO";
    defparam add_1120_27.INJECT1_1 = "NO";
    CCU2D add_1120_25 (.A0(d_d8[58]), .B0(n6556), .C0(n6557[22]), .D0(d8[58]), 
          .A1(d_d8[59]), .B1(n6556), .C1(n6557[23]), .D1(d8[59]), .CIN(n11478), 
          .COUT(n11479), .S0(d9_71__N_1675[58]), .S1(d9_71__N_1675[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1120_25.INIT0 = 16'hb874;
    defparam add_1120_25.INIT1 = 16'hb874;
    defparam add_1120_25.INJECT1_0 = "NO";
    defparam add_1120_25.INJECT1_1 = "NO";
    CCU2D add_1120_23 (.A0(d_d8[56]), .B0(n6556), .C0(n6557[20]), .D0(d8[56]), 
          .A1(d_d8[57]), .B1(n6556), .C1(n6557[21]), .D1(d8[57]), .CIN(n11477), 
          .COUT(n11478), .S0(d9_71__N_1675[56]), .S1(d9_71__N_1675[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1120_23.INIT0 = 16'hb874;
    defparam add_1120_23.INIT1 = 16'hb874;
    defparam add_1120_23.INJECT1_0 = "NO";
    defparam add_1120_23.INJECT1_1 = "NO";
    CCU2D add_1120_21 (.A0(d_d8[54]), .B0(n6556), .C0(n6557[18]), .D0(d8[54]), 
          .A1(d_d8[55]), .B1(n6556), .C1(n6557[19]), .D1(d8[55]), .CIN(n11476), 
          .COUT(n11477), .S0(d9_71__N_1675[54]), .S1(d9_71__N_1675[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1120_21.INIT0 = 16'hb874;
    defparam add_1120_21.INIT1 = 16'hb874;
    defparam add_1120_21.INJECT1_0 = "NO";
    defparam add_1120_21.INJECT1_1 = "NO";
    CCU2D add_1120_19 (.A0(d_d8[52]), .B0(n6556), .C0(n6557[16]), .D0(d8[52]), 
          .A1(d_d8[53]), .B1(n6556), .C1(n6557[17]), .D1(d8[53]), .CIN(n11475), 
          .COUT(n11476), .S0(d9_71__N_1675[52]), .S1(d9_71__N_1675[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1120_19.INIT0 = 16'hb874;
    defparam add_1120_19.INIT1 = 16'hb874;
    defparam add_1120_19.INJECT1_0 = "NO";
    defparam add_1120_19.INJECT1_1 = "NO";
    CCU2D add_1120_17 (.A0(d_d8[50]), .B0(n6556), .C0(n6557[14]), .D0(d8[50]), 
          .A1(d_d8[51]), .B1(n6556), .C1(n6557[15]), .D1(d8[51]), .CIN(n11474), 
          .COUT(n11475), .S0(d9_71__N_1675[50]), .S1(d9_71__N_1675[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1120_17.INIT0 = 16'hb874;
    defparam add_1120_17.INIT1 = 16'hb874;
    defparam add_1120_17.INJECT1_0 = "NO";
    defparam add_1120_17.INJECT1_1 = "NO";
    CCU2D add_1120_15 (.A0(d_d8[48]), .B0(n6556), .C0(n6557[12]), .D0(d8[48]), 
          .A1(d_d8[49]), .B1(n6556), .C1(n6557[13]), .D1(d8[49]), .CIN(n11473), 
          .COUT(n11474), .S0(d9_71__N_1675[48]), .S1(d9_71__N_1675[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1120_15.INIT0 = 16'hb874;
    defparam add_1120_15.INIT1 = 16'hb874;
    defparam add_1120_15.INJECT1_0 = "NO";
    defparam add_1120_15.INJECT1_1 = "NO";
    CCU2D add_1120_13 (.A0(d_d8[46]), .B0(n6556), .C0(n6557[10]), .D0(d8[46]), 
          .A1(d_d8[47]), .B1(n6556), .C1(n6557[11]), .D1(d8[47]), .CIN(n11472), 
          .COUT(n11473), .S0(d9_71__N_1675[46]), .S1(d9_71__N_1675[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1120_13.INIT0 = 16'hb874;
    defparam add_1120_13.INIT1 = 16'hb874;
    defparam add_1120_13.INJECT1_0 = "NO";
    defparam add_1120_13.INJECT1_1 = "NO";
    CCU2D add_1120_11 (.A0(d_d8[44]), .B0(n6556), .C0(n6557[8]), .D0(d8[44]), 
          .A1(d_d8[45]), .B1(n6556), .C1(n6557[9]), .D1(d8[45]), .CIN(n11471), 
          .COUT(n11472), .S0(d9_71__N_1675[44]), .S1(d9_71__N_1675[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1120_11.INIT0 = 16'hb874;
    defparam add_1120_11.INIT1 = 16'hb874;
    defparam add_1120_11.INJECT1_0 = "NO";
    defparam add_1120_11.INJECT1_1 = "NO";
    CCU2D add_1120_9 (.A0(d_d8[42]), .B0(n6556), .C0(n6557[6]), .D0(d8[42]), 
          .A1(d_d8[43]), .B1(n6556), .C1(n6557[7]), .D1(d8[43]), .CIN(n11470), 
          .COUT(n11471), .S0(d9_71__N_1675[42]), .S1(d9_71__N_1675[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1120_9.INIT0 = 16'hb874;
    defparam add_1120_9.INIT1 = 16'hb874;
    defparam add_1120_9.INJECT1_0 = "NO";
    defparam add_1120_9.INJECT1_1 = "NO";
    CCU2D add_1120_7 (.A0(d_d8[40]), .B0(n6556), .C0(n6557[4]), .D0(d8[40]), 
          .A1(d_d8[41]), .B1(n6556), .C1(n6557[5]), .D1(d8[41]), .CIN(n11469), 
          .COUT(n11470), .S0(d9_71__N_1675[40]), .S1(d9_71__N_1675[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1120_7.INIT0 = 16'hb874;
    defparam add_1120_7.INIT1 = 16'hb874;
    defparam add_1120_7.INJECT1_0 = "NO";
    defparam add_1120_7.INJECT1_1 = "NO";
    CCU2D add_1120_5 (.A0(d_d8[38]), .B0(n6556), .C0(n6557[2]), .D0(d8[38]), 
          .A1(d_d8[39]), .B1(n6556), .C1(n6557[3]), .D1(d8[39]), .CIN(n11468), 
          .COUT(n11469), .S0(d9_71__N_1675[38]), .S1(d9_71__N_1675[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1120_5.INIT0 = 16'hb874;
    defparam add_1120_5.INIT1 = 16'hb874;
    defparam add_1120_5.INJECT1_0 = "NO";
    defparam add_1120_5.INJECT1_1 = "NO";
    CCU2D add_1120_3 (.A0(d_d8[36]), .B0(n6556), .C0(n6557[0]), .D0(d8[36]), 
          .A1(d_d8[37]), .B1(n6556), .C1(n6557[1]), .D1(d8[37]), .CIN(n11467), 
          .COUT(n11468), .S0(d9_71__N_1675[36]), .S1(d9_71__N_1675[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1120_3.INIT0 = 16'hb874;
    defparam add_1120_3.INIT1 = 16'hb874;
    defparam add_1120_3.INJECT1_0 = "NO";
    defparam add_1120_3.INJECT1_1 = "NO";
    CCU2D add_1120_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n6556), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11467));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1120_1.INIT0 = 16'hF000;
    defparam add_1120_1.INIT1 = 16'h0555;
    defparam add_1120_1.INJECT1_0 = "NO";
    defparam add_1120_1.INJECT1_1 = "NO";
    CCU2D add_1124_37 (.A0(d9[71]), .B0(d_d9[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11463), 
          .S0(n6709[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1124_37.INIT0 = 16'h5999;
    defparam add_1124_37.INIT1 = 16'h0000;
    defparam add_1124_37.INJECT1_0 = "NO";
    defparam add_1124_37.INJECT1_1 = "NO";
    CCU2D add_1124_35 (.A0(d9[69]), .B0(d_d9[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[70]), .B1(d_d9[70]), .C1(GND_net), .D1(GND_net), .CIN(n11462), 
          .COUT(n11463), .S0(n6709[33]), .S1(n6709[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1124_35.INIT0 = 16'h5999;
    defparam add_1124_35.INIT1 = 16'h5999;
    defparam add_1124_35.INJECT1_0 = "NO";
    defparam add_1124_35.INJECT1_1 = "NO";
    CCU2D add_1124_33 (.A0(d9[67]), .B0(d_d9[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[68]), .B1(d_d9[68]), .C1(GND_net), .D1(GND_net), .CIN(n11461), 
          .COUT(n11462), .S0(n6709[31]), .S1(n6709[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1124_33.INIT0 = 16'h5999;
    defparam add_1124_33.INIT1 = 16'h5999;
    defparam add_1124_33.INJECT1_0 = "NO";
    defparam add_1124_33.INJECT1_1 = "NO";
    CCU2D add_1124_31 (.A0(d9[65]), .B0(d_d9[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[66]), .B1(d_d9[66]), .C1(GND_net), .D1(GND_net), .CIN(n11460), 
          .COUT(n11461), .S0(n6709[29]), .S1(n6709[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1124_31.INIT0 = 16'h5999;
    defparam add_1124_31.INIT1 = 16'h5999;
    defparam add_1124_31.INJECT1_0 = "NO";
    defparam add_1124_31.INJECT1_1 = "NO";
    CCU2D add_1124_29 (.A0(d9[63]), .B0(d_d9[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[64]), .B1(d_d9[64]), .C1(GND_net), .D1(GND_net), .CIN(n11459), 
          .COUT(n11460), .S0(n6709[27]), .S1(n6709[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1124_29.INIT0 = 16'h5999;
    defparam add_1124_29.INIT1 = 16'h5999;
    defparam add_1124_29.INJECT1_0 = "NO";
    defparam add_1124_29.INJECT1_1 = "NO";
    CCU2D add_1124_27 (.A0(d9[61]), .B0(d_d9[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[62]), .B1(d_d9[62]), .C1(GND_net), .D1(GND_net), .CIN(n11458), 
          .COUT(n11459), .S0(n6709[25]), .S1(n6709[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1124_27.INIT0 = 16'h5999;
    defparam add_1124_27.INIT1 = 16'h5999;
    defparam add_1124_27.INJECT1_0 = "NO";
    defparam add_1124_27.INJECT1_1 = "NO";
    CCU2D add_1124_25 (.A0(d9[59]), .B0(d_d9[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[60]), .B1(d_d9[60]), .C1(GND_net), .D1(GND_net), .CIN(n11457), 
          .COUT(n11458), .S0(n6709[23]), .S1(n6709[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1124_25.INIT0 = 16'h5999;
    defparam add_1124_25.INIT1 = 16'h5999;
    defparam add_1124_25.INJECT1_0 = "NO";
    defparam add_1124_25.INJECT1_1 = "NO";
    CCU2D add_1124_23 (.A0(d9[57]), .B0(d_d9[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[58]), .B1(d_d9[58]), .C1(GND_net), .D1(GND_net), .CIN(n11456), 
          .COUT(n11457), .S0(n6709[21]), .S1(n6709[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1124_23.INIT0 = 16'h5999;
    defparam add_1124_23.INIT1 = 16'h5999;
    defparam add_1124_23.INJECT1_0 = "NO";
    defparam add_1124_23.INJECT1_1 = "NO";
    CCU2D add_1124_21 (.A0(d9[55]), .B0(d_d9[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[56]), .B1(d_d9[56]), .C1(GND_net), .D1(GND_net), .CIN(n11455), 
          .COUT(n11456));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1124_21.INIT0 = 16'h5999;
    defparam add_1124_21.INIT1 = 16'h5999;
    defparam add_1124_21.INJECT1_0 = "NO";
    defparam add_1124_21.INJECT1_1 = "NO";
    CCU2D add_1124_19 (.A0(d9[53]), .B0(d_d9[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[54]), .B1(d_d9[54]), .C1(GND_net), .D1(GND_net), .CIN(n11454), 
          .COUT(n11455));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1124_19.INIT0 = 16'h5999;
    defparam add_1124_19.INIT1 = 16'h5999;
    defparam add_1124_19.INJECT1_0 = "NO";
    defparam add_1124_19.INJECT1_1 = "NO";
    CCU2D add_1124_17 (.A0(d9[51]), .B0(d_d9[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[52]), .B1(d_d9[52]), .C1(GND_net), .D1(GND_net), .CIN(n11453), 
          .COUT(n11454));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1124_17.INIT0 = 16'h5999;
    defparam add_1124_17.INIT1 = 16'h5999;
    defparam add_1124_17.INJECT1_0 = "NO";
    defparam add_1124_17.INJECT1_1 = "NO";
    CCU2D add_1124_15 (.A0(d9[49]), .B0(d_d9[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[50]), .B1(d_d9[50]), .C1(GND_net), .D1(GND_net), .CIN(n11452), 
          .COUT(n11453));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1124_15.INIT0 = 16'h5999;
    defparam add_1124_15.INIT1 = 16'h5999;
    defparam add_1124_15.INJECT1_0 = "NO";
    defparam add_1124_15.INJECT1_1 = "NO";
    CCU2D add_1124_13 (.A0(d9[47]), .B0(d_d9[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[48]), .B1(d_d9[48]), .C1(GND_net), .D1(GND_net), .CIN(n11451), 
          .COUT(n11452));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1124_13.INIT0 = 16'h5999;
    defparam add_1124_13.INIT1 = 16'h5999;
    defparam add_1124_13.INJECT1_0 = "NO";
    defparam add_1124_13.INJECT1_1 = "NO";
    CCU2D add_1124_11 (.A0(d9[45]), .B0(d_d9[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[46]), .B1(d_d9[46]), .C1(GND_net), .D1(GND_net), .CIN(n11450), 
          .COUT(n11451));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1124_11.INIT0 = 16'h5999;
    defparam add_1124_11.INIT1 = 16'h5999;
    defparam add_1124_11.INJECT1_0 = "NO";
    defparam add_1124_11.INJECT1_1 = "NO";
    CCU2D add_1124_9 (.A0(d9[43]), .B0(d_d9[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[44]), .B1(d_d9[44]), .C1(GND_net), .D1(GND_net), .CIN(n11449), 
          .COUT(n11450));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1124_9.INIT0 = 16'h5999;
    defparam add_1124_9.INIT1 = 16'h5999;
    defparam add_1124_9.INJECT1_0 = "NO";
    defparam add_1124_9.INJECT1_1 = "NO";
    CCU2D add_1124_7 (.A0(d9[41]), .B0(d_d9[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[42]), .B1(d_d9[42]), .C1(GND_net), .D1(GND_net), .CIN(n11448), 
          .COUT(n11449));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1124_7.INIT0 = 16'h5999;
    defparam add_1124_7.INIT1 = 16'h5999;
    defparam add_1124_7.INJECT1_0 = "NO";
    defparam add_1124_7.INJECT1_1 = "NO";
    CCU2D add_1124_5 (.A0(d9[39]), .B0(d_d9[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[40]), .B1(d_d9[40]), .C1(GND_net), .D1(GND_net), .CIN(n11447), 
          .COUT(n11448));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1124_5.INIT0 = 16'h5999;
    defparam add_1124_5.INIT1 = 16'h5999;
    defparam add_1124_5.INJECT1_0 = "NO";
    defparam add_1124_5.INJECT1_1 = "NO";
    CCU2D add_1124_3 (.A0(d9[37]), .B0(d_d9[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[38]), .B1(d_d9[38]), .C1(GND_net), .D1(GND_net), .CIN(n11446), 
          .COUT(n11447));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1124_3.INIT0 = 16'h5999;
    defparam add_1124_3.INIT1 = 16'h5999;
    defparam add_1124_3.INJECT1_0 = "NO";
    defparam add_1124_3.INJECT1_1 = "NO";
    CCU2D add_1124_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d9[36]), .B1(d_d9[36]), .C1(GND_net), .D1(GND_net), .COUT(n11446));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1124_1.INIT0 = 16'hF000;
    defparam add_1124_1.INIT1 = 16'h5999;
    defparam add_1124_1.INJECT1_0 = "NO";
    defparam add_1124_1.INJECT1_1 = "NO";
    CCU2D add_1125_37 (.A0(d9[71]), .B0(d_d9[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11445), 
          .S0(n6747[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1125_37.INIT0 = 16'h5999;
    defparam add_1125_37.INIT1 = 16'h0000;
    defparam add_1125_37.INJECT1_0 = "NO";
    defparam add_1125_37.INJECT1_1 = "NO";
    CCU2D add_1125_35 (.A0(d9[69]), .B0(d_d9[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[70]), .B1(d_d9[70]), .C1(GND_net), .D1(GND_net), .CIN(n11444), 
          .COUT(n11445), .S0(n6747[33]), .S1(n6747[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1125_35.INIT0 = 16'h5999;
    defparam add_1125_35.INIT1 = 16'h5999;
    defparam add_1125_35.INJECT1_0 = "NO";
    defparam add_1125_35.INJECT1_1 = "NO";
    CCU2D add_1125_33 (.A0(d9[67]), .B0(d_d9[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[68]), .B1(d_d9[68]), .C1(GND_net), .D1(GND_net), .CIN(n11443), 
          .COUT(n11444), .S0(n6747[31]), .S1(n6747[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1125_33.INIT0 = 16'h5999;
    defparam add_1125_33.INIT1 = 16'h5999;
    defparam add_1125_33.INJECT1_0 = "NO";
    defparam add_1125_33.INJECT1_1 = "NO";
    CCU2D add_1125_31 (.A0(d9[65]), .B0(d_d9[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[66]), .B1(d_d9[66]), .C1(GND_net), .D1(GND_net), .CIN(n11442), 
          .COUT(n11443), .S0(n6747[29]), .S1(n6747[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1125_31.INIT0 = 16'h5999;
    defparam add_1125_31.INIT1 = 16'h5999;
    defparam add_1125_31.INJECT1_0 = "NO";
    defparam add_1125_31.INJECT1_1 = "NO";
    CCU2D add_1125_29 (.A0(d9[63]), .B0(d_d9[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[64]), .B1(d_d9[64]), .C1(GND_net), .D1(GND_net), .CIN(n11441), 
          .COUT(n11442), .S0(n6747[27]), .S1(n6747[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1125_29.INIT0 = 16'h5999;
    defparam add_1125_29.INIT1 = 16'h5999;
    defparam add_1125_29.INJECT1_0 = "NO";
    defparam add_1125_29.INJECT1_1 = "NO";
    CCU2D add_1125_27 (.A0(d9[61]), .B0(d_d9[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[62]), .B1(d_d9[62]), .C1(GND_net), .D1(GND_net), .CIN(n11440), 
          .COUT(n11441), .S0(n6747[25]), .S1(n6747[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1125_27.INIT0 = 16'h5999;
    defparam add_1125_27.INIT1 = 16'h5999;
    defparam add_1125_27.INJECT1_0 = "NO";
    defparam add_1125_27.INJECT1_1 = "NO";
    CCU2D add_1125_25 (.A0(d9[59]), .B0(d_d9[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[60]), .B1(d_d9[60]), .C1(GND_net), .D1(GND_net), .CIN(n11439), 
          .COUT(n11440), .S0(n6747[23]), .S1(n6747[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1125_25.INIT0 = 16'h5999;
    defparam add_1125_25.INIT1 = 16'h5999;
    defparam add_1125_25.INJECT1_0 = "NO";
    defparam add_1125_25.INJECT1_1 = "NO";
    CCU2D add_1125_23 (.A0(d9[57]), .B0(d_d9[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[58]), .B1(d_d9[58]), .C1(GND_net), .D1(GND_net), .CIN(n11438), 
          .COUT(n11439), .S0(n6747[21]), .S1(n6747[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1125_23.INIT0 = 16'h5999;
    defparam add_1125_23.INIT1 = 16'h5999;
    defparam add_1125_23.INJECT1_0 = "NO";
    defparam add_1125_23.INJECT1_1 = "NO";
    CCU2D add_1125_21 (.A0(d9[55]), .B0(d_d9[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[56]), .B1(d_d9[56]), .C1(GND_net), .D1(GND_net), .CIN(n11437), 
          .COUT(n11438));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1125_21.INIT0 = 16'h5999;
    defparam add_1125_21.INIT1 = 16'h5999;
    defparam add_1125_21.INJECT1_0 = "NO";
    defparam add_1125_21.INJECT1_1 = "NO";
    CCU2D add_1125_19 (.A0(d9[53]), .B0(d_d9[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[54]), .B1(d_d9[54]), .C1(GND_net), .D1(GND_net), .CIN(n11436), 
          .COUT(n11437));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1125_19.INIT0 = 16'h5999;
    defparam add_1125_19.INIT1 = 16'h5999;
    defparam add_1125_19.INJECT1_0 = "NO";
    defparam add_1125_19.INJECT1_1 = "NO";
    CCU2D add_1125_17 (.A0(d9[51]), .B0(d_d9[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[52]), .B1(d_d9[52]), .C1(GND_net), .D1(GND_net), .CIN(n11435), 
          .COUT(n11436));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1125_17.INIT0 = 16'h5999;
    defparam add_1125_17.INIT1 = 16'h5999;
    defparam add_1125_17.INJECT1_0 = "NO";
    defparam add_1125_17.INJECT1_1 = "NO";
    CCU2D add_1125_15 (.A0(d9[49]), .B0(d_d9[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[50]), .B1(d_d9[50]), .C1(GND_net), .D1(GND_net), .CIN(n11434), 
          .COUT(n11435));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1125_15.INIT0 = 16'h5999;
    defparam add_1125_15.INIT1 = 16'h5999;
    defparam add_1125_15.INJECT1_0 = "NO";
    defparam add_1125_15.INJECT1_1 = "NO";
    CCU2D add_1125_13 (.A0(d9[47]), .B0(d_d9[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[48]), .B1(d_d9[48]), .C1(GND_net), .D1(GND_net), .CIN(n11433), 
          .COUT(n11434));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1125_13.INIT0 = 16'h5999;
    defparam add_1125_13.INIT1 = 16'h5999;
    defparam add_1125_13.INJECT1_0 = "NO";
    defparam add_1125_13.INJECT1_1 = "NO";
    CCU2D add_1125_11 (.A0(d9[45]), .B0(d_d9[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[46]), .B1(d_d9[46]), .C1(GND_net), .D1(GND_net), .CIN(n11432), 
          .COUT(n11433));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1125_11.INIT0 = 16'h5999;
    defparam add_1125_11.INIT1 = 16'h5999;
    defparam add_1125_11.INJECT1_0 = "NO";
    defparam add_1125_11.INJECT1_1 = "NO";
    CCU2D add_1125_9 (.A0(d9[43]), .B0(d_d9[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[44]), .B1(d_d9[44]), .C1(GND_net), .D1(GND_net), .CIN(n11431), 
          .COUT(n11432));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1125_9.INIT0 = 16'h5999;
    defparam add_1125_9.INIT1 = 16'h5999;
    defparam add_1125_9.INJECT1_0 = "NO";
    defparam add_1125_9.INJECT1_1 = "NO";
    CCU2D add_1125_7 (.A0(d9[41]), .B0(d_d9[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[42]), .B1(d_d9[42]), .C1(GND_net), .D1(GND_net), .CIN(n11430), 
          .COUT(n11431));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1125_7.INIT0 = 16'h5999;
    defparam add_1125_7.INIT1 = 16'h5999;
    defparam add_1125_7.INJECT1_0 = "NO";
    defparam add_1125_7.INJECT1_1 = "NO";
    CCU2D add_1125_5 (.A0(d9[39]), .B0(d_d9[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[40]), .B1(d_d9[40]), .C1(GND_net), .D1(GND_net), .CIN(n11429), 
          .COUT(n11430));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1125_5.INIT0 = 16'h5999;
    defparam add_1125_5.INIT1 = 16'h5999;
    defparam add_1125_5.INJECT1_0 = "NO";
    defparam add_1125_5.INJECT1_1 = "NO";
    CCU2D add_1125_3 (.A0(d9[37]), .B0(d_d9[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[38]), .B1(d_d9[38]), .C1(GND_net), .D1(GND_net), .CIN(n11428), 
          .COUT(n11429));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1125_3.INIT0 = 16'h5999;
    defparam add_1125_3.INIT1 = 16'h5999;
    defparam add_1125_3.INJECT1_0 = "NO";
    defparam add_1125_3.INJECT1_1 = "NO";
    CCU2D add_1125_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d9[36]), .B1(d_d9[36]), .C1(GND_net), .D1(GND_net), .COUT(n11428));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1125_1.INIT0 = 16'h0000;
    defparam add_1125_1.INIT1 = 16'h5999;
    defparam add_1125_1.INJECT1_0 = "NO";
    defparam add_1125_1.INJECT1_1 = "NO";
    FD1S3IX count__i2 (.D(n375[2]), .CK(osc_clk), .CD(n8387), .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n375[3]), .CK(osc_clk), .CD(n8387), .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n375[4]), .CK(osc_clk), .CD(n8387), .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n375[5]), .CK(osc_clk), .CD(n8387), .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n375[6]), .CK(osc_clk), .CD(n8387), .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n375[7]), .CK(osc_clk), .CD(n8387), .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n375[8]), .CK(osc_clk), .CD(n8387), .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n375[9]), .CK(osc_clk), .CD(n8387), .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n375[10]), .CK(osc_clk), .CD(n8387), .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_15__N_1442[11]), .CK(osc_clk), .CD(count_15__N_1458), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(n375[12]), .CK(osc_clk), .CD(n8387), .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(n375[13]), .CK(osc_clk), .CD(n8387), .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(n375[14]), .CK(osc_clk), .CD(n8387), .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(n375[15]), .CK(osc_clk), .CD(n8387), .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i15.GSR = "ENABLED";
    CCU2D add_10_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11231), 
          .S0(n375[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_17.INIT0 = 16'h5aaa;
    defparam add_10_17.INIT1 = 16'h0000;
    defparam add_10_17.INJECT1_0 = "NO";
    defparam add_10_17.INJECT1_1 = "NO";
    CCU2D add_10_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11230), .COUT(n11231), .S0(n375[13]), .S1(n375[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_15.INIT0 = 16'h5aaa;
    defparam add_10_15.INIT1 = 16'h5aaa;
    defparam add_10_15.INJECT1_0 = "NO";
    defparam add_10_15.INJECT1_1 = "NO";
    CCU2D add_10_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11229), .COUT(n11230), .S0(n375[11]), .S1(n375[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_13.INIT0 = 16'h5aaa;
    defparam add_10_13.INIT1 = 16'h5aaa;
    defparam add_10_13.INJECT1_0 = "NO";
    defparam add_10_13.INJECT1_1 = "NO";
    CCU2D add_10_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11228), .COUT(n11229), .S0(n375[9]), .S1(n375[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_11.INIT0 = 16'h5aaa;
    defparam add_10_11.INIT1 = 16'h5aaa;
    defparam add_10_11.INJECT1_0 = "NO";
    defparam add_10_11.INJECT1_1 = "NO";
    CCU2D add_10_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11227), 
          .COUT(n11228), .S0(n375[7]), .S1(n375[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_9.INIT0 = 16'h5aaa;
    defparam add_10_9.INIT1 = 16'h5aaa;
    defparam add_10_9.INJECT1_0 = "NO";
    defparam add_10_9.INJECT1_1 = "NO";
    CCU2D add_10_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11226), 
          .COUT(n11227), .S0(n375[5]), .S1(n375[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_7.INIT0 = 16'h5aaa;
    defparam add_10_7.INIT1 = 16'h5aaa;
    defparam add_10_7.INJECT1_0 = "NO";
    defparam add_10_7.INJECT1_1 = "NO";
    CCU2D add_10_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11225), 
          .COUT(n11226), .S0(n375[3]), .S1(n375[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_5.INIT0 = 16'h5aaa;
    defparam add_10_5.INIT1 = 16'h5aaa;
    defparam add_10_5.INJECT1_0 = "NO";
    defparam add_10_5.INJECT1_1 = "NO";
    CCU2D add_10_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11224), 
          .COUT(n11225), .S0(n375[1]), .S1(n375[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_3.INIT0 = 16'h5aaa;
    defparam add_10_3.INIT1 = 16'h5aaa;
    defparam add_10_3.INJECT1_0 = "NO";
    defparam add_10_3.INJECT1_1 = "NO";
    CCU2D add_10_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11224), 
          .S1(n375[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_1.INIT0 = 16'hF000;
    defparam add_10_1.INIT1 = 16'h5555;
    defparam add_10_1.INJECT1_0 = "NO";
    defparam add_10_1.INJECT1_1 = "NO";
    CCU2D add_1088_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11205), 
          .S0(n5644));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1088_cout.INIT0 = 16'h0000;
    defparam add_1088_cout.INIT1 = 16'h0000;
    defparam add_1088_cout.INJECT1_0 = "NO";
    defparam add_1088_cout.INJECT1_1 = "NO";
    CCU2D add_1088_36 (.A0(d4[34]), .B0(d5[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[35]), .B1(d5[35]), .C1(GND_net), .D1(GND_net), .CIN(n11204), 
          .COUT(n11205), .S0(d5_71__N_706[34]), .S1(d5_71__N_706[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1088_36.INIT0 = 16'h5666;
    defparam add_1088_36.INIT1 = 16'h5666;
    defparam add_1088_36.INJECT1_0 = "NO";
    defparam add_1088_36.INJECT1_1 = "NO";
    CCU2D add_1088_34 (.A0(d4[32]), .B0(d5[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[33]), .B1(d5[33]), .C1(GND_net), .D1(GND_net), .CIN(n11203), 
          .COUT(n11204), .S0(d5_71__N_706[32]), .S1(d5_71__N_706[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1088_34.INIT0 = 16'h5666;
    defparam add_1088_34.INIT1 = 16'h5666;
    defparam add_1088_34.INJECT1_0 = "NO";
    defparam add_1088_34.INJECT1_1 = "NO";
    CCU2D add_1088_32 (.A0(d4[30]), .B0(d5[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[31]), .B1(d5[31]), .C1(GND_net), .D1(GND_net), .CIN(n11202), 
          .COUT(n11203), .S0(d5_71__N_706[30]), .S1(d5_71__N_706[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1088_32.INIT0 = 16'h5666;
    defparam add_1088_32.INIT1 = 16'h5666;
    defparam add_1088_32.INJECT1_0 = "NO";
    defparam add_1088_32.INJECT1_1 = "NO";
    CCU2D add_1088_30 (.A0(d4[28]), .B0(d5[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[29]), .B1(d5[29]), .C1(GND_net), .D1(GND_net), .CIN(n11201), 
          .COUT(n11202), .S0(d5_71__N_706[28]), .S1(d5_71__N_706[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1088_30.INIT0 = 16'h5666;
    defparam add_1088_30.INIT1 = 16'h5666;
    defparam add_1088_30.INJECT1_0 = "NO";
    defparam add_1088_30.INJECT1_1 = "NO";
    CCU2D add_1088_28 (.A0(d4[26]), .B0(d5[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[27]), .B1(d5[27]), .C1(GND_net), .D1(GND_net), .CIN(n11200), 
          .COUT(n11201), .S0(d5_71__N_706[26]), .S1(d5_71__N_706[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1088_28.INIT0 = 16'h5666;
    defparam add_1088_28.INIT1 = 16'h5666;
    defparam add_1088_28.INJECT1_0 = "NO";
    defparam add_1088_28.INJECT1_1 = "NO";
    CCU2D add_1088_26 (.A0(d4[24]), .B0(d5[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[25]), .B1(d5[25]), .C1(GND_net), .D1(GND_net), .CIN(n11199), 
          .COUT(n11200), .S0(d5_71__N_706[24]), .S1(d5_71__N_706[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1088_26.INIT0 = 16'h5666;
    defparam add_1088_26.INIT1 = 16'h5666;
    defparam add_1088_26.INJECT1_0 = "NO";
    defparam add_1088_26.INJECT1_1 = "NO";
    CCU2D add_1088_24 (.A0(d4[22]), .B0(d5[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[23]), .B1(d5[23]), .C1(GND_net), .D1(GND_net), .CIN(n11198), 
          .COUT(n11199), .S0(d5_71__N_706[22]), .S1(d5_71__N_706[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1088_24.INIT0 = 16'h5666;
    defparam add_1088_24.INIT1 = 16'h5666;
    defparam add_1088_24.INJECT1_0 = "NO";
    defparam add_1088_24.INJECT1_1 = "NO";
    CCU2D add_1088_22 (.A0(d4[20]), .B0(d5[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[21]), .B1(d5[21]), .C1(GND_net), .D1(GND_net), .CIN(n11197), 
          .COUT(n11198), .S0(d5_71__N_706[20]), .S1(d5_71__N_706[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1088_22.INIT0 = 16'h5666;
    defparam add_1088_22.INIT1 = 16'h5666;
    defparam add_1088_22.INJECT1_0 = "NO";
    defparam add_1088_22.INJECT1_1 = "NO";
    CCU2D add_1088_20 (.A0(d4[18]), .B0(d5[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[19]), .B1(d5[19]), .C1(GND_net), .D1(GND_net), .CIN(n11196), 
          .COUT(n11197), .S0(d5_71__N_706[18]), .S1(d5_71__N_706[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1088_20.INIT0 = 16'h5666;
    defparam add_1088_20.INIT1 = 16'h5666;
    defparam add_1088_20.INJECT1_0 = "NO";
    defparam add_1088_20.INJECT1_1 = "NO";
    CCU2D add_1088_18 (.A0(d4[16]), .B0(d5[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[17]), .B1(d5[17]), .C1(GND_net), .D1(GND_net), .CIN(n11195), 
          .COUT(n11196), .S0(d5_71__N_706[16]), .S1(d5_71__N_706[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1088_18.INIT0 = 16'h5666;
    defparam add_1088_18.INIT1 = 16'h5666;
    defparam add_1088_18.INJECT1_0 = "NO";
    defparam add_1088_18.INJECT1_1 = "NO";
    CCU2D add_1088_16 (.A0(d4[14]), .B0(d5[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[15]), .B1(d5[15]), .C1(GND_net), .D1(GND_net), .CIN(n11194), 
          .COUT(n11195), .S0(d5_71__N_706[14]), .S1(d5_71__N_706[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1088_16.INIT0 = 16'h5666;
    defparam add_1088_16.INIT1 = 16'h5666;
    defparam add_1088_16.INJECT1_0 = "NO";
    defparam add_1088_16.INJECT1_1 = "NO";
    CCU2D add_1088_14 (.A0(d4[12]), .B0(d5[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[13]), .B1(d5[13]), .C1(GND_net), .D1(GND_net), .CIN(n11193), 
          .COUT(n11194), .S0(d5_71__N_706[12]), .S1(d5_71__N_706[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1088_14.INIT0 = 16'h5666;
    defparam add_1088_14.INIT1 = 16'h5666;
    defparam add_1088_14.INJECT1_0 = "NO";
    defparam add_1088_14.INJECT1_1 = "NO";
    CCU2D add_1088_12 (.A0(d4[10]), .B0(d5[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[11]), .B1(d5[11]), .C1(GND_net), .D1(GND_net), .CIN(n11192), 
          .COUT(n11193), .S0(d5_71__N_706[10]), .S1(d5_71__N_706[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1088_12.INIT0 = 16'h5666;
    defparam add_1088_12.INIT1 = 16'h5666;
    defparam add_1088_12.INJECT1_0 = "NO";
    defparam add_1088_12.INJECT1_1 = "NO";
    CCU2D add_1088_10 (.A0(d4[8]), .B0(d5[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[9]), .B1(d5[9]), .C1(GND_net), .D1(GND_net), .CIN(n11191), 
          .COUT(n11192), .S0(d5_71__N_706[8]), .S1(d5_71__N_706[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1088_10.INIT0 = 16'h5666;
    defparam add_1088_10.INIT1 = 16'h5666;
    defparam add_1088_10.INJECT1_0 = "NO";
    defparam add_1088_10.INJECT1_1 = "NO";
    CCU2D add_1088_8 (.A0(d4[6]), .B0(d5[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[7]), .B1(d5[7]), .C1(GND_net), .D1(GND_net), .CIN(n11190), 
          .COUT(n11191), .S0(d5_71__N_706[6]), .S1(d5_71__N_706[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1088_8.INIT0 = 16'h5666;
    defparam add_1088_8.INIT1 = 16'h5666;
    defparam add_1088_8.INJECT1_0 = "NO";
    defparam add_1088_8.INJECT1_1 = "NO";
    CCU2D add_1088_6 (.A0(d4[4]), .B0(d5[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[5]), .B1(d5[5]), .C1(GND_net), .D1(GND_net), .CIN(n11189), 
          .COUT(n11190), .S0(d5_71__N_706[4]), .S1(d5_71__N_706[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1088_6.INIT0 = 16'h5666;
    defparam add_1088_6.INIT1 = 16'h5666;
    defparam add_1088_6.INJECT1_0 = "NO";
    defparam add_1088_6.INJECT1_1 = "NO";
    CCU2D add_1088_4 (.A0(d4[2]), .B0(d5[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[3]), .B1(d5[3]), .C1(GND_net), .D1(GND_net), .CIN(n11188), 
          .COUT(n11189), .S0(d5_71__N_706[2]), .S1(d5_71__N_706[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1088_4.INIT0 = 16'h5666;
    defparam add_1088_4.INIT1 = 16'h5666;
    defparam add_1088_4.INJECT1_0 = "NO";
    defparam add_1088_4.INJECT1_1 = "NO";
    CCU2D add_1088_2 (.A0(d4[0]), .B0(d5[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[1]), .B1(d5[1]), .C1(GND_net), .D1(GND_net), .COUT(n11188), 
          .S1(d5_71__N_706[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1088_2.INIT0 = 16'h7000;
    defparam add_1088_2.INIT1 = 16'h5666;
    defparam add_1088_2.INJECT1_0 = "NO";
    defparam add_1088_2.INJECT1_1 = "NO";
    CCU2D add_1083_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11186), 
          .S0(n5492));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1083_cout.INIT0 = 16'h0000;
    defparam add_1083_cout.INIT1 = 16'h0000;
    defparam add_1083_cout.INJECT1_0 = "NO";
    defparam add_1083_cout.INJECT1_1 = "NO";
    CCU2D add_1083_36 (.A0(d3[34]), .B0(d4[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[35]), .B1(d4[35]), .C1(GND_net), .D1(GND_net), .CIN(n11185), 
          .COUT(n11186), .S0(d4_71__N_634[34]), .S1(d4_71__N_634[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1083_36.INIT0 = 16'h5666;
    defparam add_1083_36.INIT1 = 16'h5666;
    defparam add_1083_36.INJECT1_0 = "NO";
    defparam add_1083_36.INJECT1_1 = "NO";
    CCU2D add_1083_34 (.A0(d3[32]), .B0(d4[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[33]), .B1(d4[33]), .C1(GND_net), .D1(GND_net), .CIN(n11184), 
          .COUT(n11185), .S0(d4_71__N_634[32]), .S1(d4_71__N_634[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1083_34.INIT0 = 16'h5666;
    defparam add_1083_34.INIT1 = 16'h5666;
    defparam add_1083_34.INJECT1_0 = "NO";
    defparam add_1083_34.INJECT1_1 = "NO";
    CCU2D add_1083_32 (.A0(d3[30]), .B0(d4[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[31]), .B1(d4[31]), .C1(GND_net), .D1(GND_net), .CIN(n11183), 
          .COUT(n11184), .S0(d4_71__N_634[30]), .S1(d4_71__N_634[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1083_32.INIT0 = 16'h5666;
    defparam add_1083_32.INIT1 = 16'h5666;
    defparam add_1083_32.INJECT1_0 = "NO";
    defparam add_1083_32.INJECT1_1 = "NO";
    CCU2D add_1083_30 (.A0(d3[28]), .B0(d4[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[29]), .B1(d4[29]), .C1(GND_net), .D1(GND_net), .CIN(n11182), 
          .COUT(n11183), .S0(d4_71__N_634[28]), .S1(d4_71__N_634[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1083_30.INIT0 = 16'h5666;
    defparam add_1083_30.INIT1 = 16'h5666;
    defparam add_1083_30.INJECT1_0 = "NO";
    defparam add_1083_30.INJECT1_1 = "NO";
    CCU2D add_1083_28 (.A0(d3[26]), .B0(d4[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[27]), .B1(d4[27]), .C1(GND_net), .D1(GND_net), .CIN(n11181), 
          .COUT(n11182), .S0(d4_71__N_634[26]), .S1(d4_71__N_634[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1083_28.INIT0 = 16'h5666;
    defparam add_1083_28.INIT1 = 16'h5666;
    defparam add_1083_28.INJECT1_0 = "NO";
    defparam add_1083_28.INJECT1_1 = "NO";
    CCU2D add_1083_26 (.A0(d3[24]), .B0(d4[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[25]), .B1(d4[25]), .C1(GND_net), .D1(GND_net), .CIN(n11180), 
          .COUT(n11181), .S0(d4_71__N_634[24]), .S1(d4_71__N_634[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1083_26.INIT0 = 16'h5666;
    defparam add_1083_26.INIT1 = 16'h5666;
    defparam add_1083_26.INJECT1_0 = "NO";
    defparam add_1083_26.INJECT1_1 = "NO";
    CCU2D add_1083_24 (.A0(d3[22]), .B0(d4[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[23]), .B1(d4[23]), .C1(GND_net), .D1(GND_net), .CIN(n11179), 
          .COUT(n11180), .S0(d4_71__N_634[22]), .S1(d4_71__N_634[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1083_24.INIT0 = 16'h5666;
    defparam add_1083_24.INIT1 = 16'h5666;
    defparam add_1083_24.INJECT1_0 = "NO";
    defparam add_1083_24.INJECT1_1 = "NO";
    CCU2D add_1083_22 (.A0(d3[20]), .B0(d4[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[21]), .B1(d4[21]), .C1(GND_net), .D1(GND_net), .CIN(n11178), 
          .COUT(n11179), .S0(d4_71__N_634[20]), .S1(d4_71__N_634[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1083_22.INIT0 = 16'h5666;
    defparam add_1083_22.INIT1 = 16'h5666;
    defparam add_1083_22.INJECT1_0 = "NO";
    defparam add_1083_22.INJECT1_1 = "NO";
    CCU2D add_1083_20 (.A0(d3[18]), .B0(d4[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[19]), .B1(d4[19]), .C1(GND_net), .D1(GND_net), .CIN(n11177), 
          .COUT(n11178), .S0(d4_71__N_634[18]), .S1(d4_71__N_634[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1083_20.INIT0 = 16'h5666;
    defparam add_1083_20.INIT1 = 16'h5666;
    defparam add_1083_20.INJECT1_0 = "NO";
    defparam add_1083_20.INJECT1_1 = "NO";
    CCU2D add_1083_18 (.A0(d3[16]), .B0(d4[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[17]), .B1(d4[17]), .C1(GND_net), .D1(GND_net), .CIN(n11176), 
          .COUT(n11177), .S0(d4_71__N_634[16]), .S1(d4_71__N_634[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1083_18.INIT0 = 16'h5666;
    defparam add_1083_18.INIT1 = 16'h5666;
    defparam add_1083_18.INJECT1_0 = "NO";
    defparam add_1083_18.INJECT1_1 = "NO";
    CCU2D add_1083_16 (.A0(d3[14]), .B0(d4[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[15]), .B1(d4[15]), .C1(GND_net), .D1(GND_net), .CIN(n11175), 
          .COUT(n11176), .S0(d4_71__N_634[14]), .S1(d4_71__N_634[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1083_16.INIT0 = 16'h5666;
    defparam add_1083_16.INIT1 = 16'h5666;
    defparam add_1083_16.INJECT1_0 = "NO";
    defparam add_1083_16.INJECT1_1 = "NO";
    CCU2D add_1083_14 (.A0(d3[12]), .B0(d4[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[13]), .B1(d4[13]), .C1(GND_net), .D1(GND_net), .CIN(n11174), 
          .COUT(n11175), .S0(d4_71__N_634[12]), .S1(d4_71__N_634[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1083_14.INIT0 = 16'h5666;
    defparam add_1083_14.INIT1 = 16'h5666;
    defparam add_1083_14.INJECT1_0 = "NO";
    defparam add_1083_14.INJECT1_1 = "NO";
    CCU2D add_1083_12 (.A0(d3[10]), .B0(d4[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[11]), .B1(d4[11]), .C1(GND_net), .D1(GND_net), .CIN(n11173), 
          .COUT(n11174), .S0(d4_71__N_634[10]), .S1(d4_71__N_634[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1083_12.INIT0 = 16'h5666;
    defparam add_1083_12.INIT1 = 16'h5666;
    defparam add_1083_12.INJECT1_0 = "NO";
    defparam add_1083_12.INJECT1_1 = "NO";
    CCU2D add_1083_10 (.A0(d3[8]), .B0(d4[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[9]), .B1(d4[9]), .C1(GND_net), .D1(GND_net), .CIN(n11172), 
          .COUT(n11173), .S0(d4_71__N_634[8]), .S1(d4_71__N_634[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1083_10.INIT0 = 16'h5666;
    defparam add_1083_10.INIT1 = 16'h5666;
    defparam add_1083_10.INJECT1_0 = "NO";
    defparam add_1083_10.INJECT1_1 = "NO";
    CCU2D add_1083_8 (.A0(d3[6]), .B0(d4[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[7]), .B1(d4[7]), .C1(GND_net), .D1(GND_net), .CIN(n11171), 
          .COUT(n11172), .S0(d4_71__N_634[6]), .S1(d4_71__N_634[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1083_8.INIT0 = 16'h5666;
    defparam add_1083_8.INIT1 = 16'h5666;
    defparam add_1083_8.INJECT1_0 = "NO";
    defparam add_1083_8.INJECT1_1 = "NO";
    CCU2D add_1083_6 (.A0(d3[4]), .B0(d4[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[5]), .B1(d4[5]), .C1(GND_net), .D1(GND_net), .CIN(n11170), 
          .COUT(n11171), .S0(d4_71__N_634[4]), .S1(d4_71__N_634[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1083_6.INIT0 = 16'h5666;
    defparam add_1083_6.INIT1 = 16'h5666;
    defparam add_1083_6.INJECT1_0 = "NO";
    defparam add_1083_6.INJECT1_1 = "NO";
    CCU2D add_1083_4 (.A0(d3[2]), .B0(d4[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[3]), .B1(d4[3]), .C1(GND_net), .D1(GND_net), .CIN(n11169), 
          .COUT(n11170), .S0(d4_71__N_634[2]), .S1(d4_71__N_634[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1083_4.INIT0 = 16'h5666;
    defparam add_1083_4.INIT1 = 16'h5666;
    defparam add_1083_4.INJECT1_0 = "NO";
    defparam add_1083_4.INJECT1_1 = "NO";
    CCU2D add_1083_2 (.A0(d3[0]), .B0(d4[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[1]), .B1(d4[1]), .C1(GND_net), .D1(GND_net), .COUT(n11169), 
          .S1(d4_71__N_634[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1083_2.INIT0 = 16'h7000;
    defparam add_1083_2.INIT1 = 16'h5666;
    defparam add_1083_2.INJECT1_0 = "NO";
    defparam add_1083_2.INJECT1_1 = "NO";
    CCU2D add_1078_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11167), 
          .S0(n5340));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1078_cout.INIT0 = 16'h0000;
    defparam add_1078_cout.INIT1 = 16'h0000;
    defparam add_1078_cout.INJECT1_0 = "NO";
    defparam add_1078_cout.INJECT1_1 = "NO";
    CCU2D add_1078_36 (.A0(d2[34]), .B0(d3[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[35]), .B1(d3[35]), .C1(GND_net), .D1(GND_net), .CIN(n11166), 
          .COUT(n11167), .S0(d3_71__N_562[34]), .S1(d3_71__N_562[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1078_36.INIT0 = 16'h5666;
    defparam add_1078_36.INIT1 = 16'h5666;
    defparam add_1078_36.INJECT1_0 = "NO";
    defparam add_1078_36.INJECT1_1 = "NO";
    CCU2D add_1078_34 (.A0(d2[32]), .B0(d3[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[33]), .B1(d3[33]), .C1(GND_net), .D1(GND_net), .CIN(n11165), 
          .COUT(n11166), .S0(d3_71__N_562[32]), .S1(d3_71__N_562[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1078_34.INIT0 = 16'h5666;
    defparam add_1078_34.INIT1 = 16'h5666;
    defparam add_1078_34.INJECT1_0 = "NO";
    defparam add_1078_34.INJECT1_1 = "NO";
    CCU2D add_1078_32 (.A0(d2[30]), .B0(d3[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[31]), .B1(d3[31]), .C1(GND_net), .D1(GND_net), .CIN(n11164), 
          .COUT(n11165), .S0(d3_71__N_562[30]), .S1(d3_71__N_562[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1078_32.INIT0 = 16'h5666;
    defparam add_1078_32.INIT1 = 16'h5666;
    defparam add_1078_32.INJECT1_0 = "NO";
    defparam add_1078_32.INJECT1_1 = "NO";
    CCU2D add_1078_30 (.A0(d2[28]), .B0(d3[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[29]), .B1(d3[29]), .C1(GND_net), .D1(GND_net), .CIN(n11163), 
          .COUT(n11164), .S0(d3_71__N_562[28]), .S1(d3_71__N_562[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1078_30.INIT0 = 16'h5666;
    defparam add_1078_30.INIT1 = 16'h5666;
    defparam add_1078_30.INJECT1_0 = "NO";
    defparam add_1078_30.INJECT1_1 = "NO";
    CCU2D add_1078_28 (.A0(d2[26]), .B0(d3[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[27]), .B1(d3[27]), .C1(GND_net), .D1(GND_net), .CIN(n11162), 
          .COUT(n11163), .S0(d3_71__N_562[26]), .S1(d3_71__N_562[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1078_28.INIT0 = 16'h5666;
    defparam add_1078_28.INIT1 = 16'h5666;
    defparam add_1078_28.INJECT1_0 = "NO";
    defparam add_1078_28.INJECT1_1 = "NO";
    CCU2D add_1078_26 (.A0(d2[24]), .B0(d3[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[25]), .B1(d3[25]), .C1(GND_net), .D1(GND_net), .CIN(n11161), 
          .COUT(n11162), .S0(d3_71__N_562[24]), .S1(d3_71__N_562[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1078_26.INIT0 = 16'h5666;
    defparam add_1078_26.INIT1 = 16'h5666;
    defparam add_1078_26.INJECT1_0 = "NO";
    defparam add_1078_26.INJECT1_1 = "NO";
    CCU2D add_1078_24 (.A0(d2[22]), .B0(d3[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[23]), .B1(d3[23]), .C1(GND_net), .D1(GND_net), .CIN(n11160), 
          .COUT(n11161), .S0(d3_71__N_562[22]), .S1(d3_71__N_562[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1078_24.INIT0 = 16'h5666;
    defparam add_1078_24.INIT1 = 16'h5666;
    defparam add_1078_24.INJECT1_0 = "NO";
    defparam add_1078_24.INJECT1_1 = "NO";
    CCU2D add_1078_22 (.A0(d2[20]), .B0(d3[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[21]), .B1(d3[21]), .C1(GND_net), .D1(GND_net), .CIN(n11159), 
          .COUT(n11160), .S0(d3_71__N_562[20]), .S1(d3_71__N_562[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1078_22.INIT0 = 16'h5666;
    defparam add_1078_22.INIT1 = 16'h5666;
    defparam add_1078_22.INJECT1_0 = "NO";
    defparam add_1078_22.INJECT1_1 = "NO";
    CCU2D add_1078_20 (.A0(d2[18]), .B0(d3[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[19]), .B1(d3[19]), .C1(GND_net), .D1(GND_net), .CIN(n11158), 
          .COUT(n11159), .S0(d3_71__N_562[18]), .S1(d3_71__N_562[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1078_20.INIT0 = 16'h5666;
    defparam add_1078_20.INIT1 = 16'h5666;
    defparam add_1078_20.INJECT1_0 = "NO";
    defparam add_1078_20.INJECT1_1 = "NO";
    CCU2D add_1078_18 (.A0(d2[16]), .B0(d3[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[17]), .B1(d3[17]), .C1(GND_net), .D1(GND_net), .CIN(n11157), 
          .COUT(n11158), .S0(d3_71__N_562[16]), .S1(d3_71__N_562[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1078_18.INIT0 = 16'h5666;
    defparam add_1078_18.INIT1 = 16'h5666;
    defparam add_1078_18.INJECT1_0 = "NO";
    defparam add_1078_18.INJECT1_1 = "NO";
    CCU2D add_1078_16 (.A0(d2[14]), .B0(d3[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[15]), .B1(d3[15]), .C1(GND_net), .D1(GND_net), .CIN(n11156), 
          .COUT(n11157), .S0(d3_71__N_562[14]), .S1(d3_71__N_562[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1078_16.INIT0 = 16'h5666;
    defparam add_1078_16.INIT1 = 16'h5666;
    defparam add_1078_16.INJECT1_0 = "NO";
    defparam add_1078_16.INJECT1_1 = "NO";
    CCU2D add_1078_14 (.A0(d2[12]), .B0(d3[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[13]), .B1(d3[13]), .C1(GND_net), .D1(GND_net), .CIN(n11155), 
          .COUT(n11156), .S0(d3_71__N_562[12]), .S1(d3_71__N_562[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1078_14.INIT0 = 16'h5666;
    defparam add_1078_14.INIT1 = 16'h5666;
    defparam add_1078_14.INJECT1_0 = "NO";
    defparam add_1078_14.INJECT1_1 = "NO";
    CCU2D add_1078_12 (.A0(d2[10]), .B0(d3[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[11]), .B1(d3[11]), .C1(GND_net), .D1(GND_net), .CIN(n11154), 
          .COUT(n11155), .S0(d3_71__N_562[10]), .S1(d3_71__N_562[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1078_12.INIT0 = 16'h5666;
    defparam add_1078_12.INIT1 = 16'h5666;
    defparam add_1078_12.INJECT1_0 = "NO";
    defparam add_1078_12.INJECT1_1 = "NO";
    CCU2D add_1078_10 (.A0(d2[8]), .B0(d3[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[9]), .B1(d3[9]), .C1(GND_net), .D1(GND_net), .CIN(n11153), 
          .COUT(n11154), .S0(d3_71__N_562[8]), .S1(d3_71__N_562[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1078_10.INIT0 = 16'h5666;
    defparam add_1078_10.INIT1 = 16'h5666;
    defparam add_1078_10.INJECT1_0 = "NO";
    defparam add_1078_10.INJECT1_1 = "NO";
    CCU2D add_1078_8 (.A0(d2[6]), .B0(d3[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[7]), .B1(d3[7]), .C1(GND_net), .D1(GND_net), .CIN(n11152), 
          .COUT(n11153), .S0(d3_71__N_562[6]), .S1(d3_71__N_562[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1078_8.INIT0 = 16'h5666;
    defparam add_1078_8.INIT1 = 16'h5666;
    defparam add_1078_8.INJECT1_0 = "NO";
    defparam add_1078_8.INJECT1_1 = "NO";
    CCU2D add_1078_6 (.A0(d2[4]), .B0(d3[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[5]), .B1(d3[5]), .C1(GND_net), .D1(GND_net), .CIN(n11151), 
          .COUT(n11152), .S0(d3_71__N_562[4]), .S1(d3_71__N_562[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1078_6.INIT0 = 16'h5666;
    defparam add_1078_6.INIT1 = 16'h5666;
    defparam add_1078_6.INJECT1_0 = "NO";
    defparam add_1078_6.INJECT1_1 = "NO";
    CCU2D add_1078_4 (.A0(d2[2]), .B0(d3[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[3]), .B1(d3[3]), .C1(GND_net), .D1(GND_net), .CIN(n11150), 
          .COUT(n11151), .S0(d3_71__N_562[2]), .S1(d3_71__N_562[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1078_4.INIT0 = 16'h5666;
    defparam add_1078_4.INIT1 = 16'h5666;
    defparam add_1078_4.INJECT1_0 = "NO";
    defparam add_1078_4.INJECT1_1 = "NO";
    CCU2D add_1078_2 (.A0(d2[0]), .B0(d3[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[1]), .B1(d3[1]), .C1(GND_net), .D1(GND_net), .COUT(n11150), 
          .S1(d3_71__N_562[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1078_2.INIT0 = 16'h7000;
    defparam add_1078_2.INIT1 = 16'h5666;
    defparam add_1078_2.INJECT1_0 = "NO";
    defparam add_1078_2.INJECT1_1 = "NO";
    CCU2D add_1073_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11148), 
          .S0(n5188));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1073_cout.INIT0 = 16'h0000;
    defparam add_1073_cout.INIT1 = 16'h0000;
    defparam add_1073_cout.INJECT1_0 = "NO";
    defparam add_1073_cout.INJECT1_1 = "NO";
    CCU2D add_1073_36 (.A0(d1[34]), .B0(d2[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[35]), .B1(d2[35]), .C1(GND_net), .D1(GND_net), .CIN(n11147), 
          .COUT(n11148), .S0(d2_71__N_490[34]), .S1(d2_71__N_490[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1073_36.INIT0 = 16'h5666;
    defparam add_1073_36.INIT1 = 16'h5666;
    defparam add_1073_36.INJECT1_0 = "NO";
    defparam add_1073_36.INJECT1_1 = "NO";
    CCU2D add_1073_34 (.A0(d1[32]), .B0(d2[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[33]), .B1(d2[33]), .C1(GND_net), .D1(GND_net), .CIN(n11146), 
          .COUT(n11147), .S0(d2_71__N_490[32]), .S1(d2_71__N_490[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1073_34.INIT0 = 16'h5666;
    defparam add_1073_34.INIT1 = 16'h5666;
    defparam add_1073_34.INJECT1_0 = "NO";
    defparam add_1073_34.INJECT1_1 = "NO";
    CCU2D add_1073_32 (.A0(d1[30]), .B0(d2[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[31]), .B1(d2[31]), .C1(GND_net), .D1(GND_net), .CIN(n11145), 
          .COUT(n11146), .S0(d2_71__N_490[30]), .S1(d2_71__N_490[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1073_32.INIT0 = 16'h5666;
    defparam add_1073_32.INIT1 = 16'h5666;
    defparam add_1073_32.INJECT1_0 = "NO";
    defparam add_1073_32.INJECT1_1 = "NO";
    CCU2D add_1073_30 (.A0(d1[28]), .B0(d2[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[29]), .B1(d2[29]), .C1(GND_net), .D1(GND_net), .CIN(n11144), 
          .COUT(n11145), .S0(d2_71__N_490[28]), .S1(d2_71__N_490[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1073_30.INIT0 = 16'h5666;
    defparam add_1073_30.INIT1 = 16'h5666;
    defparam add_1073_30.INJECT1_0 = "NO";
    defparam add_1073_30.INJECT1_1 = "NO";
    CCU2D add_1073_28 (.A0(d1[26]), .B0(d2[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[27]), .B1(d2[27]), .C1(GND_net), .D1(GND_net), .CIN(n11143), 
          .COUT(n11144), .S0(d2_71__N_490[26]), .S1(d2_71__N_490[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1073_28.INIT0 = 16'h5666;
    defparam add_1073_28.INIT1 = 16'h5666;
    defparam add_1073_28.INJECT1_0 = "NO";
    defparam add_1073_28.INJECT1_1 = "NO";
    CCU2D add_1073_26 (.A0(d1[24]), .B0(d2[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[25]), .B1(d2[25]), .C1(GND_net), .D1(GND_net), .CIN(n11142), 
          .COUT(n11143), .S0(d2_71__N_490[24]), .S1(d2_71__N_490[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1073_26.INIT0 = 16'h5666;
    defparam add_1073_26.INIT1 = 16'h5666;
    defparam add_1073_26.INJECT1_0 = "NO";
    defparam add_1073_26.INJECT1_1 = "NO";
    CCU2D add_1073_24 (.A0(d1[22]), .B0(d2[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[23]), .B1(d2[23]), .C1(GND_net), .D1(GND_net), .CIN(n11141), 
          .COUT(n11142), .S0(d2_71__N_490[22]), .S1(d2_71__N_490[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1073_24.INIT0 = 16'h5666;
    defparam add_1073_24.INIT1 = 16'h5666;
    defparam add_1073_24.INJECT1_0 = "NO";
    defparam add_1073_24.INJECT1_1 = "NO";
    CCU2D add_1073_22 (.A0(d1[20]), .B0(d2[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[21]), .B1(d2[21]), .C1(GND_net), .D1(GND_net), .CIN(n11140), 
          .COUT(n11141), .S0(d2_71__N_490[20]), .S1(d2_71__N_490[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1073_22.INIT0 = 16'h5666;
    defparam add_1073_22.INIT1 = 16'h5666;
    defparam add_1073_22.INJECT1_0 = "NO";
    defparam add_1073_22.INJECT1_1 = "NO";
    CCU2D add_1073_20 (.A0(d1[18]), .B0(d2[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[19]), .B1(d2[19]), .C1(GND_net), .D1(GND_net), .CIN(n11139), 
          .COUT(n11140), .S0(d2_71__N_490[18]), .S1(d2_71__N_490[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1073_20.INIT0 = 16'h5666;
    defparam add_1073_20.INIT1 = 16'h5666;
    defparam add_1073_20.INJECT1_0 = "NO";
    defparam add_1073_20.INJECT1_1 = "NO";
    CCU2D add_1073_18 (.A0(d1[16]), .B0(d2[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[17]), .B1(d2[17]), .C1(GND_net), .D1(GND_net), .CIN(n11138), 
          .COUT(n11139), .S0(d2_71__N_490[16]), .S1(d2_71__N_490[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1073_18.INIT0 = 16'h5666;
    defparam add_1073_18.INIT1 = 16'h5666;
    defparam add_1073_18.INJECT1_0 = "NO";
    defparam add_1073_18.INJECT1_1 = "NO";
    CCU2D add_1073_16 (.A0(d1[14]), .B0(d2[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[15]), .B1(d2[15]), .C1(GND_net), .D1(GND_net), .CIN(n11137), 
          .COUT(n11138), .S0(d2_71__N_490[14]), .S1(d2_71__N_490[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1073_16.INIT0 = 16'h5666;
    defparam add_1073_16.INIT1 = 16'h5666;
    defparam add_1073_16.INJECT1_0 = "NO";
    defparam add_1073_16.INJECT1_1 = "NO";
    CCU2D add_1073_14 (.A0(d1[12]), .B0(d2[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[13]), .B1(d2[13]), .C1(GND_net), .D1(GND_net), .CIN(n11136), 
          .COUT(n11137), .S0(d2_71__N_490[12]), .S1(d2_71__N_490[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1073_14.INIT0 = 16'h5666;
    defparam add_1073_14.INIT1 = 16'h5666;
    defparam add_1073_14.INJECT1_0 = "NO";
    defparam add_1073_14.INJECT1_1 = "NO";
    CCU2D add_1073_12 (.A0(d1[10]), .B0(d2[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[11]), .B1(d2[11]), .C1(GND_net), .D1(GND_net), .CIN(n11135), 
          .COUT(n11136), .S0(d2_71__N_490[10]), .S1(d2_71__N_490[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1073_12.INIT0 = 16'h5666;
    defparam add_1073_12.INIT1 = 16'h5666;
    defparam add_1073_12.INJECT1_0 = "NO";
    defparam add_1073_12.INJECT1_1 = "NO";
    CCU2D add_1073_10 (.A0(d1[8]), .B0(d2[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[9]), .B1(d2[9]), .C1(GND_net), .D1(GND_net), .CIN(n11134), 
          .COUT(n11135), .S0(d2_71__N_490[8]), .S1(d2_71__N_490[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1073_10.INIT0 = 16'h5666;
    defparam add_1073_10.INIT1 = 16'h5666;
    defparam add_1073_10.INJECT1_0 = "NO";
    defparam add_1073_10.INJECT1_1 = "NO";
    CCU2D add_1073_8 (.A0(d1[6]), .B0(d2[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[7]), .B1(d2[7]), .C1(GND_net), .D1(GND_net), .CIN(n11133), 
          .COUT(n11134), .S0(d2_71__N_490[6]), .S1(d2_71__N_490[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1073_8.INIT0 = 16'h5666;
    defparam add_1073_8.INIT1 = 16'h5666;
    defparam add_1073_8.INJECT1_0 = "NO";
    defparam add_1073_8.INJECT1_1 = "NO";
    CCU2D add_1073_6 (.A0(d1[4]), .B0(d2[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[5]), .B1(d2[5]), .C1(GND_net), .D1(GND_net), .CIN(n11132), 
          .COUT(n11133), .S0(d2_71__N_490[4]), .S1(d2_71__N_490[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1073_6.INIT0 = 16'h5666;
    defparam add_1073_6.INIT1 = 16'h5666;
    defparam add_1073_6.INJECT1_0 = "NO";
    defparam add_1073_6.INJECT1_1 = "NO";
    CCU2D add_1073_4 (.A0(d1[2]), .B0(d2[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[3]), .B1(d2[3]), .C1(GND_net), .D1(GND_net), .CIN(n11131), 
          .COUT(n11132), .S0(d2_71__N_490[2]), .S1(d2_71__N_490[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1073_4.INIT0 = 16'h5666;
    defparam add_1073_4.INIT1 = 16'h5666;
    defparam add_1073_4.INJECT1_0 = "NO";
    defparam add_1073_4.INJECT1_1 = "NO";
    CCU2D add_1073_2 (.A0(d1[0]), .B0(d2[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[1]), .B1(d2[1]), .C1(GND_net), .D1(GND_net), .COUT(n11131), 
          .S1(d2_71__N_490[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1073_2.INIT0 = 16'h7000;
    defparam add_1073_2.INIT1 = 16'h5666;
    defparam add_1073_2.INJECT1_0 = "NO";
    defparam add_1073_2.INJECT1_1 = "NO";
    CCU2D add_1068_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11091), 
          .S0(n5036));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1068_cout.INIT0 = 16'h0000;
    defparam add_1068_cout.INIT1 = 16'h0000;
    defparam add_1068_cout.INJECT1_0 = "NO";
    defparam add_1068_cout.INJECT1_1 = "NO";
    CCU2D add_1068_36 (.A0(MixerOutCos[11]), .B0(d1[34]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[35]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11090), .COUT(n11091), .S0(d1_71__N_418[34]), 
          .S1(d1_71__N_418[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1068_36.INIT0 = 16'h5666;
    defparam add_1068_36.INIT1 = 16'h5666;
    defparam add_1068_36.INJECT1_0 = "NO";
    defparam add_1068_36.INJECT1_1 = "NO";
    CCU2D add_1068_34 (.A0(MixerOutCos[11]), .B0(d1[32]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[33]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11089), .COUT(n11090), .S0(d1_71__N_418[32]), 
          .S1(d1_71__N_418[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1068_34.INIT0 = 16'h5666;
    defparam add_1068_34.INIT1 = 16'h5666;
    defparam add_1068_34.INJECT1_0 = "NO";
    defparam add_1068_34.INJECT1_1 = "NO";
    CCU2D add_1068_32 (.A0(MixerOutCos[11]), .B0(d1[30]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11088), .COUT(n11089), .S0(d1_71__N_418[30]), 
          .S1(d1_71__N_418[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1068_32.INIT0 = 16'h5666;
    defparam add_1068_32.INIT1 = 16'h5666;
    defparam add_1068_32.INJECT1_0 = "NO";
    defparam add_1068_32.INJECT1_1 = "NO";
    CCU2D add_1068_30 (.A0(MixerOutCos[11]), .B0(d1[28]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11087), .COUT(n11088), .S0(d1_71__N_418[28]), 
          .S1(d1_71__N_418[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1068_30.INIT0 = 16'h5666;
    defparam add_1068_30.INIT1 = 16'h5666;
    defparam add_1068_30.INJECT1_0 = "NO";
    defparam add_1068_30.INJECT1_1 = "NO";
    CCU2D add_1068_28 (.A0(MixerOutCos[11]), .B0(d1[26]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11086), .COUT(n11087), .S0(d1_71__N_418[26]), 
          .S1(d1_71__N_418[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1068_28.INIT0 = 16'h5666;
    defparam add_1068_28.INIT1 = 16'h5666;
    defparam add_1068_28.INJECT1_0 = "NO";
    defparam add_1068_28.INJECT1_1 = "NO";
    CCU2D add_1068_26 (.A0(MixerOutCos[11]), .B0(d1[24]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11085), .COUT(n11086), .S0(d1_71__N_418[24]), 
          .S1(d1_71__N_418[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1068_26.INIT0 = 16'h5666;
    defparam add_1068_26.INIT1 = 16'h5666;
    defparam add_1068_26.INJECT1_0 = "NO";
    defparam add_1068_26.INJECT1_1 = "NO";
    CCU2D add_1068_24 (.A0(MixerOutCos[11]), .B0(d1[22]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11084), .COUT(n11085), .S0(d1_71__N_418[22]), 
          .S1(d1_71__N_418[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1068_24.INIT0 = 16'h5666;
    defparam add_1068_24.INIT1 = 16'h5666;
    defparam add_1068_24.INJECT1_0 = "NO";
    defparam add_1068_24.INJECT1_1 = "NO";
    CCU2D add_1068_22 (.A0(MixerOutCos[11]), .B0(d1[20]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11083), .COUT(n11084), .S0(d1_71__N_418[20]), 
          .S1(d1_71__N_418[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1068_22.INIT0 = 16'h5666;
    defparam add_1068_22.INIT1 = 16'h5666;
    defparam add_1068_22.INJECT1_0 = "NO";
    defparam add_1068_22.INJECT1_1 = "NO";
    CCU2D add_1068_20 (.A0(MixerOutCos[11]), .B0(d1[18]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11082), .COUT(n11083), .S0(d1_71__N_418[18]), 
          .S1(d1_71__N_418[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1068_20.INIT0 = 16'h5666;
    defparam add_1068_20.INIT1 = 16'h5666;
    defparam add_1068_20.INJECT1_0 = "NO";
    defparam add_1068_20.INJECT1_1 = "NO";
    CCU2D add_1068_18 (.A0(MixerOutCos[11]), .B0(d1[16]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11081), .COUT(n11082), .S0(d1_71__N_418[16]), 
          .S1(d1_71__N_418[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1068_18.INIT0 = 16'h5666;
    defparam add_1068_18.INIT1 = 16'h5666;
    defparam add_1068_18.INJECT1_0 = "NO";
    defparam add_1068_18.INJECT1_1 = "NO";
    CCU2D add_1068_16 (.A0(MixerOutCos[11]), .B0(d1[14]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11080), .COUT(n11081), .S0(d1_71__N_418[14]), 
          .S1(d1_71__N_418[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1068_16.INIT0 = 16'h5666;
    defparam add_1068_16.INIT1 = 16'h5666;
    defparam add_1068_16.INJECT1_0 = "NO";
    defparam add_1068_16.INJECT1_1 = "NO";
    CCU2D add_1068_14 (.A0(MixerOutCos[11]), .B0(d1[12]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11079), .COUT(n11080), .S0(d1_71__N_418[12]), 
          .S1(d1_71__N_418[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1068_14.INIT0 = 16'h5666;
    defparam add_1068_14.INIT1 = 16'h5666;
    defparam add_1068_14.INJECT1_0 = "NO";
    defparam add_1068_14.INJECT1_1 = "NO";
    CCU2D add_1068_12 (.A0(MixerOutCos[10]), .B0(d1[10]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11078), .COUT(n11079), .S0(d1_71__N_418[10]), 
          .S1(d1_71__N_418[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1068_12.INIT0 = 16'h5666;
    defparam add_1068_12.INIT1 = 16'h5666;
    defparam add_1068_12.INJECT1_0 = "NO";
    defparam add_1068_12.INJECT1_1 = "NO";
    CCU2D add_1068_10 (.A0(MixerOutCos[8]), .B0(d1[8]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[9]), .B1(d1[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11077), .COUT(n11078), .S0(d1_71__N_418[8]), 
          .S1(d1_71__N_418[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1068_10.INIT0 = 16'h5666;
    defparam add_1068_10.INIT1 = 16'h5666;
    defparam add_1068_10.INJECT1_0 = "NO";
    defparam add_1068_10.INJECT1_1 = "NO";
    CCU2D add_1068_8 (.A0(MixerOutCos[6]), .B0(d1[6]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutCos[7]), .B1(d1[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11076), .COUT(n11077), .S0(d1_71__N_418[6]), .S1(d1_71__N_418[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1068_8.INIT0 = 16'h5666;
    defparam add_1068_8.INIT1 = 16'h5666;
    defparam add_1068_8.INJECT1_0 = "NO";
    defparam add_1068_8.INJECT1_1 = "NO";
    CCU2D add_1068_6 (.A0(MixerOutCos[4]), .B0(d1[4]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutCos[5]), .B1(d1[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11075), .COUT(n11076), .S0(d1_71__N_418[4]), .S1(d1_71__N_418[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1068_6.INIT0 = 16'h5666;
    defparam add_1068_6.INIT1 = 16'h5666;
    defparam add_1068_6.INJECT1_0 = "NO";
    defparam add_1068_6.INJECT1_1 = "NO";
    CCU2D add_1068_4 (.A0(MixerOutCos[2]), .B0(d1[2]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutCos[3]), .B1(d1[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11074), .COUT(n11075), .S0(d1_71__N_418[2]), .S1(d1_71__N_418[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1068_4.INIT0 = 16'h5666;
    defparam add_1068_4.INIT1 = 16'h5666;
    defparam add_1068_4.INJECT1_0 = "NO";
    defparam add_1068_4.INJECT1_1 = "NO";
    CCU2D add_1068_2 (.A0(MixerOutCos[0]), .B0(d1[0]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutCos[1]), .B1(d1[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n11074), .S1(d1_71__N_418[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1068_2.INIT0 = 16'h7000;
    defparam add_1068_2.INIT1 = 16'h5666;
    defparam add_1068_2.INJECT1_0 = "NO";
    defparam add_1068_2.INJECT1_1 = "NO";
    LUT4 i4914_2_lut (.A(d2[0]), .B(d3[0]), .Z(d3_71__N_562[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4914_2_lut.init = 16'h6666;
    CCU2D add_1123_37 (.A0(d9[35]), .B0(d_d9[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11745), 
          .S1(n6708));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1123_37.INIT0 = 16'h5999;
    defparam add_1123_37.INIT1 = 16'h0000;
    defparam add_1123_37.INJECT1_0 = "NO";
    defparam add_1123_37.INJECT1_1 = "NO";
    CCU2D add_1123_35 (.A0(d9[33]), .B0(d_d9[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[34]), .B1(d_d9[34]), .C1(GND_net), .D1(GND_net), .CIN(n11744), 
          .COUT(n11745));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1123_35.INIT0 = 16'h5999;
    defparam add_1123_35.INIT1 = 16'h5999;
    defparam add_1123_35.INJECT1_0 = "NO";
    defparam add_1123_35.INJECT1_1 = "NO";
    CCU2D add_1123_33 (.A0(d9[31]), .B0(d_d9[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[32]), .B1(d_d9[32]), .C1(GND_net), .D1(GND_net), .CIN(n11743), 
          .COUT(n11744));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1123_33.INIT0 = 16'h5999;
    defparam add_1123_33.INIT1 = 16'h5999;
    defparam add_1123_33.INJECT1_0 = "NO";
    defparam add_1123_33.INJECT1_1 = "NO";
    CCU2D add_1123_31 (.A0(d9[29]), .B0(d_d9[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[30]), .B1(d_d9[30]), .C1(GND_net), .D1(GND_net), .CIN(n11742), 
          .COUT(n11743));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1123_31.INIT0 = 16'h5999;
    defparam add_1123_31.INIT1 = 16'h5999;
    defparam add_1123_31.INJECT1_0 = "NO";
    defparam add_1123_31.INJECT1_1 = "NO";
    CCU2D add_1123_29 (.A0(d9[27]), .B0(d_d9[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[28]), .B1(d_d9[28]), .C1(GND_net), .D1(GND_net), .CIN(n11741), 
          .COUT(n11742));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1123_29.INIT0 = 16'h5999;
    defparam add_1123_29.INIT1 = 16'h5999;
    defparam add_1123_29.INJECT1_0 = "NO";
    defparam add_1123_29.INJECT1_1 = "NO";
    CCU2D add_1123_27 (.A0(d9[25]), .B0(d_d9[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[26]), .B1(d_d9[26]), .C1(GND_net), .D1(GND_net), .CIN(n11740), 
          .COUT(n11741));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1123_27.INIT0 = 16'h5999;
    defparam add_1123_27.INIT1 = 16'h5999;
    defparam add_1123_27.INJECT1_0 = "NO";
    defparam add_1123_27.INJECT1_1 = "NO";
    CCU2D add_1123_25 (.A0(d9[23]), .B0(d_d9[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[24]), .B1(d_d9[24]), .C1(GND_net), .D1(GND_net), .CIN(n11739), 
          .COUT(n11740));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1123_25.INIT0 = 16'h5999;
    defparam add_1123_25.INIT1 = 16'h5999;
    defparam add_1123_25.INJECT1_0 = "NO";
    defparam add_1123_25.INJECT1_1 = "NO";
    CCU2D add_1123_23 (.A0(d9[21]), .B0(d_d9[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[22]), .B1(d_d9[22]), .C1(GND_net), .D1(GND_net), .CIN(n11738), 
          .COUT(n11739));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1123_23.INIT0 = 16'h5999;
    defparam add_1123_23.INIT1 = 16'h5999;
    defparam add_1123_23.INJECT1_0 = "NO";
    defparam add_1123_23.INJECT1_1 = "NO";
    CCU2D add_1123_21 (.A0(d9[19]), .B0(d_d9[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[20]), .B1(d_d9[20]), .C1(GND_net), .D1(GND_net), .CIN(n11737), 
          .COUT(n11738));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1123_21.INIT0 = 16'h5999;
    defparam add_1123_21.INIT1 = 16'h5999;
    defparam add_1123_21.INJECT1_0 = "NO";
    defparam add_1123_21.INJECT1_1 = "NO";
    CCU2D add_1123_19 (.A0(d9[17]), .B0(d_d9[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[18]), .B1(d_d9[18]), .C1(GND_net), .D1(GND_net), .CIN(n11736), 
          .COUT(n11737));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1123_19.INIT0 = 16'h5999;
    defparam add_1123_19.INIT1 = 16'h5999;
    defparam add_1123_19.INJECT1_0 = "NO";
    defparam add_1123_19.INJECT1_1 = "NO";
    CCU2D add_1123_17 (.A0(d9[15]), .B0(d_d9[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[16]), .B1(d_d9[16]), .C1(GND_net), .D1(GND_net), .CIN(n11735), 
          .COUT(n11736));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1123_17.INIT0 = 16'h5999;
    defparam add_1123_17.INIT1 = 16'h5999;
    defparam add_1123_17.INJECT1_0 = "NO";
    defparam add_1123_17.INJECT1_1 = "NO";
    CCU2D add_1123_15 (.A0(d9[13]), .B0(d_d9[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[14]), .B1(d_d9[14]), .C1(GND_net), .D1(GND_net), .CIN(n11734), 
          .COUT(n11735));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1123_15.INIT0 = 16'h5999;
    defparam add_1123_15.INIT1 = 16'h5999;
    defparam add_1123_15.INJECT1_0 = "NO";
    defparam add_1123_15.INJECT1_1 = "NO";
    CCU2D add_1123_13 (.A0(d9[11]), .B0(d_d9[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[12]), .B1(d_d9[12]), .C1(GND_net), .D1(GND_net), .CIN(n11733), 
          .COUT(n11734));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1123_13.INIT0 = 16'h5999;
    defparam add_1123_13.INIT1 = 16'h5999;
    defparam add_1123_13.INJECT1_0 = "NO";
    defparam add_1123_13.INJECT1_1 = "NO";
    CCU2D add_1123_11 (.A0(d9[9]), .B0(d_d9[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[10]), .B1(d_d9[10]), .C1(GND_net), .D1(GND_net), .CIN(n11732), 
          .COUT(n11733));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1123_11.INIT0 = 16'h5999;
    defparam add_1123_11.INIT1 = 16'h5999;
    defparam add_1123_11.INJECT1_0 = "NO";
    defparam add_1123_11.INJECT1_1 = "NO";
    CCU2D add_1123_9 (.A0(d9[7]), .B0(d_d9[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[8]), .B1(d_d9[8]), .C1(GND_net), .D1(GND_net), .CIN(n11731), 
          .COUT(n11732));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1123_9.INIT0 = 16'h5999;
    defparam add_1123_9.INIT1 = 16'h5999;
    defparam add_1123_9.INJECT1_0 = "NO";
    defparam add_1123_9.INJECT1_1 = "NO";
    CCU2D add_1123_7 (.A0(d9[5]), .B0(d_d9[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[6]), .B1(d_d9[6]), .C1(GND_net), .D1(GND_net), .CIN(n11730), 
          .COUT(n11731));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1123_7.INIT0 = 16'h5999;
    defparam add_1123_7.INIT1 = 16'h5999;
    defparam add_1123_7.INJECT1_0 = "NO";
    defparam add_1123_7.INJECT1_1 = "NO";
    CCU2D add_1123_5 (.A0(d9[3]), .B0(d_d9[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[4]), .B1(d_d9[4]), .C1(GND_net), .D1(GND_net), .CIN(n11729), 
          .COUT(n11730));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1123_5.INIT0 = 16'h5999;
    defparam add_1123_5.INIT1 = 16'h5999;
    defparam add_1123_5.INJECT1_0 = "NO";
    defparam add_1123_5.INJECT1_1 = "NO";
    CCU2D add_1123_3 (.A0(d9[1]), .B0(d_d9[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[2]), .B1(d_d9[2]), .C1(GND_net), .D1(GND_net), .CIN(n11728), 
          .COUT(n11729));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1123_3.INIT0 = 16'h5999;
    defparam add_1123_3.INIT1 = 16'h5999;
    defparam add_1123_3.INJECT1_0 = "NO";
    defparam add_1123_3.INJECT1_1 = "NO";
    CCU2D add_1123_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d9[0]), .B1(d_d9[0]), .C1(GND_net), .D1(GND_net), .COUT(n11728));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1123_1.INIT0 = 16'h0000;
    defparam add_1123_1.INIT1 = 16'h5999;
    defparam add_1123_1.INJECT1_0 = "NO";
    defparam add_1123_1.INJECT1_1 = "NO";
    CCU2D add_1118_37 (.A0(d8[35]), .B0(d_d8[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11727), 
          .S0(d9_71__N_1675[35]), .S1(n6556));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1118_37.INIT0 = 16'h5999;
    defparam add_1118_37.INIT1 = 16'h0000;
    defparam add_1118_37.INJECT1_0 = "NO";
    defparam add_1118_37.INJECT1_1 = "NO";
    CCU2D add_1118_35 (.A0(d8[33]), .B0(d_d8[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[34]), .B1(d_d8[34]), .C1(GND_net), .D1(GND_net), .CIN(n11726), 
          .COUT(n11727), .S0(d9_71__N_1675[33]), .S1(d9_71__N_1675[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1118_35.INIT0 = 16'h5999;
    defparam add_1118_35.INIT1 = 16'h5999;
    defparam add_1118_35.INJECT1_0 = "NO";
    defparam add_1118_35.INJECT1_1 = "NO";
    CCU2D add_1118_33 (.A0(d8[31]), .B0(d_d8[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[32]), .B1(d_d8[32]), .C1(GND_net), .D1(GND_net), .CIN(n11725), 
          .COUT(n11726), .S0(d9_71__N_1675[31]), .S1(d9_71__N_1675[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1118_33.INIT0 = 16'h5999;
    defparam add_1118_33.INIT1 = 16'h5999;
    defparam add_1118_33.INJECT1_0 = "NO";
    defparam add_1118_33.INJECT1_1 = "NO";
    CCU2D add_1118_31 (.A0(d8[29]), .B0(d_d8[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[30]), .B1(d_d8[30]), .C1(GND_net), .D1(GND_net), .CIN(n11724), 
          .COUT(n11725), .S0(d9_71__N_1675[29]), .S1(d9_71__N_1675[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1118_31.INIT0 = 16'h5999;
    defparam add_1118_31.INIT1 = 16'h5999;
    defparam add_1118_31.INJECT1_0 = "NO";
    defparam add_1118_31.INJECT1_1 = "NO";
    CCU2D add_1118_29 (.A0(d8[27]), .B0(d_d8[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[28]), .B1(d_d8[28]), .C1(GND_net), .D1(GND_net), .CIN(n11723), 
          .COUT(n11724), .S0(d9_71__N_1675[27]), .S1(d9_71__N_1675[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1118_29.INIT0 = 16'h5999;
    defparam add_1118_29.INIT1 = 16'h5999;
    defparam add_1118_29.INJECT1_0 = "NO";
    defparam add_1118_29.INJECT1_1 = "NO";
    CCU2D add_1118_27 (.A0(d8[25]), .B0(d_d8[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[26]), .B1(d_d8[26]), .C1(GND_net), .D1(GND_net), .CIN(n11722), 
          .COUT(n11723), .S0(d9_71__N_1675[25]), .S1(d9_71__N_1675[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1118_27.INIT0 = 16'h5999;
    defparam add_1118_27.INIT1 = 16'h5999;
    defparam add_1118_27.INJECT1_0 = "NO";
    defparam add_1118_27.INJECT1_1 = "NO";
    CCU2D add_1118_25 (.A0(d8[23]), .B0(d_d8[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[24]), .B1(d_d8[24]), .C1(GND_net), .D1(GND_net), .CIN(n11721), 
          .COUT(n11722), .S0(d9_71__N_1675[23]), .S1(d9_71__N_1675[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1118_25.INIT0 = 16'h5999;
    defparam add_1118_25.INIT1 = 16'h5999;
    defparam add_1118_25.INJECT1_0 = "NO";
    defparam add_1118_25.INJECT1_1 = "NO";
    CCU2D add_1118_23 (.A0(d8[21]), .B0(d_d8[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[22]), .B1(d_d8[22]), .C1(GND_net), .D1(GND_net), .CIN(n11720), 
          .COUT(n11721), .S0(d9_71__N_1675[21]), .S1(d9_71__N_1675[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1118_23.INIT0 = 16'h5999;
    defparam add_1118_23.INIT1 = 16'h5999;
    defparam add_1118_23.INJECT1_0 = "NO";
    defparam add_1118_23.INJECT1_1 = "NO";
    CCU2D add_1118_21 (.A0(d8[19]), .B0(d_d8[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[20]), .B1(d_d8[20]), .C1(GND_net), .D1(GND_net), .CIN(n11719), 
          .COUT(n11720), .S0(d9_71__N_1675[19]), .S1(d9_71__N_1675[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1118_21.INIT0 = 16'h5999;
    defparam add_1118_21.INIT1 = 16'h5999;
    defparam add_1118_21.INJECT1_0 = "NO";
    defparam add_1118_21.INJECT1_1 = "NO";
    CCU2D add_1118_19 (.A0(d8[17]), .B0(d_d8[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[18]), .B1(d_d8[18]), .C1(GND_net), .D1(GND_net), .CIN(n11718), 
          .COUT(n11719), .S0(d9_71__N_1675[17]), .S1(d9_71__N_1675[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1118_19.INIT0 = 16'h5999;
    defparam add_1118_19.INIT1 = 16'h5999;
    defparam add_1118_19.INJECT1_0 = "NO";
    defparam add_1118_19.INJECT1_1 = "NO";
    CCU2D add_1118_17 (.A0(d8[15]), .B0(d_d8[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[16]), .B1(d_d8[16]), .C1(GND_net), .D1(GND_net), .CIN(n11717), 
          .COUT(n11718), .S0(d9_71__N_1675[15]), .S1(d9_71__N_1675[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1118_17.INIT0 = 16'h5999;
    defparam add_1118_17.INIT1 = 16'h5999;
    defparam add_1118_17.INJECT1_0 = "NO";
    defparam add_1118_17.INJECT1_1 = "NO";
    CCU2D add_1118_15 (.A0(d8[13]), .B0(d_d8[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[14]), .B1(d_d8[14]), .C1(GND_net), .D1(GND_net), .CIN(n11716), 
          .COUT(n11717), .S0(d9_71__N_1675[13]), .S1(d9_71__N_1675[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1118_15.INIT0 = 16'h5999;
    defparam add_1118_15.INIT1 = 16'h5999;
    defparam add_1118_15.INJECT1_0 = "NO";
    defparam add_1118_15.INJECT1_1 = "NO";
    CCU2D add_1118_13 (.A0(d8[11]), .B0(d_d8[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[12]), .B1(d_d8[12]), .C1(GND_net), .D1(GND_net), .CIN(n11715), 
          .COUT(n11716), .S0(d9_71__N_1675[11]), .S1(d9_71__N_1675[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1118_13.INIT0 = 16'h5999;
    defparam add_1118_13.INIT1 = 16'h5999;
    defparam add_1118_13.INJECT1_0 = "NO";
    defparam add_1118_13.INJECT1_1 = "NO";
    CCU2D add_1118_11 (.A0(d8[9]), .B0(d_d8[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[10]), .B1(d_d8[10]), .C1(GND_net), .D1(GND_net), .CIN(n11714), 
          .COUT(n11715), .S0(d9_71__N_1675[9]), .S1(d9_71__N_1675[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1118_11.INIT0 = 16'h5999;
    defparam add_1118_11.INIT1 = 16'h5999;
    defparam add_1118_11.INJECT1_0 = "NO";
    defparam add_1118_11.INJECT1_1 = "NO";
    CCU2D add_1118_9 (.A0(d8[7]), .B0(d_d8[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[8]), .B1(d_d8[8]), .C1(GND_net), .D1(GND_net), .CIN(n11713), 
          .COUT(n11714), .S0(d9_71__N_1675[7]), .S1(d9_71__N_1675[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1118_9.INIT0 = 16'h5999;
    defparam add_1118_9.INIT1 = 16'h5999;
    defparam add_1118_9.INJECT1_0 = "NO";
    defparam add_1118_9.INJECT1_1 = "NO";
    CCU2D add_1118_7 (.A0(d8[5]), .B0(d_d8[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[6]), .B1(d_d8[6]), .C1(GND_net), .D1(GND_net), .CIN(n11712), 
          .COUT(n11713), .S0(d9_71__N_1675[5]), .S1(d9_71__N_1675[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1118_7.INIT0 = 16'h5999;
    defparam add_1118_7.INIT1 = 16'h5999;
    defparam add_1118_7.INJECT1_0 = "NO";
    defparam add_1118_7.INJECT1_1 = "NO";
    CCU2D add_1118_5 (.A0(d8[3]), .B0(d_d8[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[4]), .B1(d_d8[4]), .C1(GND_net), .D1(GND_net), .CIN(n11711), 
          .COUT(n11712), .S0(d9_71__N_1675[3]), .S1(d9_71__N_1675[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1118_5.INIT0 = 16'h5999;
    defparam add_1118_5.INIT1 = 16'h5999;
    defparam add_1118_5.INJECT1_0 = "NO";
    defparam add_1118_5.INJECT1_1 = "NO";
    CCU2D add_1118_3 (.A0(d8[1]), .B0(d_d8[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[2]), .B1(d_d8[2]), .C1(GND_net), .D1(GND_net), .CIN(n11710), 
          .COUT(n11711), .S0(d9_71__N_1675[1]), .S1(d9_71__N_1675[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1118_3.INIT0 = 16'h5999;
    defparam add_1118_3.INIT1 = 16'h5999;
    defparam add_1118_3.INJECT1_0 = "NO";
    defparam add_1118_3.INJECT1_1 = "NO";
    CCU2D add_1118_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d8[0]), .B1(d_d8[0]), .C1(GND_net), .D1(GND_net), .COUT(n11710), 
          .S1(d9_71__N_1675[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1118_1.INIT0 = 16'h0000;
    defparam add_1118_1.INIT1 = 16'h5999;
    defparam add_1118_1.INJECT1_0 = "NO";
    defparam add_1118_1.INJECT1_1 = "NO";
    CCU2D add_1113_37 (.A0(d7[35]), .B0(d_d7[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11709), 
          .S0(d8_71__N_1603[35]), .S1(n6404));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1113_37.INIT0 = 16'h5999;
    defparam add_1113_37.INIT1 = 16'h0000;
    defparam add_1113_37.INJECT1_0 = "NO";
    defparam add_1113_37.INJECT1_1 = "NO";
    CCU2D add_1113_35 (.A0(d7[33]), .B0(d_d7[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[34]), .B1(d_d7[34]), .C1(GND_net), .D1(GND_net), .CIN(n11708), 
          .COUT(n11709), .S0(d8_71__N_1603[33]), .S1(d8_71__N_1603[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1113_35.INIT0 = 16'h5999;
    defparam add_1113_35.INIT1 = 16'h5999;
    defparam add_1113_35.INJECT1_0 = "NO";
    defparam add_1113_35.INJECT1_1 = "NO";
    CCU2D add_1113_33 (.A0(d7[31]), .B0(d_d7[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[32]), .B1(d_d7[32]), .C1(GND_net), .D1(GND_net), .CIN(n11707), 
          .COUT(n11708), .S0(d8_71__N_1603[31]), .S1(d8_71__N_1603[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1113_33.INIT0 = 16'h5999;
    defparam add_1113_33.INIT1 = 16'h5999;
    defparam add_1113_33.INJECT1_0 = "NO";
    defparam add_1113_33.INJECT1_1 = "NO";
    CCU2D add_1113_31 (.A0(d7[29]), .B0(d_d7[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[30]), .B1(d_d7[30]), .C1(GND_net), .D1(GND_net), .CIN(n11706), 
          .COUT(n11707), .S0(d8_71__N_1603[29]), .S1(d8_71__N_1603[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1113_31.INIT0 = 16'h5999;
    defparam add_1113_31.INIT1 = 16'h5999;
    defparam add_1113_31.INJECT1_0 = "NO";
    defparam add_1113_31.INJECT1_1 = "NO";
    CCU2D add_1113_29 (.A0(d7[27]), .B0(d_d7[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[28]), .B1(d_d7[28]), .C1(GND_net), .D1(GND_net), .CIN(n11705), 
          .COUT(n11706), .S0(d8_71__N_1603[27]), .S1(d8_71__N_1603[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1113_29.INIT0 = 16'h5999;
    defparam add_1113_29.INIT1 = 16'h5999;
    defparam add_1113_29.INJECT1_0 = "NO";
    defparam add_1113_29.INJECT1_1 = "NO";
    CCU2D add_1113_27 (.A0(d7[25]), .B0(d_d7[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[26]), .B1(d_d7[26]), .C1(GND_net), .D1(GND_net), .CIN(n11704), 
          .COUT(n11705), .S0(d8_71__N_1603[25]), .S1(d8_71__N_1603[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1113_27.INIT0 = 16'h5999;
    defparam add_1113_27.INIT1 = 16'h5999;
    defparam add_1113_27.INJECT1_0 = "NO";
    defparam add_1113_27.INJECT1_1 = "NO";
    CCU2D add_1113_25 (.A0(d7[23]), .B0(d_d7[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[24]), .B1(d_d7[24]), .C1(GND_net), .D1(GND_net), .CIN(n11703), 
          .COUT(n11704), .S0(d8_71__N_1603[23]), .S1(d8_71__N_1603[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1113_25.INIT0 = 16'h5999;
    defparam add_1113_25.INIT1 = 16'h5999;
    defparam add_1113_25.INJECT1_0 = "NO";
    defparam add_1113_25.INJECT1_1 = "NO";
    CCU2D add_1113_23 (.A0(d7[21]), .B0(d_d7[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[22]), .B1(d_d7[22]), .C1(GND_net), .D1(GND_net), .CIN(n11702), 
          .COUT(n11703), .S0(d8_71__N_1603[21]), .S1(d8_71__N_1603[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1113_23.INIT0 = 16'h5999;
    defparam add_1113_23.INIT1 = 16'h5999;
    defparam add_1113_23.INJECT1_0 = "NO";
    defparam add_1113_23.INJECT1_1 = "NO";
    CCU2D add_1113_21 (.A0(d7[19]), .B0(d_d7[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[20]), .B1(d_d7[20]), .C1(GND_net), .D1(GND_net), .CIN(n11701), 
          .COUT(n11702), .S0(d8_71__N_1603[19]), .S1(d8_71__N_1603[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1113_21.INIT0 = 16'h5999;
    defparam add_1113_21.INIT1 = 16'h5999;
    defparam add_1113_21.INJECT1_0 = "NO";
    defparam add_1113_21.INJECT1_1 = "NO";
    CCU2D add_1113_19 (.A0(d7[17]), .B0(d_d7[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[18]), .B1(d_d7[18]), .C1(GND_net), .D1(GND_net), .CIN(n11700), 
          .COUT(n11701), .S0(d8_71__N_1603[17]), .S1(d8_71__N_1603[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1113_19.INIT0 = 16'h5999;
    defparam add_1113_19.INIT1 = 16'h5999;
    defparam add_1113_19.INJECT1_0 = "NO";
    defparam add_1113_19.INJECT1_1 = "NO";
    CCU2D add_1113_17 (.A0(d7[15]), .B0(d_d7[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[16]), .B1(d_d7[16]), .C1(GND_net), .D1(GND_net), .CIN(n11699), 
          .COUT(n11700), .S0(d8_71__N_1603[15]), .S1(d8_71__N_1603[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1113_17.INIT0 = 16'h5999;
    defparam add_1113_17.INIT1 = 16'h5999;
    defparam add_1113_17.INJECT1_0 = "NO";
    defparam add_1113_17.INJECT1_1 = "NO";
    CCU2D add_1113_15 (.A0(d7[13]), .B0(d_d7[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[14]), .B1(d_d7[14]), .C1(GND_net), .D1(GND_net), .CIN(n11698), 
          .COUT(n11699), .S0(d8_71__N_1603[13]), .S1(d8_71__N_1603[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1113_15.INIT0 = 16'h5999;
    defparam add_1113_15.INIT1 = 16'h5999;
    defparam add_1113_15.INJECT1_0 = "NO";
    defparam add_1113_15.INJECT1_1 = "NO";
    CCU2D add_1113_13 (.A0(d7[11]), .B0(d_d7[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[12]), .B1(d_d7[12]), .C1(GND_net), .D1(GND_net), .CIN(n11697), 
          .COUT(n11698), .S0(d8_71__N_1603[11]), .S1(d8_71__N_1603[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1113_13.INIT0 = 16'h5999;
    defparam add_1113_13.INIT1 = 16'h5999;
    defparam add_1113_13.INJECT1_0 = "NO";
    defparam add_1113_13.INJECT1_1 = "NO";
    CCU2D add_1113_11 (.A0(d7[9]), .B0(d_d7[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[10]), .B1(d_d7[10]), .C1(GND_net), .D1(GND_net), .CIN(n11696), 
          .COUT(n11697), .S0(d8_71__N_1603[9]), .S1(d8_71__N_1603[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1113_11.INIT0 = 16'h5999;
    defparam add_1113_11.INIT1 = 16'h5999;
    defparam add_1113_11.INJECT1_0 = "NO";
    defparam add_1113_11.INJECT1_1 = "NO";
    CCU2D add_1113_9 (.A0(d7[7]), .B0(d_d7[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[8]), .B1(d_d7[8]), .C1(GND_net), .D1(GND_net), .CIN(n11695), 
          .COUT(n11696), .S0(d8_71__N_1603[7]), .S1(d8_71__N_1603[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1113_9.INIT0 = 16'h5999;
    defparam add_1113_9.INIT1 = 16'h5999;
    defparam add_1113_9.INJECT1_0 = "NO";
    defparam add_1113_9.INJECT1_1 = "NO";
    CCU2D add_1113_7 (.A0(d7[5]), .B0(d_d7[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[6]), .B1(d_d7[6]), .C1(GND_net), .D1(GND_net), .CIN(n11694), 
          .COUT(n11695), .S0(d8_71__N_1603[5]), .S1(d8_71__N_1603[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1113_7.INIT0 = 16'h5999;
    defparam add_1113_7.INIT1 = 16'h5999;
    defparam add_1113_7.INJECT1_0 = "NO";
    defparam add_1113_7.INJECT1_1 = "NO";
    CCU2D add_1113_5 (.A0(d7[3]), .B0(d_d7[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[4]), .B1(d_d7[4]), .C1(GND_net), .D1(GND_net), .CIN(n11693), 
          .COUT(n11694), .S0(d8_71__N_1603[3]), .S1(d8_71__N_1603[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1113_5.INIT0 = 16'h5999;
    defparam add_1113_5.INIT1 = 16'h5999;
    defparam add_1113_5.INJECT1_0 = "NO";
    defparam add_1113_5.INJECT1_1 = "NO";
    CCU2D add_1113_3 (.A0(d7[1]), .B0(d_d7[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[2]), .B1(d_d7[2]), .C1(GND_net), .D1(GND_net), .CIN(n11692), 
          .COUT(n11693), .S0(d8_71__N_1603[1]), .S1(d8_71__N_1603[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1113_3.INIT0 = 16'h5999;
    defparam add_1113_3.INIT1 = 16'h5999;
    defparam add_1113_3.INJECT1_0 = "NO";
    defparam add_1113_3.INJECT1_1 = "NO";
    CCU2D add_1113_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d7[0]), .B1(d_d7[0]), .C1(GND_net), .D1(GND_net), .COUT(n11692), 
          .S1(d8_71__N_1603[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1113_1.INIT0 = 16'h0000;
    defparam add_1113_1.INIT1 = 16'h5999;
    defparam add_1113_1.INJECT1_0 = "NO";
    defparam add_1113_1.INJECT1_1 = "NO";
    CCU2D add_1108_37 (.A0(d6[35]), .B0(d_d6[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11691), 
          .S0(d7_71__N_1531[35]), .S1(n6252));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1108_37.INIT0 = 16'h5999;
    defparam add_1108_37.INIT1 = 16'h0000;
    defparam add_1108_37.INJECT1_0 = "NO";
    defparam add_1108_37.INJECT1_1 = "NO";
    CCU2D add_1108_35 (.A0(d6[33]), .B0(d_d6[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[34]), .B1(d_d6[34]), .C1(GND_net), .D1(GND_net), .CIN(n11690), 
          .COUT(n11691), .S0(d7_71__N_1531[33]), .S1(d7_71__N_1531[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1108_35.INIT0 = 16'h5999;
    defparam add_1108_35.INIT1 = 16'h5999;
    defparam add_1108_35.INJECT1_0 = "NO";
    defparam add_1108_35.INJECT1_1 = "NO";
    CCU2D add_1108_33 (.A0(d6[31]), .B0(d_d6[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[32]), .B1(d_d6[32]), .C1(GND_net), .D1(GND_net), .CIN(n11689), 
          .COUT(n11690), .S0(d7_71__N_1531[31]), .S1(d7_71__N_1531[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1108_33.INIT0 = 16'h5999;
    defparam add_1108_33.INIT1 = 16'h5999;
    defparam add_1108_33.INJECT1_0 = "NO";
    defparam add_1108_33.INJECT1_1 = "NO";
    CCU2D add_1108_31 (.A0(d6[29]), .B0(d_d6[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[30]), .B1(d_d6[30]), .C1(GND_net), .D1(GND_net), .CIN(n11688), 
          .COUT(n11689), .S0(d7_71__N_1531[29]), .S1(d7_71__N_1531[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1108_31.INIT0 = 16'h5999;
    defparam add_1108_31.INIT1 = 16'h5999;
    defparam add_1108_31.INJECT1_0 = "NO";
    defparam add_1108_31.INJECT1_1 = "NO";
    CCU2D add_1108_29 (.A0(d6[27]), .B0(d_d6[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[28]), .B1(d_d6[28]), .C1(GND_net), .D1(GND_net), .CIN(n11687), 
          .COUT(n11688), .S0(d7_71__N_1531[27]), .S1(d7_71__N_1531[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1108_29.INIT0 = 16'h5999;
    defparam add_1108_29.INIT1 = 16'h5999;
    defparam add_1108_29.INJECT1_0 = "NO";
    defparam add_1108_29.INJECT1_1 = "NO";
    CCU2D add_1108_27 (.A0(d6[25]), .B0(d_d6[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[26]), .B1(d_d6[26]), .C1(GND_net), .D1(GND_net), .CIN(n11686), 
          .COUT(n11687), .S0(d7_71__N_1531[25]), .S1(d7_71__N_1531[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1108_27.INIT0 = 16'h5999;
    defparam add_1108_27.INIT1 = 16'h5999;
    defparam add_1108_27.INJECT1_0 = "NO";
    defparam add_1108_27.INJECT1_1 = "NO";
    CCU2D add_1108_25 (.A0(d6[23]), .B0(d_d6[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[24]), .B1(d_d6[24]), .C1(GND_net), .D1(GND_net), .CIN(n11685), 
          .COUT(n11686), .S0(d7_71__N_1531[23]), .S1(d7_71__N_1531[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1108_25.INIT0 = 16'h5999;
    defparam add_1108_25.INIT1 = 16'h5999;
    defparam add_1108_25.INJECT1_0 = "NO";
    defparam add_1108_25.INJECT1_1 = "NO";
    CCU2D add_1108_23 (.A0(d6[21]), .B0(d_d6[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[22]), .B1(d_d6[22]), .C1(GND_net), .D1(GND_net), .CIN(n11684), 
          .COUT(n11685), .S0(d7_71__N_1531[21]), .S1(d7_71__N_1531[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1108_23.INIT0 = 16'h5999;
    defparam add_1108_23.INIT1 = 16'h5999;
    defparam add_1108_23.INJECT1_0 = "NO";
    defparam add_1108_23.INJECT1_1 = "NO";
    CCU2D add_1108_21 (.A0(d6[19]), .B0(d_d6[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[20]), .B1(d_d6[20]), .C1(GND_net), .D1(GND_net), .CIN(n11683), 
          .COUT(n11684), .S0(d7_71__N_1531[19]), .S1(d7_71__N_1531[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1108_21.INIT0 = 16'h5999;
    defparam add_1108_21.INIT1 = 16'h5999;
    defparam add_1108_21.INJECT1_0 = "NO";
    defparam add_1108_21.INJECT1_1 = "NO";
    CCU2D add_1108_19 (.A0(d6[17]), .B0(d_d6[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[18]), .B1(d_d6[18]), .C1(GND_net), .D1(GND_net), .CIN(n11682), 
          .COUT(n11683), .S0(d7_71__N_1531[17]), .S1(d7_71__N_1531[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1108_19.INIT0 = 16'h5999;
    defparam add_1108_19.INIT1 = 16'h5999;
    defparam add_1108_19.INJECT1_0 = "NO";
    defparam add_1108_19.INJECT1_1 = "NO";
    CCU2D add_1108_17 (.A0(d6[15]), .B0(d_d6[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[16]), .B1(d_d6[16]), .C1(GND_net), .D1(GND_net), .CIN(n11681), 
          .COUT(n11682), .S0(d7_71__N_1531[15]), .S1(d7_71__N_1531[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1108_17.INIT0 = 16'h5999;
    defparam add_1108_17.INIT1 = 16'h5999;
    defparam add_1108_17.INJECT1_0 = "NO";
    defparam add_1108_17.INJECT1_1 = "NO";
    CCU2D add_1108_15 (.A0(d6[13]), .B0(d_d6[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[14]), .B1(d_d6[14]), .C1(GND_net), .D1(GND_net), .CIN(n11680), 
          .COUT(n11681), .S0(d7_71__N_1531[13]), .S1(d7_71__N_1531[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1108_15.INIT0 = 16'h5999;
    defparam add_1108_15.INIT1 = 16'h5999;
    defparam add_1108_15.INJECT1_0 = "NO";
    defparam add_1108_15.INJECT1_1 = "NO";
    CCU2D add_1108_13 (.A0(d6[11]), .B0(d_d6[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[12]), .B1(d_d6[12]), .C1(GND_net), .D1(GND_net), .CIN(n11679), 
          .COUT(n11680), .S0(d7_71__N_1531[11]), .S1(d7_71__N_1531[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1108_13.INIT0 = 16'h5999;
    defparam add_1108_13.INIT1 = 16'h5999;
    defparam add_1108_13.INJECT1_0 = "NO";
    defparam add_1108_13.INJECT1_1 = "NO";
    CCU2D add_1108_11 (.A0(d6[9]), .B0(d_d6[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[10]), .B1(d_d6[10]), .C1(GND_net), .D1(GND_net), .CIN(n11678), 
          .COUT(n11679), .S0(d7_71__N_1531[9]), .S1(d7_71__N_1531[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1108_11.INIT0 = 16'h5999;
    defparam add_1108_11.INIT1 = 16'h5999;
    defparam add_1108_11.INJECT1_0 = "NO";
    defparam add_1108_11.INJECT1_1 = "NO";
    CCU2D add_1108_9 (.A0(d6[7]), .B0(d_d6[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[8]), .B1(d_d6[8]), .C1(GND_net), .D1(GND_net), .CIN(n11677), 
          .COUT(n11678), .S0(d7_71__N_1531[7]), .S1(d7_71__N_1531[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1108_9.INIT0 = 16'h5999;
    defparam add_1108_9.INIT1 = 16'h5999;
    defparam add_1108_9.INJECT1_0 = "NO";
    defparam add_1108_9.INJECT1_1 = "NO";
    CCU2D add_1108_7 (.A0(d6[5]), .B0(d_d6[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[6]), .B1(d_d6[6]), .C1(GND_net), .D1(GND_net), .CIN(n11676), 
          .COUT(n11677), .S0(d7_71__N_1531[5]), .S1(d7_71__N_1531[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1108_7.INIT0 = 16'h5999;
    defparam add_1108_7.INIT1 = 16'h5999;
    defparam add_1108_7.INJECT1_0 = "NO";
    defparam add_1108_7.INJECT1_1 = "NO";
    CCU2D add_1108_5 (.A0(d6[3]), .B0(d_d6[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[4]), .B1(d_d6[4]), .C1(GND_net), .D1(GND_net), .CIN(n11675), 
          .COUT(n11676), .S0(d7_71__N_1531[3]), .S1(d7_71__N_1531[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1108_5.INIT0 = 16'h5999;
    defparam add_1108_5.INIT1 = 16'h5999;
    defparam add_1108_5.INJECT1_0 = "NO";
    defparam add_1108_5.INJECT1_1 = "NO";
    CCU2D add_1108_3 (.A0(d6[1]), .B0(d_d6[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[2]), .B1(d_d6[2]), .C1(GND_net), .D1(GND_net), .CIN(n11674), 
          .COUT(n11675), .S0(d7_71__N_1531[1]), .S1(d7_71__N_1531[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1108_3.INIT0 = 16'h5999;
    defparam add_1108_3.INIT1 = 16'h5999;
    defparam add_1108_3.INJECT1_0 = "NO";
    defparam add_1108_3.INJECT1_1 = "NO";
    CCU2D add_1108_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d6[0]), .B1(d_d6[0]), .C1(GND_net), .D1(GND_net), .COUT(n11674), 
          .S1(d7_71__N_1531[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1108_1.INIT0 = 16'h0000;
    defparam add_1108_1.INIT1 = 16'h5999;
    defparam add_1108_1.INJECT1_0 = "NO";
    defparam add_1108_1.INJECT1_1 = "NO";
    CCU2D add_1103_37 (.A0(d_tmp[35]), .B0(d_d_tmp[35]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11673), .S0(d6_71__N_1459[35]), .S1(n6100));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1103_37.INIT0 = 16'h5999;
    defparam add_1103_37.INIT1 = 16'h0000;
    defparam add_1103_37.INJECT1_0 = "NO";
    defparam add_1103_37.INJECT1_1 = "NO";
    CCU2D add_1103_35 (.A0(d_tmp[33]), .B0(d_d_tmp[33]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[34]), .B1(d_d_tmp[34]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11672), .COUT(n11673), .S0(d6_71__N_1459[33]), 
          .S1(d6_71__N_1459[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1103_35.INIT0 = 16'h5999;
    defparam add_1103_35.INIT1 = 16'h5999;
    defparam add_1103_35.INJECT1_0 = "NO";
    defparam add_1103_35.INJECT1_1 = "NO";
    CCU2D add_1103_33 (.A0(d_tmp[31]), .B0(d_d_tmp[31]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[32]), .B1(d_d_tmp[32]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11671), .COUT(n11672), .S0(d6_71__N_1459[31]), 
          .S1(d6_71__N_1459[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1103_33.INIT0 = 16'h5999;
    defparam add_1103_33.INIT1 = 16'h5999;
    defparam add_1103_33.INJECT1_0 = "NO";
    defparam add_1103_33.INJECT1_1 = "NO";
    CCU2D add_1103_31 (.A0(d_tmp[29]), .B0(d_d_tmp[29]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[30]), .B1(d_d_tmp[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11670), .COUT(n11671), .S0(d6_71__N_1459[29]), 
          .S1(d6_71__N_1459[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1103_31.INIT0 = 16'h5999;
    defparam add_1103_31.INIT1 = 16'h5999;
    defparam add_1103_31.INJECT1_0 = "NO";
    defparam add_1103_31.INJECT1_1 = "NO";
    CCU2D add_1103_29 (.A0(d_tmp[27]), .B0(d_d_tmp[27]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[28]), .B1(d_d_tmp[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11669), .COUT(n11670), .S0(d6_71__N_1459[27]), 
          .S1(d6_71__N_1459[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1103_29.INIT0 = 16'h5999;
    defparam add_1103_29.INIT1 = 16'h5999;
    defparam add_1103_29.INJECT1_0 = "NO";
    defparam add_1103_29.INJECT1_1 = "NO";
    CCU2D add_1103_27 (.A0(d_tmp[25]), .B0(d_d_tmp[25]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[26]), .B1(d_d_tmp[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11668), .COUT(n11669), .S0(d6_71__N_1459[25]), 
          .S1(d6_71__N_1459[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1103_27.INIT0 = 16'h5999;
    defparam add_1103_27.INIT1 = 16'h5999;
    defparam add_1103_27.INJECT1_0 = "NO";
    defparam add_1103_27.INJECT1_1 = "NO";
    CCU2D add_1103_25 (.A0(d_tmp[23]), .B0(d_d_tmp[23]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[24]), .B1(d_d_tmp[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11667), .COUT(n11668), .S0(d6_71__N_1459[23]), 
          .S1(d6_71__N_1459[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1103_25.INIT0 = 16'h5999;
    defparam add_1103_25.INIT1 = 16'h5999;
    defparam add_1103_25.INJECT1_0 = "NO";
    defparam add_1103_25.INJECT1_1 = "NO";
    CCU2D add_1103_23 (.A0(d_tmp[21]), .B0(d_d_tmp[21]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[22]), .B1(d_d_tmp[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11666), .COUT(n11667), .S0(d6_71__N_1459[21]), 
          .S1(d6_71__N_1459[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1103_23.INIT0 = 16'h5999;
    defparam add_1103_23.INIT1 = 16'h5999;
    defparam add_1103_23.INJECT1_0 = "NO";
    defparam add_1103_23.INJECT1_1 = "NO";
    CCU2D add_1103_21 (.A0(d_tmp[19]), .B0(d_d_tmp[19]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[20]), .B1(d_d_tmp[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11665), .COUT(n11666), .S0(d6_71__N_1459[19]), 
          .S1(d6_71__N_1459[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1103_21.INIT0 = 16'h5999;
    defparam add_1103_21.INIT1 = 16'h5999;
    defparam add_1103_21.INJECT1_0 = "NO";
    defparam add_1103_21.INJECT1_1 = "NO";
    CCU2D add_1103_19 (.A0(d_tmp[17]), .B0(d_d_tmp[17]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[18]), .B1(d_d_tmp[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11664), .COUT(n11665), .S0(d6_71__N_1459[17]), 
          .S1(d6_71__N_1459[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1103_19.INIT0 = 16'h5999;
    defparam add_1103_19.INIT1 = 16'h5999;
    defparam add_1103_19.INJECT1_0 = "NO";
    defparam add_1103_19.INJECT1_1 = "NO";
    CCU2D add_1103_17 (.A0(d_tmp[15]), .B0(d_d_tmp[15]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[16]), .B1(d_d_tmp[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11663), .COUT(n11664), .S0(d6_71__N_1459[15]), 
          .S1(d6_71__N_1459[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1103_17.INIT0 = 16'h5999;
    defparam add_1103_17.INIT1 = 16'h5999;
    defparam add_1103_17.INJECT1_0 = "NO";
    defparam add_1103_17.INJECT1_1 = "NO";
    CCU2D add_1103_15 (.A0(d_tmp[13]), .B0(d_d_tmp[13]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[14]), .B1(d_d_tmp[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11662), .COUT(n11663), .S0(d6_71__N_1459[13]), 
          .S1(d6_71__N_1459[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1103_15.INIT0 = 16'h5999;
    defparam add_1103_15.INIT1 = 16'h5999;
    defparam add_1103_15.INJECT1_0 = "NO";
    defparam add_1103_15.INJECT1_1 = "NO";
    CCU2D add_1103_13 (.A0(d_tmp[11]), .B0(d_d_tmp[11]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[12]), .B1(d_d_tmp[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11661), .COUT(n11662), .S0(d6_71__N_1459[11]), 
          .S1(d6_71__N_1459[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1103_13.INIT0 = 16'h5999;
    defparam add_1103_13.INIT1 = 16'h5999;
    defparam add_1103_13.INJECT1_0 = "NO";
    defparam add_1103_13.INJECT1_1 = "NO";
    CCU2D add_1103_11 (.A0(d_tmp[9]), .B0(d_d_tmp[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[10]), .B1(d_d_tmp[10]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11660), .COUT(n11661), .S0(d6_71__N_1459[9]), .S1(d6_71__N_1459[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1103_11.INIT0 = 16'h5999;
    defparam add_1103_11.INIT1 = 16'h5999;
    defparam add_1103_11.INJECT1_0 = "NO";
    defparam add_1103_11.INJECT1_1 = "NO";
    CCU2D add_1103_9 (.A0(d_tmp[7]), .B0(d_d_tmp[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[8]), .B1(d_d_tmp[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11659), .COUT(n11660), .S0(d6_71__N_1459[7]), .S1(d6_71__N_1459[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1103_9.INIT0 = 16'h5999;
    defparam add_1103_9.INIT1 = 16'h5999;
    defparam add_1103_9.INJECT1_0 = "NO";
    defparam add_1103_9.INJECT1_1 = "NO";
    CCU2D add_1103_7 (.A0(d_tmp[5]), .B0(d_d_tmp[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[6]), .B1(d_d_tmp[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11658), .COUT(n11659), .S0(d6_71__N_1459[5]), .S1(d6_71__N_1459[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1103_7.INIT0 = 16'h5999;
    defparam add_1103_7.INIT1 = 16'h5999;
    defparam add_1103_7.INJECT1_0 = "NO";
    defparam add_1103_7.INJECT1_1 = "NO";
    CCU2D add_1103_5 (.A0(d_tmp[3]), .B0(d_d_tmp[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[4]), .B1(d_d_tmp[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11657), .COUT(n11658), .S0(d6_71__N_1459[3]), .S1(d6_71__N_1459[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1103_5.INIT0 = 16'h5999;
    defparam add_1103_5.INIT1 = 16'h5999;
    defparam add_1103_5.INJECT1_0 = "NO";
    defparam add_1103_5.INJECT1_1 = "NO";
    CCU2D add_1103_3 (.A0(d_tmp[1]), .B0(d_d_tmp[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[2]), .B1(d_d_tmp[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11656), .COUT(n11657), .S0(d6_71__N_1459[1]), .S1(d6_71__N_1459[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1103_3.INIT0 = 16'h5999;
    defparam add_1103_3.INIT1 = 16'h5999;
    defparam add_1103_3.INJECT1_0 = "NO";
    defparam add_1103_3.INJECT1_1 = "NO";
    CCU2D add_1103_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[0]), .B1(d_d_tmp[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n11656), .S1(d6_71__N_1459[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1103_1.INIT0 = 16'h0000;
    defparam add_1103_1.INIT1 = 16'h5999;
    defparam add_1103_1.INJECT1_0 = "NO";
    defparam add_1103_1.INJECT1_1 = "NO";
    LUT4 i4915_2_lut (.A(d3[0]), .B(d4[0]), .Z(d4_71__N_634[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4915_2_lut.init = 16'h6666;
    FD1S3AX v_comb_66_rep_100 (.D(osc_clk_enable_744), .CK(osc_clk), .Q(osc_clk_enable_784)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_100.GSR = "ENABLED";
    LUT4 i4916_2_lut (.A(d4[0]), .B(d5[0]), .Z(d5_71__N_706[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4916_2_lut.init = 16'h6666;
    LUT4 mux_1236_i2_3_lut (.A(n6709[21]), .B(n6747[21]), .C(n6708), .Z(d10_71__N_1747[57])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1236_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1236_i3_3_lut (.A(n6709[22]), .B(n6747[22]), .C(n6708), .Z(d10_71__N_1747[58])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1236_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1236_i4_3_lut (.A(n6709[23]), .B(n6747[23]), .C(n6708), .Z(d10_71__N_1747[59])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1236_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1236_i5_3_lut (.A(n6709[24]), .B(n6747[24]), .C(n6708), .Z(d10_71__N_1747[60])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1236_i5_3_lut.init = 16'hcaca;
    LUT4 i4951_2_lut (.A(d1[36]), .B(d2[36]), .Z(n5189[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4951_2_lut.init = 16'h6666;
    LUT4 mux_1236_i6_3_lut (.A(n6709[25]), .B(n6747[25]), .C(n6708), .Z(d10_71__N_1747[61])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1236_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1236_i7_3_lut (.A(n6709[26]), .B(n6747[26]), .C(n6708), .Z(d10_71__N_1747[62])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1236_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1236_i8_3_lut (.A(n6709[27]), .B(n6747[27]), .C(n6708), .Z(d10_71__N_1747[63])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1236_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1236_i9_3_lut (.A(n6709[28]), .B(n6747[28]), .C(n6708), .Z(d10_71__N_1747[64])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1236_i9_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i61_3_lut (.A(\d10[60] ), .B(\d10[61] ), .C(\CICGain[0] ), 
         .Z(n61)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i61_3_lut.init = 16'hcaca;
    LUT4 mux_1236_i10_3_lut (.A(n6709[29]), .B(n6747[29]), .C(n6708), 
         .Z(d10_71__N_1747[65])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1236_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1236_i11_3_lut (.A(n6709[30]), .B(n6747[30]), .C(n6708), 
         .Z(d10_71__N_1747[66])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1236_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1236_i12_3_lut (.A(n6709[31]), .B(n6747[31]), .C(n6708), 
         .Z(d10_71__N_1747[67])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1236_i12_3_lut.init = 16'hcaca;
    FD1S3AX v_comb_66_rep_112 (.D(osc_clk_enable_744), .CK(osc_clk), .Q(osc_clk_enable_1384)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_112.GSR = "ENABLED";
    LUT4 mux_1236_i13_3_lut (.A(n6709[32]), .B(n6747[32]), .C(n6708), 
         .Z(d10_71__N_1747[68])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1236_i13_3_lut.init = 16'hcaca;
    LUT4 i4954_2_lut (.A(MixerOutCos[11]), .B(d1[36]), .Z(n5037[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4954_2_lut.init = 16'h6666;
    LUT4 mux_1236_i14_3_lut (.A(n6709[33]), .B(n6747[33]), .C(n6708), 
         .Z(d10_71__N_1747[69])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1236_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1236_i15_3_lut (.A(n6709[34]), .B(n6747[34]), .C(n6708), 
         .Z(d10_71__N_1747[70])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1236_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1236_i16_3_lut (.A(n6709[35]), .B(n6747[35]), .C(n6708), 
         .Z(d10_71__N_1747[71])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1236_i16_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i70_3_lut (.A(\d10[69] ), .B(\d10[70] ), .C(\CICGain[0] ), 
         .Z(n70)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i70_3_lut.init = 16'hcaca;
    LUT4 i5767_then_3_lut (.A(\CICGain[1] ), .B(\d10[59] ), .C(d10[57]), 
         .Z(n13404)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i5767_then_3_lut.init = 16'he4e4;
    LUT4 i5767_else_3_lut (.A(n61), .B(\CICGain[1] ), .C(d10[58]), .Z(n13403)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i5767_else_3_lut.init = 16'he2e2;
    LUT4 i5760_then_3_lut (.A(\CICGain[1] ), .B(\d10[60] ), .C(d10[58]), 
         .Z(n13407)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i5760_then_3_lut.init = 16'he4e4;
    LUT4 i5760_else_3_lut (.A(n62), .B(\CICGain[1] ), .C(\d10[59] ), .Z(n13406)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i5760_else_3_lut.init = 16'he2e2;
    LUT4 i4945_2_lut (.A(d3[36]), .B(d4[36]), .Z(n5493[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4945_2_lut.init = 16'h6666;
    LUT4 shift_right_31_i62_3_lut (.A(\d10[61] ), .B(\d10[62] ), .C(\CICGain[0] ), 
         .Z(n62)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i62_3_lut.init = 16'hcaca;
    FD1S3AX v_comb_66_rep_111 (.D(osc_clk_enable_744), .CK(osc_clk), .Q(osc_clk_enable_1334)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_111.GSR = "ENABLED";
    LUT4 shift_right_31_i63_3_lut (.A(\d10[62] ), .B(\d10[63] ), .C(\CICGain[0] ), 
         .Z(n63)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i63_3_lut.init = 16'hcaca;
    FD1S3AX v_comb_66_rep_110 (.D(osc_clk_enable_744), .CK(osc_clk), .Q(osc_clk_enable_1284)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_110.GSR = "ENABLED";
    LUT4 shift_right_31_i64_3_lut (.A(\d10[63] ), .B(\d10[64] ), .C(\CICGain[0] ), 
         .Z(n64)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i64_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i65_3_lut (.A(\d10[64] ), .B(\d10[65] ), .C(\CICGain[0] ), 
         .Z(n65)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i65_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i66_3_lut (.A(\d10[65] ), .B(\d10[66] ), .C(\CICGain[0] ), 
         .Z(n66)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i66_3_lut.init = 16'hcaca;
    CCU2D add_1070_17 (.A0(d1[50]), .B0(n5036), .C0(n5037[14]), .D0(MixerOutCos[11]), 
          .A1(d1[51]), .B1(n5036), .C1(n5037[15]), .D1(MixerOutCos[11]), 
          .CIN(n12055), .COUT(n12056), .S0(d1_71__N_418[50]), .S1(d1_71__N_418[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1070_17.INIT0 = 16'h74b8;
    defparam add_1070_17.INIT1 = 16'h74b8;
    defparam add_1070_17.INJECT1_0 = "NO";
    defparam add_1070_17.INJECT1_1 = "NO";
    CCU2D add_1089_18 (.A0(d4[52]), .B0(d5[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[53]), .B1(d5[53]), .C1(GND_net), .D1(GND_net), .CIN(n11911), 
          .COUT(n11912), .S0(n5645[16]), .S1(n5645[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1089_18.INIT0 = 16'h5666;
    defparam add_1089_18.INIT1 = 16'h5666;
    defparam add_1089_18.INJECT1_0 = "NO";
    defparam add_1089_18.INJECT1_1 = "NO";
    CCU2D add_1070_25 (.A0(d1[58]), .B0(n5036), .C0(n5037[22]), .D0(MixerOutCos[11]), 
          .A1(d1[59]), .B1(n5036), .C1(n5037[23]), .D1(MixerOutCos[11]), 
          .CIN(n12059), .COUT(n12060), .S0(d1_71__N_418[58]), .S1(d1_71__N_418[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1070_25.INIT0 = 16'h74b8;
    defparam add_1070_25.INIT1 = 16'h74b8;
    defparam add_1070_25.INJECT1_0 = "NO";
    defparam add_1070_25.INJECT1_1 = "NO";
    CCU2D add_1089_16 (.A0(d4[50]), .B0(d5[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[51]), .B1(d5[51]), .C1(GND_net), .D1(GND_net), .CIN(n11910), 
          .COUT(n11911), .S0(n5645[14]), .S1(n5645[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1089_16.INIT0 = 16'h5666;
    defparam add_1089_16.INIT1 = 16'h5666;
    defparam add_1089_16.INJECT1_0 = "NO";
    defparam add_1089_16.INJECT1_1 = "NO";
    CCU2D add_1069_10 (.A0(MixerOutCos[11]), .B0(d1[44]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[45]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12071), .COUT(n12072), .S0(n5037[8]), 
          .S1(n5037[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1069_10.INIT0 = 16'h5666;
    defparam add_1069_10.INIT1 = 16'h5666;
    defparam add_1069_10.INJECT1_0 = "NO";
    defparam add_1069_10.INJECT1_1 = "NO";
    CCU2D add_1069_8 (.A0(MixerOutCos[11]), .B0(d1[42]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[43]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12070), .COUT(n12071), .S0(n5037[6]), 
          .S1(n5037[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1069_8.INIT0 = 16'h5666;
    defparam add_1069_8.INIT1 = 16'h5666;
    defparam add_1069_8.INJECT1_0 = "NO";
    defparam add_1069_8.INJECT1_1 = "NO";
    CCU2D add_1069_6 (.A0(MixerOutCos[11]), .B0(d1[40]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[41]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12069), .COUT(n12070), .S0(n5037[4]), 
          .S1(n5037[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1069_6.INIT0 = 16'h5666;
    defparam add_1069_6.INIT1 = 16'h5666;
    defparam add_1069_6.INJECT1_0 = "NO";
    defparam add_1069_6.INJECT1_1 = "NO";
    CCU2D add_1069_4 (.A0(MixerOutCos[11]), .B0(d1[38]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[39]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12068), .COUT(n12069), .S0(n5037[2]), 
          .S1(n5037[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1069_4.INIT0 = 16'h5666;
    defparam add_1069_4.INIT1 = 16'h5666;
    defparam add_1069_4.INJECT1_0 = "NO";
    defparam add_1069_4.INJECT1_1 = "NO";
    CCU2D add_1069_2 (.A0(MixerOutCos[11]), .B0(d1[36]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[37]), .C1(GND_net), 
          .D1(GND_net), .COUT(n12068), .S1(n5037[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1069_2.INIT0 = 16'h7000;
    defparam add_1069_2.INIT1 = 16'h5666;
    defparam add_1069_2.INJECT1_0 = "NO";
    defparam add_1069_2.INJECT1_1 = "NO";
    LUT4 shift_right_31_i67_3_lut (.A(\d10[66] ), .B(\d10[67] ), .C(\CICGain[0] ), 
         .Z(n67)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i67_3_lut.init = 16'hcaca;
    CCU2D add_1070_37 (.A0(d1[70]), .B0(n5036), .C0(n5037[34]), .D0(MixerOutCos[11]), 
          .A1(d1[71]), .B1(n5036), .C1(n5037[35]), .D1(MixerOutCos[11]), 
          .CIN(n12065), .S0(d1_71__N_418[70]), .S1(d1_71__N_418[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1070_37.INIT0 = 16'h74b8;
    defparam add_1070_37.INIT1 = 16'h74b8;
    defparam add_1070_37.INJECT1_0 = "NO";
    defparam add_1070_37.INJECT1_1 = "NO";
    CCU2D add_1070_35 (.A0(d1[68]), .B0(n5036), .C0(n5037[32]), .D0(MixerOutCos[11]), 
          .A1(d1[69]), .B1(n5036), .C1(n5037[33]), .D1(MixerOutCos[11]), 
          .CIN(n12064), .COUT(n12065), .S0(d1_71__N_418[68]), .S1(d1_71__N_418[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1070_35.INIT0 = 16'h74b8;
    defparam add_1070_35.INIT1 = 16'h74b8;
    defparam add_1070_35.INJECT1_0 = "NO";
    defparam add_1070_35.INJECT1_1 = "NO";
    FD1S3IX count__i1 (.D(n375[1]), .CK(osc_clk), .CD(n8387), .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i1.GSR = "ENABLED";
    LUT4 i5728_2_lut (.A(n31), .B(n13507), .Z(n8387)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam i5728_2_lut.init = 16'hdddd;
    LUT4 i2906_2_lut (.A(n375[11]), .B(n31), .Z(count_15__N_1442[11])) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(86[13] 89[16])
    defparam i2906_2_lut.init = 16'hbbbb;
    LUT4 shift_right_31_i68_3_lut (.A(\d10[67] ), .B(\d10[68] ), .C(\CICGain[0] ), 
         .Z(n68)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i68_3_lut.init = 16'hcaca;
    CCU2D add_1070_33 (.A0(d1[66]), .B0(n5036), .C0(n5037[30]), .D0(MixerOutCos[11]), 
          .A1(d1[67]), .B1(n5036), .C1(n5037[31]), .D1(MixerOutCos[11]), 
          .CIN(n12063), .COUT(n12064), .S0(d1_71__N_418[66]), .S1(d1_71__N_418[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1070_33.INIT0 = 16'h74b8;
    defparam add_1070_33.INIT1 = 16'h74b8;
    defparam add_1070_33.INJECT1_0 = "NO";
    defparam add_1070_33.INJECT1_1 = "NO";
    CCU2D add_1070_31 (.A0(d1[64]), .B0(n5036), .C0(n5037[28]), .D0(MixerOutCos[11]), 
          .A1(d1[65]), .B1(n5036), .C1(n5037[29]), .D1(MixerOutCos[11]), 
          .CIN(n12062), .COUT(n12063), .S0(d1_71__N_418[64]), .S1(d1_71__N_418[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1070_31.INIT0 = 16'h74b8;
    defparam add_1070_31.INIT1 = 16'h74b8;
    defparam add_1070_31.INJECT1_0 = "NO";
    defparam add_1070_31.INJECT1_1 = "NO";
    FD1S3AX v_comb_66_rep_109 (.D(osc_clk_enable_744), .CK(osc_clk), .Q(osc_clk_enable_1234)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_109.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_108 (.D(osc_clk_enable_744), .CK(osc_clk), .Q(osc_clk_enable_1184)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_108.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_107 (.D(osc_clk_enable_744), .CK(osc_clk), .Q(osc_clk_enable_1134)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_107.GSR = "ENABLED";
    PFUMX i5802 (.BLUT(n13406), .ALUT(n13407), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[1]));
    FD1S3AX v_comb_66_rep_106 (.D(osc_clk_enable_744), .CK(osc_clk), .Q(osc_clk_enable_1084)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_106.GSR = "ENABLED";
    PFUMX i5800 (.BLUT(n13403), .ALUT(n13404), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[0]));
    CCU2D add_1070_23 (.A0(d1[56]), .B0(n5036), .C0(n5037[20]), .D0(MixerOutCos[11]), 
          .A1(d1[57]), .B1(n5036), .C1(n5037[21]), .D1(MixerOutCos[11]), 
          .CIN(n12058), .COUT(n12059), .S0(d1_71__N_418[56]), .S1(d1_71__N_418[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1070_23.INIT0 = 16'h74b8;
    defparam add_1070_23.INIT1 = 16'h74b8;
    defparam add_1070_23.INJECT1_0 = "NO";
    defparam add_1070_23.INJECT1_1 = "NO";
    FD1S3AX v_comb_66_rep_105 (.D(osc_clk_enable_744), .CK(osc_clk), .Q(osc_clk_enable_1034)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_105.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_104 (.D(osc_clk_enable_744), .CK(osc_clk), .Q(osc_clk_enable_984)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_104.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_103 (.D(osc_clk_enable_744), .CK(osc_clk), .Q(osc_clk_enable_934)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_103.GSR = "ENABLED";
    CCU2D add_1070_21 (.A0(d1[54]), .B0(n5036), .C0(n5037[18]), .D0(MixerOutCos[11]), 
          .A1(d1[55]), .B1(n5036), .C1(n5037[19]), .D1(MixerOutCos[11]), 
          .CIN(n12057), .COUT(n12058), .S0(d1_71__N_418[54]), .S1(d1_71__N_418[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1070_21.INIT0 = 16'h74b8;
    defparam add_1070_21.INIT1 = 16'h74b8;
    defparam add_1070_21.INJECT1_0 = "NO";
    defparam add_1070_21.INJECT1_1 = "NO";
    FD1S3AX v_comb_66_rep_102 (.D(osc_clk_enable_744), .CK(osc_clk), .Q(osc_clk_enable_884)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_102.GSR = "ENABLED";
    CCU2D add_1070_19 (.A0(d1[52]), .B0(n5036), .C0(n5037[16]), .D0(MixerOutCos[11]), 
          .A1(d1[53]), .B1(n5036), .C1(n5037[17]), .D1(MixerOutCos[11]), 
          .CIN(n12056), .COUT(n12057), .S0(d1_71__N_418[52]), .S1(d1_71__N_418[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1070_19.INIT0 = 16'h74b8;
    defparam add_1070_19.INIT1 = 16'h74b8;
    defparam add_1070_19.INJECT1_0 = "NO";
    defparam add_1070_19.INJECT1_1 = "NO";
    CCU2D add_1070_29 (.A0(d1[62]), .B0(n5036), .C0(n5037[26]), .D0(MixerOutCos[11]), 
          .A1(d1[63]), .B1(n5036), .C1(n5037[27]), .D1(MixerOutCos[11]), 
          .CIN(n12061), .COUT(n12062), .S0(d1_71__N_418[62]), .S1(d1_71__N_418[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1070_29.INIT0 = 16'h74b8;
    defparam add_1070_29.INIT1 = 16'h74b8;
    defparam add_1070_29.INJECT1_0 = "NO";
    defparam add_1070_29.INJECT1_1 = "NO";
    CCU2D add_1070_27 (.A0(d1[60]), .B0(n5036), .C0(n5037[24]), .D0(MixerOutCos[11]), 
          .A1(d1[61]), .B1(n5036), .C1(n5037[25]), .D1(MixerOutCos[11]), 
          .CIN(n12060), .COUT(n12061), .S0(d1_71__N_418[60]), .S1(d1_71__N_418[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1070_27.INIT0 = 16'h74b8;
    defparam add_1070_27.INIT1 = 16'h74b8;
    defparam add_1070_27.INJECT1_0 = "NO";
    defparam add_1070_27.INJECT1_1 = "NO";
    CCU2D add_1075_25 (.A0(d2[58]), .B0(n5188), .C0(n5189[22]), .D0(d1[58]), 
          .A1(d2[59]), .B1(n5188), .C1(n5189[23]), .D1(d1[59]), .CIN(n12018), 
          .COUT(n12019), .S0(d2_71__N_490[58]), .S1(d2_71__N_490[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1075_25.INIT0 = 16'h74b8;
    defparam add_1075_25.INIT1 = 16'h74b8;
    defparam add_1075_25.INJECT1_0 = "NO";
    defparam add_1075_25.INJECT1_1 = "NO";
    CCU2D add_1069_36 (.A0(MixerOutCos[11]), .B0(d1[70]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[71]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12084), .S0(n5037[34]), .S1(n5037[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1069_36.INIT0 = 16'h5666;
    defparam add_1069_36.INIT1 = 16'h5666;
    defparam add_1069_36.INJECT1_0 = "NO";
    defparam add_1069_36.INJECT1_1 = "NO";
    CCU2D add_1069_34 (.A0(MixerOutCos[11]), .B0(d1[68]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[69]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12083), .COUT(n12084), .S0(n5037[32]), 
          .S1(n5037[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1069_34.INIT0 = 16'h5666;
    defparam add_1069_34.INIT1 = 16'h5666;
    defparam add_1069_34.INJECT1_0 = "NO";
    defparam add_1069_34.INJECT1_1 = "NO";
    CCU2D add_1069_32 (.A0(MixerOutCos[11]), .B0(d1[66]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[67]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12082), .COUT(n12083), .S0(n5037[30]), 
          .S1(n5037[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1069_32.INIT0 = 16'h5666;
    defparam add_1069_32.INIT1 = 16'h5666;
    defparam add_1069_32.INJECT1_0 = "NO";
    defparam add_1069_32.INJECT1_1 = "NO";
    CCU2D add_1069_30 (.A0(MixerOutCos[11]), .B0(d1[64]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[65]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12081), .COUT(n12082), .S0(n5037[28]), 
          .S1(n5037[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1069_30.INIT0 = 16'h5666;
    defparam add_1069_30.INIT1 = 16'h5666;
    defparam add_1069_30.INJECT1_0 = "NO";
    defparam add_1069_30.INJECT1_1 = "NO";
    FD1S3AX v_comb_66_rep_101 (.D(osc_clk_enable_744), .CK(osc_clk), .Q(osc_clk_enable_834)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=183 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_101.GSR = "ENABLED";
    CCU2D add_1069_28 (.A0(MixerOutCos[11]), .B0(d1[62]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[63]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12080), .COUT(n12081), .S0(n5037[26]), 
          .S1(n5037[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1069_28.INIT0 = 16'h5666;
    defparam add_1069_28.INIT1 = 16'h5666;
    defparam add_1069_28.INJECT1_0 = "NO";
    defparam add_1069_28.INJECT1_1 = "NO";
    CCU2D add_1069_26 (.A0(MixerOutCos[11]), .B0(d1[60]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[61]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12079), .COUT(n12080), .S0(n5037[24]), 
          .S1(n5037[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1069_26.INIT0 = 16'h5666;
    defparam add_1069_26.INIT1 = 16'h5666;
    defparam add_1069_26.INJECT1_0 = "NO";
    defparam add_1069_26.INJECT1_1 = "NO";
    CCU2D add_1069_24 (.A0(MixerOutCos[11]), .B0(d1[58]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[59]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12078), .COUT(n12079), .S0(n5037[22]), 
          .S1(n5037[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1069_24.INIT0 = 16'h5666;
    defparam add_1069_24.INIT1 = 16'h5666;
    defparam add_1069_24.INJECT1_0 = "NO";
    defparam add_1069_24.INJECT1_1 = "NO";
    CCU2D add_1069_22 (.A0(MixerOutCos[11]), .B0(d1[56]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[57]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12077), .COUT(n12078), .S0(n5037[20]), 
          .S1(n5037[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1069_22.INIT0 = 16'h5666;
    defparam add_1069_22.INIT1 = 16'h5666;
    defparam add_1069_22.INJECT1_0 = "NO";
    defparam add_1069_22.INJECT1_1 = "NO";
    CCU2D add_1069_20 (.A0(MixerOutCos[11]), .B0(d1[54]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[55]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12076), .COUT(n12077), .S0(n5037[18]), 
          .S1(n5037[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1069_20.INIT0 = 16'h5666;
    defparam add_1069_20.INIT1 = 16'h5666;
    defparam add_1069_20.INJECT1_0 = "NO";
    defparam add_1069_20.INJECT1_1 = "NO";
    CCU2D add_1069_18 (.A0(MixerOutCos[11]), .B0(d1[52]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[53]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12075), .COUT(n12076), .S0(n5037[16]), 
          .S1(n5037[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1069_18.INIT0 = 16'h5666;
    defparam add_1069_18.INIT1 = 16'h5666;
    defparam add_1069_18.INJECT1_0 = "NO";
    defparam add_1069_18.INJECT1_1 = "NO";
    CCU2D add_1069_16 (.A0(MixerOutCos[11]), .B0(d1[50]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[51]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12074), .COUT(n12075), .S0(n5037[14]), 
          .S1(n5037[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1069_16.INIT0 = 16'h5666;
    defparam add_1069_16.INIT1 = 16'h5666;
    defparam add_1069_16.INJECT1_0 = "NO";
    defparam add_1069_16.INJECT1_1 = "NO";
    CCU2D add_1069_14 (.A0(MixerOutCos[11]), .B0(d1[48]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[49]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12073), .COUT(n12074), .S0(n5037[12]), 
          .S1(n5037[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1069_14.INIT0 = 16'h5666;
    defparam add_1069_14.INIT1 = 16'h5666;
    defparam add_1069_14.INJECT1_0 = "NO";
    defparam add_1069_14.INJECT1_1 = "NO";
    CCU2D add_1069_12 (.A0(MixerOutCos[11]), .B0(d1[46]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[47]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12072), .COUT(n12073), .S0(n5037[10]), 
          .S1(n5037[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1069_12.INIT0 = 16'h5666;
    defparam add_1069_12.INIT1 = 16'h5666;
    defparam add_1069_12.INJECT1_0 = "NO";
    defparam add_1069_12.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module AMDemodulator
//

module AMDemodulator (CIC1_out_clkSin, \CIC1_outSin[0] , CIC1_outCos, 
            \DataInReg_11__N_1856[0] , GND_net, \CIC1_outSin[1] , \CIC1_outSin[2] , 
            \CIC1_outSin[3] , \CIC1_outSin[4] , \CIC1_outSin[5] , MYLED_c_0, 
            MYLED_c_1, MYLED_c_2, MYLED_c_3, MYLED_c_4, MYLED_c_5, 
            \DataInReg_11__N_1856[1] , \DataInReg_11__N_1856[2] , \DataInReg_11__N_1856[3] , 
            \DataInReg_11__N_1856[4] , \DataInReg_11__N_1856[5] , \DataInReg_11__N_1856[6] , 
            \DataInReg_11__N_1856[7] , \DataInReg_11__N_1856[8] , \DemodOut[9] , 
            VCC_net) /* synthesis syn_module_defined=1 */ ;
    input CIC1_out_clkSin;
    input \CIC1_outSin[0] ;
    input [11:0]CIC1_outCos;
    output \DataInReg_11__N_1856[0] ;
    input GND_net;
    input \CIC1_outSin[1] ;
    input \CIC1_outSin[2] ;
    input \CIC1_outSin[3] ;
    input \CIC1_outSin[4] ;
    input \CIC1_outSin[5] ;
    input MYLED_c_0;
    input MYLED_c_1;
    input MYLED_c_2;
    input MYLED_c_3;
    input MYLED_c_4;
    input MYLED_c_5;
    output \DataInReg_11__N_1856[1] ;
    output \DataInReg_11__N_1856[2] ;
    output \DataInReg_11__N_1856[3] ;
    output \DataInReg_11__N_1856[4] ;
    output \DataInReg_11__N_1856[5] ;
    output \DataInReg_11__N_1856[6] ;
    output \DataInReg_11__N_1856[7] ;
    output \DataInReg_11__N_1856[8] ;
    output \DemodOut[9] ;
    input VCC_net;
    
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(82[6:21])
    wire [11:0]MultDataB;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(29[21:30])
    wire [11:0]MultDataC;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(33[21:30])
    wire [31:0]ISquare;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(24[14:21])
    wire [31:0]ISquare_31__N_1895;
    wire [15:0]d_out_d;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(20[21:28])
    wire [23:0]MultResult1;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(30[22:33])
    wire [23:0]MultResult2;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(35[22:33])
    wire [17:0]d_out_d_11__N_1894;
    
    wire n11796;
    wire [17:0]d_out_d_11__N_1874;
    
    wire d_out_d_11__N_1873;
    wire [17:0]d_out_d_11__N_1876;
    
    wire n11795, n11794, n11793, n11792;
    wire [17:0]d_out_d_11__N_1872;
    
    wire n11791, n12451;
    wire [17:0]d_out_d_11__N_2335;
    wire [17:0]d_out_d_11__N_2353;
    wire [17:0]d_out_d_11__N_1892;
    
    wire n11785, d_out_d_11__N_1891, n11244, n11243, n11242, n11241, 
        n11240, n11239, n11238, n11237, n11236, n11235, n11234, 
        n11233, n10995, d_out_d_11__N_1871, n10994, n10993, n10992, 
        n12447, n10991, d_out_d_11__N_1889, d_out_d_11__N_1887, d_out_d_11__N_1885, 
        d_out_d_11__N_1883, d_out_d_11__N_1881, d_out_d_11__N_1879, d_out_d_11__N_1877, 
        d_out_d_11__N_1875, n12450, n209, n12449, n12445;
    wire [17:0]d_out_d_11__N_1878;
    wire [17:0]d_out_d_11__N_1880;
    
    wire n12444, n12443, n12442, n11784, n12441, n12440, n12439, 
        n12438, n12432, n12431, n12430, n12429, n12428, n12427;
    wire [17:0]d_out_d_11__N_1884;
    wire [17:0]d_out_d_11__N_1882;
    
    wire n12426;
    wire [17:0]d_out_d_11__N_1888;
    wire [17:0]d_out_d_11__N_1886;
    
    wire n12425;
    wire [17:0]d_out_d_11__N_1890;
    
    wire n11783, n11782, n11781, n11780, n11779, n11778, n11758, 
        n11757, n11756, n11755, n11754, n11753, n11752, n11751, 
        n11750, n11654, n11653, n11652, n11651, n11650, n11649, 
        n11648, n11647, n11646, n12397, n12396, n12395, n12394, 
        n12393, n12392, n12391, n12390, n12389, n12383, n12382, 
        n12381, n12380, n12379, n12378, n12377, n12376, n12375, 
        n12369, n12368, n12367, n12366, n12365, n12364, n12363, 
        n12362, n12361, n12355, n12354, n12353, n12352, n12351, 
        n12350, n12349, n12348, n12347, n12341, n12340, n12339, 
        n12338, n12337, n12336, n12335;
    
    FD1S3AX MultDataB_i0 (.D(\CIC1_outSin[0] ), .CK(CIC1_out_clkSin), .Q(MultDataB[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i0.GSR = "ENABLED";
    FD1S3AX MultDataC_i0 (.D(CIC1_outCos[0]), .CK(CIC1_out_clkSin), .Q(MultDataC[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i0.GSR = "ENABLED";
    FD1S3AX ISquare_i1 (.D(ISquare_31__N_1895[0]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i1.GSR = "ENABLED";
    FD1S3AX d_out_i1 (.D(d_out_d[0]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i1.GSR = "ENABLED";
    LUT4 i4917_2_lut (.A(MultResult1[0]), .B(MultResult2[0]), .Z(ISquare_31__N_1895[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4917_2_lut.init = 16'h6666;
    FD1S3AX d_out_d__0_i1 (.D(d_out_d_11__N_1894[17]), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i1.GSR = "ENABLED";
    CCU2D add_453_13 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1873), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1874[17]), .B1(d_out_d_11__N_1873), 
          .C1(GND_net), .D1(GND_net), .CIN(n11796), .S0(d_out_d_11__N_1876[9]), 
          .S1(d_out_d_11__N_1876[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_453_13.INIT0 = 16'h5666;
    defparam add_453_13.INIT1 = 16'h5666;
    defparam add_453_13.INJECT1_0 = "NO";
    defparam add_453_13.INJECT1_1 = "NO";
    FD1S3AX MultDataB_i1 (.D(\CIC1_outSin[1] ), .CK(CIC1_out_clkSin), .Q(MultDataB[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i1.GSR = "ENABLED";
    FD1S3AX MultDataB_i2 (.D(\CIC1_outSin[2] ), .CK(CIC1_out_clkSin), .Q(MultDataB[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i2.GSR = "ENABLED";
    FD1S3AX MultDataB_i3 (.D(\CIC1_outSin[3] ), .CK(CIC1_out_clkSin), .Q(MultDataB[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i3.GSR = "ENABLED";
    FD1S3AX MultDataB_i4 (.D(\CIC1_outSin[4] ), .CK(CIC1_out_clkSin), .Q(MultDataB[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i4.GSR = "ENABLED";
    FD1S3AX MultDataB_i5 (.D(\CIC1_outSin[5] ), .CK(CIC1_out_clkSin), .Q(MultDataB[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i5.GSR = "ENABLED";
    FD1S3AX MultDataB_i6 (.D(MYLED_c_0), .CK(CIC1_out_clkSin), .Q(MultDataB[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i6.GSR = "ENABLED";
    FD1S3AX MultDataB_i7 (.D(MYLED_c_1), .CK(CIC1_out_clkSin), .Q(MultDataB[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i7.GSR = "ENABLED";
    FD1S3AX MultDataB_i8 (.D(MYLED_c_2), .CK(CIC1_out_clkSin), .Q(MultDataB[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i8.GSR = "ENABLED";
    FD1S3AX MultDataB_i9 (.D(MYLED_c_3), .CK(CIC1_out_clkSin), .Q(MultDataB[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i9.GSR = "ENABLED";
    FD1S3AX MultDataB_i10 (.D(MYLED_c_4), .CK(CIC1_out_clkSin), .Q(MultDataB[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i10.GSR = "ENABLED";
    FD1S3AX MultDataB_i11 (.D(MYLED_c_5), .CK(CIC1_out_clkSin), .Q(MultDataB[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i11.GSR = "ENABLED";
    FD1S3AX MultDataC_i1 (.D(CIC1_outCos[1]), .CK(CIC1_out_clkSin), .Q(MultDataC[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i1.GSR = "ENABLED";
    FD1S3AX MultDataC_i2 (.D(CIC1_outCos[2]), .CK(CIC1_out_clkSin), .Q(MultDataC[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i2.GSR = "ENABLED";
    FD1S3AX MultDataC_i3 (.D(CIC1_outCos[3]), .CK(CIC1_out_clkSin), .Q(MultDataC[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i3.GSR = "ENABLED";
    FD1S3AX MultDataC_i4 (.D(CIC1_outCos[4]), .CK(CIC1_out_clkSin), .Q(MultDataC[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i4.GSR = "ENABLED";
    FD1S3AX MultDataC_i5 (.D(CIC1_outCos[5]), .CK(CIC1_out_clkSin), .Q(MultDataC[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i5.GSR = "ENABLED";
    FD1S3AX MultDataC_i6 (.D(CIC1_outCos[6]), .CK(CIC1_out_clkSin), .Q(MultDataC[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i6.GSR = "ENABLED";
    FD1S3AX MultDataC_i7 (.D(CIC1_outCos[7]), .CK(CIC1_out_clkSin), .Q(MultDataC[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i7.GSR = "ENABLED";
    FD1S3AX MultDataC_i8 (.D(CIC1_outCos[8]), .CK(CIC1_out_clkSin), .Q(MultDataC[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i8.GSR = "ENABLED";
    FD1S3AX MultDataC_i9 (.D(CIC1_outCos[9]), .CK(CIC1_out_clkSin), .Q(MultDataC[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i9.GSR = "ENABLED";
    FD1S3AX MultDataC_i10 (.D(CIC1_outCos[10]), .CK(CIC1_out_clkSin), .Q(MultDataC[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i10.GSR = "ENABLED";
    FD1S3AX MultDataC_i11 (.D(CIC1_outCos[11]), .CK(CIC1_out_clkSin), .Q(MultDataC[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i11.GSR = "ENABLED";
    FD1S3AX ISquare_i2 (.D(ISquare_31__N_1895[1]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i2.GSR = "ENABLED";
    FD1S3AX ISquare_i3 (.D(ISquare_31__N_1895[2]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i3.GSR = "ENABLED";
    FD1S3AX ISquare_i4 (.D(ISquare_31__N_1895[3]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i4.GSR = "ENABLED";
    FD1S3AX ISquare_i5 (.D(ISquare_31__N_1895[4]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i5.GSR = "ENABLED";
    FD1S3AX ISquare_i6 (.D(ISquare_31__N_1895[5]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i6.GSR = "ENABLED";
    FD1S3AX ISquare_i7 (.D(ISquare_31__N_1895[6]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i7.GSR = "ENABLED";
    FD1S3AX ISquare_i8 (.D(ISquare_31__N_1895[7]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i8.GSR = "ENABLED";
    FD1S3AX ISquare_i9 (.D(ISquare_31__N_1895[8]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i9.GSR = "ENABLED";
    FD1S3AX ISquare_i10 (.D(ISquare_31__N_1895[9]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i10.GSR = "ENABLED";
    FD1S3AX ISquare_i11 (.D(ISquare_31__N_1895[10]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i11.GSR = "ENABLED";
    FD1S3AX ISquare_i12 (.D(ISquare_31__N_1895[11]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i12.GSR = "ENABLED";
    FD1S3AX ISquare_i13 (.D(ISquare_31__N_1895[12]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i13.GSR = "ENABLED";
    FD1S3AX ISquare_i14 (.D(ISquare_31__N_1895[13]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i14.GSR = "ENABLED";
    FD1S3AX ISquare_i15 (.D(ISquare_31__N_1895[14]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i15.GSR = "ENABLED";
    FD1S3AX ISquare_i16 (.D(ISquare_31__N_1895[15]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i16.GSR = "ENABLED";
    FD1S3AX ISquare_i17 (.D(ISquare_31__N_1895[16]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i17.GSR = "ENABLED";
    FD1S3AX ISquare_i18 (.D(ISquare_31__N_1895[17]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i18.GSR = "ENABLED";
    FD1S3AX ISquare_i19 (.D(ISquare_31__N_1895[18]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i19.GSR = "ENABLED";
    FD1S3AX ISquare_i20 (.D(ISquare_31__N_1895[19]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i20.GSR = "ENABLED";
    FD1S3AX ISquare_i21 (.D(ISquare_31__N_1895[20]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i21.GSR = "ENABLED";
    FD1S3AX ISquare_i22 (.D(ISquare_31__N_1895[21]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i22.GSR = "ENABLED";
    FD1S3AX ISquare_i23 (.D(ISquare_31__N_1895[22]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i23.GSR = "ENABLED";
    FD1S3AX ISquare_i24 (.D(ISquare_31__N_1895[23]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i24.GSR = "ENABLED";
    FD1S3AX ISquare_i25 (.D(ISquare_31__N_1895[24]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i25.GSR = "ENABLED";
    FD1S3AX d_out_i2 (.D(d_out_d[1]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i2.GSR = "ENABLED";
    FD1S3AX d_out_i3 (.D(d_out_d[2]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i3.GSR = "ENABLED";
    FD1S3AX d_out_i4 (.D(d_out_d[3]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i4.GSR = "ENABLED";
    FD1S3AX d_out_i5 (.D(d_out_d[4]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i5.GSR = "ENABLED";
    FD1S3AX d_out_i6 (.D(d_out_d[5]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i6.GSR = "ENABLED";
    FD1S3AX d_out_i7 (.D(d_out_d[6]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i7.GSR = "ENABLED";
    FD1S3AX d_out_i8 (.D(d_out_d[7]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i8.GSR = "ENABLED";
    FD1S3AX d_out_i9 (.D(d_out_d[8]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i9.GSR = "ENABLED";
    FD1S3AX d_out_i10 (.D(d_out_d[9]), .CK(CIC1_out_clkSin), .Q(\DemodOut[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=209, LSE_RLINE=214 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i10.GSR = "ENABLED";
    CCU2D add_453_11 (.A0(d_out_d_11__N_1874[6]), .B0(d_out_d_11__N_1874[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1874[7]), .B1(d_out_d_11__N_1874[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11795), .COUT(n11796), .S0(d_out_d_11__N_1876[7]), 
          .S1(d_out_d_11__N_1876[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_453_11.INIT0 = 16'h5999;
    defparam add_453_11.INIT1 = 16'h5999;
    defparam add_453_11.INJECT1_0 = "NO";
    defparam add_453_11.INJECT1_1 = "NO";
    CCU2D add_453_9 (.A0(ISquare[31]), .B0(d_out_d_11__N_1874[17]), .C0(d_out_d_11__N_1874[4]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1874[17]), 
          .C1(d_out_d_11__N_1874[5]), .D1(GND_net), .CIN(n11794), .COUT(n11795), 
          .S0(d_out_d_11__N_1876[5]), .S1(d_out_d_11__N_1876[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_453_9.INIT0 = 16'h6969;
    defparam add_453_9.INIT1 = 16'h6969;
    defparam add_453_9.INJECT1_0 = "NO";
    defparam add_453_9.INJECT1_1 = "NO";
    CCU2D add_453_7 (.A0(d_out_d_11__N_1874[2]), .B0(d_out_d_11__N_1874[17]), 
          .C0(GND_net), .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1874[17]), 
          .C1(d_out_d_11__N_1874[3]), .D1(GND_net), .CIN(n11793), .COUT(n11794), 
          .S0(d_out_d_11__N_1876[3]), .S1(d_out_d_11__N_1876[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_453_7.INIT0 = 16'h5999;
    defparam add_453_7.INIT1 = 16'h6969;
    defparam add_453_7.INJECT1_0 = "NO";
    defparam add_453_7.INJECT1_1 = "NO";
    CCU2D add_453_5 (.A0(d_out_d_11__N_1874[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1872[17]), .B1(d_out_d_11__N_1874[17]), 
          .C1(d_out_d_11__N_1874[1]), .D1(GND_net), .CIN(n11792), .COUT(n11793), 
          .S0(d_out_d_11__N_1876[1]), .S1(d_out_d_11__N_1876[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_453_5.INIT0 = 16'h5aaa;
    defparam add_453_5.INIT1 = 16'h9696;
    defparam add_453_5.INJECT1_0 = "NO";
    defparam add_453_5.INJECT1_1 = "NO";
    CCU2D add_453_3 (.A0(ISquare[18]), .B0(d_out_d_11__N_1874[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11791), .COUT(n11792), .S1(d_out_d_11__N_1876[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_453_3.INIT0 = 16'h5666;
    defparam add_453_3.INIT1 = 16'h5555;
    defparam add_453_3.INJECT1_0 = "NO";
    defparam add_453_3.INJECT1_1 = "NO";
    CCU2D add_3441_8 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n12451), 
          .S0(d_out_d_11__N_1872[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_3441_8.INIT0 = 16'h0fff;
    defparam add_3441_8.INIT1 = 16'h0000;
    defparam add_3441_8.INJECT1_0 = "NO";
    defparam add_3441_8.INJECT1_1 = "NO";
    CCU2D add_453_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1874[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n11791));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_453_1.INIT0 = 16'hF000;
    defparam add_453_1.INIT1 = 16'h0aaa;
    defparam add_453_1.INJECT1_0 = "NO";
    defparam add_453_1.INJECT1_1 = "NO";
    LUT4 mux_78_i1_3_lut (.A(d_out_d_11__N_2335[17]), .B(d_out_d_11__N_2353[17]), 
         .C(d_out_d_11__N_1892[17]), .Z(d_out_d_11__N_1894[17])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam mux_78_i1_3_lut.init = 16'h3535;
    CCU2D sub_78_add_2_18 (.A0(d_out_d_11__N_1892[14]), .B0(ISquare[31]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[15]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n11785), .S1(d_out_d_11__N_2335[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_18.INIT0 = 16'h5999;
    defparam sub_78_add_2_18.INIT1 = 16'h5555;
    defparam sub_78_add_2_18.INJECT1_0 = "NO";
    defparam sub_78_add_2_18.INJECT1_1 = "NO";
    FD1S3AX d_out_d__0_i2 (.D(d_out_d_11__N_1891), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[1]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i2.GSR = "ENABLED";
    CCU2D MultResult1_23__I_0_26 (.A0(MultResult1[23]), .B0(MultResult2[23]), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11244), .S0(ISquare_31__N_1895[24]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_26.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_26.INIT1 = 16'h0000;
    defparam MultResult1_23__I_0_26.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_26.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_24 (.A0(MultResult1[22]), .B0(MultResult2[22]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[23]), .B1(MultResult2[23]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11243), .COUT(n11244), .S0(ISquare_31__N_1895[22]), 
          .S1(ISquare_31__N_1895[23]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_24.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_24.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_24.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_24.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_22 (.A0(MultResult1[20]), .B0(MultResult2[20]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[21]), .B1(MultResult2[21]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11242), .COUT(n11243), .S0(ISquare_31__N_1895[20]), 
          .S1(ISquare_31__N_1895[21]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_22.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_22.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_22.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_22.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_20 (.A0(MultResult1[18]), .B0(MultResult2[18]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[19]), .B1(MultResult2[19]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11241), .COUT(n11242), .S0(ISquare_31__N_1895[18]), 
          .S1(ISquare_31__N_1895[19]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_20.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_20.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_20.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_20.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_18 (.A0(MultResult1[16]), .B0(MultResult2[16]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[17]), .B1(MultResult2[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11240), .COUT(n11241), .S0(ISquare_31__N_1895[16]), 
          .S1(ISquare_31__N_1895[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_18.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_18.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_18.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_18.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_16 (.A0(MultResult1[14]), .B0(MultResult2[14]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[15]), .B1(MultResult2[15]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11239), .COUT(n11240), .S0(ISquare_31__N_1895[14]), 
          .S1(ISquare_31__N_1895[15]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_16.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_16.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_16.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_16.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_14 (.A0(MultResult1[12]), .B0(MultResult2[12]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[13]), .B1(MultResult2[13]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11238), .COUT(n11239), .S0(ISquare_31__N_1895[12]), 
          .S1(ISquare_31__N_1895[13]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_14.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_14.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_14.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_14.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_12 (.A0(MultResult1[10]), .B0(MultResult2[10]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[11]), .B1(MultResult2[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11237), .COUT(n11238), .S0(ISquare_31__N_1895[10]), 
          .S1(ISquare_31__N_1895[11]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_12.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_12.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_12.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_12.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_10 (.A0(MultResult1[8]), .B0(MultResult2[8]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[9]), .B1(MultResult2[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11236), .COUT(n11237), .S0(ISquare_31__N_1895[8]), 
          .S1(ISquare_31__N_1895[9]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_10.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_10.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_10.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_10.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_8 (.A0(MultResult1[6]), .B0(MultResult2[6]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[7]), .B1(MultResult2[7]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11235), .COUT(n11236), .S0(ISquare_31__N_1895[6]), 
          .S1(ISquare_31__N_1895[7]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_8.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_8.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_8.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_8.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_6 (.A0(MultResult1[4]), .B0(MultResult2[4]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[5]), .B1(MultResult2[5]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11234), .COUT(n11235), .S0(ISquare_31__N_1895[4]), 
          .S1(ISquare_31__N_1895[5]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_6.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_6.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_6.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_6.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_4 (.A0(MultResult1[2]), .B0(MultResult2[2]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[3]), .B1(MultResult2[3]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11233), .COUT(n11234), .S0(ISquare_31__N_1895[2]), 
          .S1(ISquare_31__N_1895[3]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_4.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_4.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_4.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_4.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_2 (.A0(MultResult1[0]), .B0(MultResult2[0]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[1]), .B1(MultResult2[1]), 
          .C1(GND_net), .D1(GND_net), .COUT(n11233), .S1(ISquare_31__N_1895[1]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_2.INIT0 = 16'h7000;
    defparam MultResult1_23__I_0_2.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_2.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_2.INJECT1_1 = "NO";
    CCU2D add_513_11 (.A0(d_out_d_11__N_1872[17]), .B0(d_out_d_11__N_1871), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1872[17]), .B1(d_out_d_11__N_1871), 
          .C1(GND_net), .D1(GND_net), .CIN(n10995), .S0(d_out_d_11__N_1874[7]), 
          .S1(d_out_d_11__N_1874[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_513_11.INIT0 = 16'h5666;
    defparam add_513_11.INIT1 = 16'h5666;
    defparam add_513_11.INJECT1_0 = "NO";
    defparam add_513_11.INJECT1_1 = "NO";
    CCU2D add_513_9 (.A0(ISquare[31]), .B0(d_out_d_11__N_1872[17]), .C0(d_out_d_11__N_1872[4]), 
          .D0(GND_net), .A1(d_out_d_11__N_1872[5]), .B1(d_out_d_11__N_1872[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10994), .COUT(n10995), .S0(d_out_d_11__N_1874[5]), 
          .S1(d_out_d_11__N_1874[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_513_9.INIT0 = 16'h6969;
    defparam add_513_9.INIT1 = 16'h5999;
    defparam add_513_9.INJECT1_0 = "NO";
    defparam add_513_9.INJECT1_1 = "NO";
    CCU2D add_513_7 (.A0(ISquare[31]), .B0(d_out_d_11__N_1872[17]), .C0(d_out_d_11__N_1872[2]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1872[17]), 
          .C1(d_out_d_11__N_1872[3]), .D1(GND_net), .CIN(n10993), .COUT(n10994), 
          .S0(d_out_d_11__N_1874[3]), .S1(d_out_d_11__N_1874[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_513_7.INIT0 = 16'h6969;
    defparam add_513_7.INIT1 = 16'h6969;
    defparam add_513_7.INJECT1_0 = "NO";
    defparam add_513_7.INJECT1_1 = "NO";
    CCU2D add_513_5 (.A0(n12447), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1872[1]), .B1(d_out_d_11__N_1872[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10992), .COUT(n10993), .S0(d_out_d_11__N_1874[1]), 
          .S1(d_out_d_11__N_1874[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_513_5.INIT0 = 16'h5aaa;
    defparam add_513_5.INIT1 = 16'h5999;
    defparam add_513_5.INJECT1_0 = "NO";
    defparam add_513_5.INJECT1_1 = "NO";
    CCU2D add_513_3 (.A0(ISquare[20]), .B0(d_out_d_11__N_1872[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10991), .COUT(n10992), .S1(d_out_d_11__N_1874[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_513_3.INIT0 = 16'h5666;
    defparam add_513_3.INIT1 = 16'h5555;
    defparam add_513_3.INJECT1_0 = "NO";
    defparam add_513_3.INJECT1_1 = "NO";
    CCU2D add_513_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1872[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n10991));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_513_1.INIT0 = 16'hF000;
    defparam add_513_1.INIT1 = 16'h0aaa;
    defparam add_513_1.INJECT1_0 = "NO";
    defparam add_513_1.INJECT1_1 = "NO";
    FD1S3AX d_out_d__0_i3 (.D(d_out_d_11__N_1889), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i3.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i4 (.D(d_out_d_11__N_1887), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[3]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i4.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i5 (.D(d_out_d_11__N_1885), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i5.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i6 (.D(d_out_d_11__N_1883), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[5]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i6.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i7 (.D(d_out_d_11__N_1881), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i7.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i8 (.D(d_out_d_11__N_1879), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[7]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i8.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i9 (.D(d_out_d_11__N_1877), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i9.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i10 (.D(d_out_d_11__N_1875), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[9]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i10.GSR = "ENABLED";
    CCU2D add_3441_6 (.A0(n209), .B0(ISquare[31]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n12450), 
          .COUT(n12451), .S0(d_out_d_11__N_1872[4]), .S1(d_out_d_11__N_1872[5]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_3441_6.INIT0 = 16'h5666;
    defparam add_3441_6.INIT1 = 16'h0fff;
    defparam add_3441_6.INJECT1_0 = "NO";
    defparam add_3441_6.INJECT1_1 = "NO";
    CCU2D add_3441_4 (.A0(n209), .B0(ISquare[31]), .C0(GND_net), .D0(GND_net), 
          .A1(ISquare[31]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12449), .COUT(n12450), .S0(d_out_d_11__N_1872[2]), .S1(d_out_d_11__N_1872[3]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_3441_4.INIT0 = 16'h5666;
    defparam add_3441_4.INIT1 = 16'h0555;
    defparam add_3441_4.INJECT1_0 = "NO";
    defparam add_3441_4.INJECT1_1 = "NO";
    CCU2D add_3441_2 (.A0(ISquare[23]), .B0(ISquare[22]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n12449), .S1(d_out_d_11__N_1872[1]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_3441_2.INIT0 = 16'h1000;
    defparam add_3441_2.INIT1 = 16'h0fff;
    defparam add_3441_2.INJECT1_0 = "NO";
    defparam add_3441_2.INJECT1_1 = "NO";
    CCU2D add_413_17 (.A0(d_out_d_11__N_1878[17]), .B0(d_out_d_11__N_1877), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1878[17]), .B1(d_out_d_11__N_1877), 
          .C1(GND_net), .D1(GND_net), .CIN(n12445), .S0(d_out_d_11__N_1880[13]), 
          .S1(d_out_d_11__N_1880[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_413_17.INIT0 = 16'h5666;
    defparam add_413_17.INIT1 = 16'h5666;
    defparam add_413_17.INJECT1_0 = "NO";
    defparam add_413_17.INJECT1_1 = "NO";
    CCU2D add_413_15 (.A0(d_out_d_11__N_1878[10]), .B0(d_out_d_11__N_1878[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1878[11]), .B1(d_out_d_11__N_1878[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12444), .COUT(n12445), .S0(d_out_d_11__N_1880[11]), 
          .S1(d_out_d_11__N_1880[12]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_413_15.INIT0 = 16'h5999;
    defparam add_413_15.INIT1 = 16'h5999;
    defparam add_413_15.INJECT1_0 = "NO";
    defparam add_413_15.INJECT1_1 = "NO";
    CCU2D add_413_13 (.A0(d_out_d_11__N_1878[8]), .B0(d_out_d_11__N_1878[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1878[9]), .B1(d_out_d_11__N_1878[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12443), .COUT(n12444), .S0(d_out_d_11__N_1880[9]), 
          .S1(d_out_d_11__N_1880[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_413_13.INIT0 = 16'h5999;
    defparam add_413_13.INIT1 = 16'h5999;
    defparam add_413_13.INJECT1_0 = "NO";
    defparam add_413_13.INJECT1_1 = "NO";
    CCU2D add_413_11 (.A0(ISquare[31]), .B0(d_out_d_11__N_1878[17]), .C0(d_out_d_11__N_1878[6]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1878[17]), 
          .C1(d_out_d_11__N_1878[7]), .D1(GND_net), .CIN(n12442), .COUT(n12443), 
          .S0(d_out_d_11__N_1880[7]), .S1(d_out_d_11__N_1880[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_413_11.INIT0 = 16'h6969;
    defparam add_413_11.INIT1 = 16'h6969;
    defparam add_413_11.INJECT1_0 = "NO";
    defparam add_413_11.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_16 (.A0(d_out_d_11__N_1892[12]), .B0(ISquare[31]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[13]), .B1(ISquare[31]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11784), .COUT(n11785));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_16.INIT0 = 16'h5999;
    defparam sub_78_add_2_16.INIT1 = 16'h5999;
    defparam sub_78_add_2_16.INJECT1_0 = "NO";
    defparam sub_78_add_2_16.INJECT1_1 = "NO";
    CCU2D add_413_9 (.A0(d_out_d_11__N_1878[4]), .B0(d_out_d_11__N_1878[17]), 
          .C0(GND_net), .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1878[17]), 
          .C1(d_out_d_11__N_1878[5]), .D1(GND_net), .CIN(n12441), .COUT(n12442), 
          .S0(d_out_d_11__N_1880[5]), .S1(d_out_d_11__N_1880[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_413_9.INIT0 = 16'h5999;
    defparam add_413_9.INIT1 = 16'h6969;
    defparam add_413_9.INJECT1_0 = "NO";
    defparam add_413_9.INJECT1_1 = "NO";
    CCU2D add_413_7 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1878[17]), 
          .C0(d_out_d_11__N_1878[2]), .D0(GND_net), .A1(d_out_d_11__N_1872[17]), 
          .B1(d_out_d_11__N_1878[17]), .C1(d_out_d_11__N_1878[3]), .D1(GND_net), 
          .CIN(n12440), .COUT(n12441), .S0(d_out_d_11__N_1880[3]), .S1(d_out_d_11__N_1880[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_413_7.INIT0 = 16'h9696;
    defparam add_413_7.INIT1 = 16'h9696;
    defparam add_413_7.INJECT1_0 = "NO";
    defparam add_413_7.INJECT1_1 = "NO";
    CCU2D add_413_5 (.A0(d_out_d_11__N_1878[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1876[17]), .B1(d_out_d_11__N_1878[17]), 
          .C1(d_out_d_11__N_1878[1]), .D1(GND_net), .CIN(n12439), .COUT(n12440), 
          .S0(d_out_d_11__N_1880[1]), .S1(d_out_d_11__N_1880[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_413_5.INIT0 = 16'h5aaa;
    defparam add_413_5.INIT1 = 16'h9696;
    defparam add_413_5.INJECT1_0 = "NO";
    defparam add_413_5.INJECT1_1 = "NO";
    CCU2D add_413_3 (.A0(ISquare[14]), .B0(d_out_d_11__N_1878[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12438), .COUT(n12439), .S1(d_out_d_11__N_1880[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_413_3.INIT0 = 16'h5666;
    defparam add_413_3.INIT1 = 16'h5555;
    defparam add_413_3.INJECT1_0 = "NO";
    defparam add_413_3.INJECT1_1 = "NO";
    CCU2D add_413_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1878[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n12438));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_413_1.INIT0 = 16'hF000;
    defparam add_413_1.INIT1 = 16'h0aaa;
    defparam add_413_1.INJECT1_0 = "NO";
    defparam add_413_1.INJECT1_1 = "NO";
    CCU2D add_140_17 (.A0(d_out_d_11__N_1892[14]), .B0(ISquare[31]), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1892[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12432), .S1(d_out_d_11__N_2353[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_140_17.INIT0 = 16'h5666;
    defparam add_140_17.INIT1 = 16'h5aaa;
    defparam add_140_17.INJECT1_0 = "NO";
    defparam add_140_17.INJECT1_1 = "NO";
    CCU2D add_140_15 (.A0(d_out_d_11__N_1892[12]), .B0(ISquare[31]), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1892[13]), .B1(ISquare[31]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12431), .COUT(n12432));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_140_15.INIT0 = 16'h5666;
    defparam add_140_15.INIT1 = 16'h5666;
    defparam add_140_15.INJECT1_0 = "NO";
    defparam add_140_15.INJECT1_1 = "NO";
    CCU2D add_140_13 (.A0(d_out_d_11__N_1892[10]), .B0(d_out_d_11__N_1872[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[11]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12430), .COUT(n12431));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_140_13.INIT0 = 16'h5999;
    defparam add_140_13.INIT1 = 16'h5aaa;
    defparam add_140_13.INJECT1_0 = "NO";
    defparam add_140_13.INJECT1_1 = "NO";
    CCU2D add_140_11 (.A0(d_out_d_11__N_1892[8]), .B0(d_out_d_11__N_1876[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[9]), .B1(d_out_d_11__N_1874[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12429), .COUT(n12430));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_140_11.INIT0 = 16'h5999;
    defparam add_140_11.INIT1 = 16'h5999;
    defparam add_140_11.INJECT1_0 = "NO";
    defparam add_140_11.INJECT1_1 = "NO";
    CCU2D add_140_9 (.A0(d_out_d_11__N_1892[6]), .B0(d_out_d_11__N_1880[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[7]), .B1(d_out_d_11__N_1878[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12428), .COUT(n12429));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_140_9.INIT0 = 16'h5999;
    defparam add_140_9.INIT1 = 16'h5999;
    defparam add_140_9.INJECT1_0 = "NO";
    defparam add_140_9.INJECT1_1 = "NO";
    CCU2D add_140_7 (.A0(d_out_d_11__N_1892[4]), .B0(d_out_d_11__N_1884[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[5]), .B1(d_out_d_11__N_1882[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12427), .COUT(n12428));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_140_7.INIT0 = 16'h5999;
    defparam add_140_7.INIT1 = 16'h5999;
    defparam add_140_7.INJECT1_0 = "NO";
    defparam add_140_7.INJECT1_1 = "NO";
    CCU2D add_140_5 (.A0(d_out_d_11__N_1892[2]), .B0(d_out_d_11__N_1888[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[3]), .B1(d_out_d_11__N_1886[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12426), .COUT(n12427));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_140_5.INIT0 = 16'h5999;
    defparam add_140_5.INIT1 = 16'h5999;
    defparam add_140_5.INJECT1_0 = "NO";
    defparam add_140_5.INJECT1_1 = "NO";
    CCU2D add_140_3 (.A0(d_out_d_11__N_1892[0]), .B0(d_out_d_11__N_1892[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[1]), .B1(d_out_d_11__N_1890[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12425), .COUT(n12426));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_140_3.INIT0 = 16'h5999;
    defparam add_140_3.INIT1 = 16'h5999;
    defparam add_140_3.INJECT1_0 = "NO";
    defparam add_140_3.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_14 (.A0(d_out_d_11__N_1892[10]), .B0(d_out_d_11__N_1872[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[11]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n11783), .COUT(n11784));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_14.INIT0 = 16'h5666;
    defparam sub_78_add_2_14.INIT1 = 16'h5555;
    defparam sub_78_add_2_14.INJECT1_0 = "NO";
    defparam sub_78_add_2_14.INJECT1_1 = "NO";
    CCU2D add_140_1 (.A0(ISquare[0]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(ISquare[1]), .B1(d_out_d_11__N_1892[17]), .C1(GND_net), 
          .D1(GND_net), .COUT(n12425));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_140_1.INIT0 = 16'h5000;
    defparam add_140_1.INIT1 = 16'h5666;
    defparam add_140_1.INJECT1_0 = "NO";
    defparam add_140_1.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_12 (.A0(d_out_d_11__N_1892[8]), .B0(d_out_d_11__N_1876[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[9]), .B1(d_out_d_11__N_1874[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11782), .COUT(n11783));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_12.INIT0 = 16'h5666;
    defparam sub_78_add_2_12.INIT1 = 16'h5666;
    defparam sub_78_add_2_12.INJECT1_0 = "NO";
    defparam sub_78_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_10 (.A0(d_out_d_11__N_1892[6]), .B0(d_out_d_11__N_1880[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[7]), .B1(d_out_d_11__N_1878[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11781), .COUT(n11782));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_10.INIT0 = 16'h5666;
    defparam sub_78_add_2_10.INIT1 = 16'h5666;
    defparam sub_78_add_2_10.INJECT1_0 = "NO";
    defparam sub_78_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_8 (.A0(d_out_d_11__N_1892[4]), .B0(d_out_d_11__N_1884[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[5]), .B1(d_out_d_11__N_1882[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11780), .COUT(n11781));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_8.INIT0 = 16'h5666;
    defparam sub_78_add_2_8.INIT1 = 16'h5666;
    defparam sub_78_add_2_8.INJECT1_0 = "NO";
    defparam sub_78_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_6 (.A0(d_out_d_11__N_1892[2]), .B0(d_out_d_11__N_1888[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[3]), .B1(d_out_d_11__N_1886[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11779), .COUT(n11780));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_6.INIT0 = 16'h5666;
    defparam sub_78_add_2_6.INIT1 = 16'h5666;
    defparam sub_78_add_2_6.INJECT1_0 = "NO";
    defparam sub_78_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_4 (.A0(d_out_d_11__N_1892[0]), .B0(d_out_d_11__N_1892[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1892[1]), .B1(d_out_d_11__N_1890[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11778), .COUT(n11779));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_4.INIT0 = 16'h5666;
    defparam sub_78_add_2_4.INIT1 = 16'h5666;
    defparam sub_78_add_2_4.INJECT1_0 = "NO";
    defparam sub_78_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_2 (.A0(ISquare[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[1]), .B1(d_out_d_11__N_1892[17]), 
          .C1(GND_net), .D1(GND_net), .COUT(n11778));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_2.INIT0 = 16'h5000;
    defparam sub_78_add_2_2.INIT1 = 16'h5999;
    defparam sub_78_add_2_2.INJECT1_0 = "NO";
    defparam sub_78_add_2_2.INJECT1_1 = "NO";
    CCU2D add_573_19 (.A0(d_out_d_11__N_1886[14]), .B0(d_out_d_11__N_1886[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1886[15]), .B1(d_out_d_11__N_1886[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11758), .S0(d_out_d_11__N_1888[15]), 
          .S1(d_out_d_11__N_1888[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_573_19.INIT0 = 16'h5999;
    defparam add_573_19.INIT1 = 16'h5999;
    defparam add_573_19.INJECT1_0 = "NO";
    defparam add_573_19.INJECT1_1 = "NO";
    CCU2D add_573_17 (.A0(d_out_d_11__N_1886[12]), .B0(d_out_d_11__N_1886[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1886[13]), .B1(d_out_d_11__N_1886[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11757), .COUT(n11758), .S0(d_out_d_11__N_1888[13]), 
          .S1(d_out_d_11__N_1888[14]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_573_17.INIT0 = 16'h5999;
    defparam add_573_17.INIT1 = 16'h5999;
    defparam add_573_17.INJECT1_0 = "NO";
    defparam add_573_17.INJECT1_1 = "NO";
    CCU2D add_573_15 (.A0(ISquare[31]), .B0(d_out_d_11__N_1886[17]), .C0(d_out_d_11__N_1886[10]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1886[17]), 
          .C1(d_out_d_11__N_1886[11]), .D1(GND_net), .CIN(n11756), .COUT(n11757), 
          .S0(d_out_d_11__N_1888[11]), .S1(d_out_d_11__N_1888[12]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_573_15.INIT0 = 16'h6969;
    defparam add_573_15.INIT1 = 16'h6969;
    defparam add_573_15.INJECT1_0 = "NO";
    defparam add_573_15.INJECT1_1 = "NO";
    CCU2D add_573_13 (.A0(d_out_d_11__N_1886[8]), .B0(d_out_d_11__N_1886[17]), 
          .C0(GND_net), .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1886[17]), 
          .C1(d_out_d_11__N_1886[9]), .D1(GND_net), .CIN(n11755), .COUT(n11756), 
          .S0(d_out_d_11__N_1888[9]), .S1(d_out_d_11__N_1888[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_573_13.INIT0 = 16'h5999;
    defparam add_573_13.INIT1 = 16'h6969;
    defparam add_573_13.INJECT1_0 = "NO";
    defparam add_573_13.INJECT1_1 = "NO";
    CCU2D add_573_11 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1886[17]), 
          .C0(d_out_d_11__N_1886[6]), .D0(GND_net), .A1(d_out_d_11__N_1872[17]), 
          .B1(d_out_d_11__N_1886[17]), .C1(d_out_d_11__N_1886[7]), .D1(GND_net), 
          .CIN(n11754), .COUT(n11755), .S0(d_out_d_11__N_1888[7]), .S1(d_out_d_11__N_1888[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_573_11.INIT0 = 16'h9696;
    defparam add_573_11.INIT1 = 16'h9696;
    defparam add_573_11.INJECT1_0 = "NO";
    defparam add_573_11.INJECT1_1 = "NO";
    CCU2D add_573_9 (.A0(d_out_d_11__N_1878[17]), .B0(d_out_d_11__N_1886[17]), 
          .C0(d_out_d_11__N_1886[4]), .D0(GND_net), .A1(d_out_d_11__N_1876[17]), 
          .B1(d_out_d_11__N_1886[17]), .C1(d_out_d_11__N_1886[5]), .D1(GND_net), 
          .CIN(n11753), .COUT(n11754), .S0(d_out_d_11__N_1888[5]), .S1(d_out_d_11__N_1888[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_573_9.INIT0 = 16'h9696;
    defparam add_573_9.INIT1 = 16'h9696;
    defparam add_573_9.INJECT1_0 = "NO";
    defparam add_573_9.INJECT1_1 = "NO";
    CCU2D add_573_7 (.A0(d_out_d_11__N_1882[17]), .B0(d_out_d_11__N_1886[17]), 
          .C0(d_out_d_11__N_1886[2]), .D0(GND_net), .A1(d_out_d_11__N_1880[17]), 
          .B1(d_out_d_11__N_1886[17]), .C1(d_out_d_11__N_1886[3]), .D1(GND_net), 
          .CIN(n11752), .COUT(n11753), .S0(d_out_d_11__N_1888[3]), .S1(d_out_d_11__N_1888[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_573_7.INIT0 = 16'h9696;
    defparam add_573_7.INIT1 = 16'h9696;
    defparam add_573_7.INJECT1_0 = "NO";
    defparam add_573_7.INJECT1_1 = "NO";
    CCU2D add_573_5 (.A0(d_out_d_11__N_1886[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1884[17]), .B1(d_out_d_11__N_1886[17]), 
          .C1(d_out_d_11__N_1886[1]), .D1(GND_net), .CIN(n11751), .COUT(n11752), 
          .S0(d_out_d_11__N_1888[1]), .S1(d_out_d_11__N_1888[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_573_5.INIT0 = 16'h5aaa;
    defparam add_573_5.INIT1 = 16'h9696;
    defparam add_573_5.INJECT1_0 = "NO";
    defparam add_573_5.INJECT1_1 = "NO";
    CCU2D add_573_3 (.A0(ISquare[6]), .B0(d_out_d_11__N_1886[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11750), .COUT(n11751), .S1(d_out_d_11__N_1888[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_573_3.INIT0 = 16'h5666;
    defparam add_573_3.INIT1 = 16'h5555;
    defparam add_573_3.INJECT1_0 = "NO";
    defparam add_573_3.INJECT1_1 = "NO";
    CCU2D add_573_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1886[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n11750));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_573_1.INIT0 = 16'hF000;
    defparam add_573_1.INIT1 = 16'h0aaa;
    defparam add_573_1.INJECT1_0 = "NO";
    defparam add_573_1.INJECT1_1 = "NO";
    CCU2D add_493_19 (.A0(d_out_d_11__N_1880[17]), .B0(d_out_d_11__N_1879), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1880[17]), .B1(d_out_d_11__N_1879), 
          .C1(GND_net), .D1(GND_net), .CIN(n11654), .S0(d_out_d_11__N_1882[15]), 
          .S1(d_out_d_11__N_1882[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_493_19.INIT0 = 16'h5666;
    defparam add_493_19.INIT1 = 16'h5666;
    defparam add_493_19.INJECT1_0 = "NO";
    defparam add_493_19.INJECT1_1 = "NO";
    CCU2D add_493_17 (.A0(d_out_d_11__N_1880[12]), .B0(d_out_d_11__N_1880[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1880[13]), .B1(d_out_d_11__N_1880[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11653), .COUT(n11654), .S0(d_out_d_11__N_1882[13]), 
          .S1(d_out_d_11__N_1882[14]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_493_17.INIT0 = 16'h5999;
    defparam add_493_17.INIT1 = 16'h5999;
    defparam add_493_17.INJECT1_0 = "NO";
    defparam add_493_17.INJECT1_1 = "NO";
    CCU2D add_493_15 (.A0(d_out_d_11__N_1880[10]), .B0(d_out_d_11__N_1880[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1880[11]), .B1(d_out_d_11__N_1880[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11652), .COUT(n11653), .S0(d_out_d_11__N_1882[11]), 
          .S1(d_out_d_11__N_1882[12]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_493_15.INIT0 = 16'h5999;
    defparam add_493_15.INIT1 = 16'h5999;
    defparam add_493_15.INJECT1_0 = "NO";
    defparam add_493_15.INJECT1_1 = "NO";
    CCU2D add_493_13 (.A0(ISquare[31]), .B0(d_out_d_11__N_1880[17]), .C0(d_out_d_11__N_1880[8]), 
          .D0(GND_net), .A1(d_out_d_11__N_1880[9]), .B1(d_out_d_11__N_1880[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11651), .COUT(n11652), .S0(d_out_d_11__N_1882[9]), 
          .S1(d_out_d_11__N_1882[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_493_13.INIT0 = 16'h6969;
    defparam add_493_13.INIT1 = 16'h5999;
    defparam add_493_13.INJECT1_0 = "NO";
    defparam add_493_13.INJECT1_1 = "NO";
    CCU2D add_493_11 (.A0(ISquare[31]), .B0(d_out_d_11__N_1880[17]), .C0(d_out_d_11__N_1880[6]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1880[17]), 
          .C1(d_out_d_11__N_1880[7]), .D1(GND_net), .CIN(n11650), .COUT(n11651), 
          .S0(d_out_d_11__N_1882[7]), .S1(d_out_d_11__N_1882[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_493_11.INIT0 = 16'h6969;
    defparam add_493_11.INIT1 = 16'h6969;
    defparam add_493_11.INJECT1_0 = "NO";
    defparam add_493_11.INJECT1_1 = "NO";
    CCU2D add_493_9 (.A0(d_out_d_11__N_1872[17]), .B0(d_out_d_11__N_1880[17]), 
          .C0(d_out_d_11__N_1880[4]), .D0(GND_net), .A1(d_out_d_11__N_1880[5]), 
          .B1(d_out_d_11__N_1880[17]), .C1(GND_net), .D1(GND_net), .CIN(n11649), 
          .COUT(n11650), .S0(d_out_d_11__N_1882[5]), .S1(d_out_d_11__N_1882[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_493_9.INIT0 = 16'h9696;
    defparam add_493_9.INIT1 = 16'h5999;
    defparam add_493_9.INJECT1_0 = "NO";
    defparam add_493_9.INJECT1_1 = "NO";
    CCU2D add_493_7 (.A0(d_out_d_11__N_1876[17]), .B0(d_out_d_11__N_1880[17]), 
          .C0(d_out_d_11__N_1880[2]), .D0(GND_net), .A1(d_out_d_11__N_1874[17]), 
          .B1(d_out_d_11__N_1880[17]), .C1(d_out_d_11__N_1880[3]), .D1(GND_net), 
          .CIN(n11648), .COUT(n11649), .S0(d_out_d_11__N_1882[3]), .S1(d_out_d_11__N_1882[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_493_7.INIT0 = 16'h9696;
    defparam add_493_7.INIT1 = 16'h9696;
    defparam add_493_7.INJECT1_0 = "NO";
    defparam add_493_7.INJECT1_1 = "NO";
    CCU2D add_493_5 (.A0(d_out_d_11__N_1880[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1878[17]), .B1(d_out_d_11__N_1880[17]), 
          .C1(d_out_d_11__N_1880[1]), .D1(GND_net), .CIN(n11647), .COUT(n11648), 
          .S0(d_out_d_11__N_1882[1]), .S1(d_out_d_11__N_1882[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_493_5.INIT0 = 16'h5aaa;
    defparam add_493_5.INIT1 = 16'h9696;
    defparam add_493_5.INJECT1_0 = "NO";
    defparam add_493_5.INJECT1_1 = "NO";
    CCU2D add_493_3 (.A0(ISquare[12]), .B0(d_out_d_11__N_1880[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11646), .COUT(n11647), .S1(d_out_d_11__N_1882[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_493_3.INIT0 = 16'h5666;
    defparam add_493_3.INIT1 = 16'h5555;
    defparam add_493_3.INJECT1_0 = "NO";
    defparam add_493_3.INJECT1_1 = "NO";
    CCU2D add_493_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1880[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n11646));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_493_1.INIT0 = 16'hF000;
    defparam add_493_1.INIT1 = 16'h0aaa;
    defparam add_493_1.INJECT1_0 = "NO";
    defparam add_493_1.INJECT1_1 = "NO";
    CCU2D add_613_19 (.A0(d_out_d_11__N_1884[14]), .B0(d_out_d_11__N_1884[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1884[15]), .B1(d_out_d_11__N_1884[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12397), .S0(d_out_d_11__N_1886[15]), 
          .S1(d_out_d_11__N_1886[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_613_19.INIT0 = 16'h5999;
    defparam add_613_19.INIT1 = 16'h5999;
    defparam add_613_19.INJECT1_0 = "NO";
    defparam add_613_19.INJECT1_1 = "NO";
    CCU2D add_613_17 (.A0(d_out_d_11__N_1884[12]), .B0(d_out_d_11__N_1884[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1884[13]), .B1(d_out_d_11__N_1884[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12396), .COUT(n12397), .S0(d_out_d_11__N_1886[13]), 
          .S1(d_out_d_11__N_1886[14]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_613_17.INIT0 = 16'h5999;
    defparam add_613_17.INIT1 = 16'h5999;
    defparam add_613_17.INJECT1_0 = "NO";
    defparam add_613_17.INJECT1_1 = "NO";
    CCU2D add_613_15 (.A0(ISquare[31]), .B0(d_out_d_11__N_1884[17]), .C0(d_out_d_11__N_1884[10]), 
          .D0(GND_net), .A1(d_out_d_11__N_1884[11]), .B1(d_out_d_11__N_1884[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12395), .COUT(n12396), .S0(d_out_d_11__N_1886[11]), 
          .S1(d_out_d_11__N_1886[12]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_613_15.INIT0 = 16'h6969;
    defparam add_613_15.INIT1 = 16'h5999;
    defparam add_613_15.INJECT1_0 = "NO";
    defparam add_613_15.INJECT1_1 = "NO";
    CCU2D add_613_13 (.A0(ISquare[31]), .B0(d_out_d_11__N_1884[17]), .C0(d_out_d_11__N_1884[8]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1884[17]), 
          .C1(d_out_d_11__N_1884[9]), .D1(GND_net), .CIN(n12394), .COUT(n12395), 
          .S0(d_out_d_11__N_1886[9]), .S1(d_out_d_11__N_1886[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_613_13.INIT0 = 16'h6969;
    defparam add_613_13.INIT1 = 16'h6969;
    defparam add_613_13.INJECT1_0 = "NO";
    defparam add_613_13.INJECT1_1 = "NO";
    CCU2D add_613_11 (.A0(d_out_d_11__N_1872[17]), .B0(d_out_d_11__N_1884[17]), 
          .C0(d_out_d_11__N_1884[6]), .D0(GND_net), .A1(d_out_d_11__N_1884[7]), 
          .B1(d_out_d_11__N_1884[17]), .C1(GND_net), .D1(GND_net), .CIN(n12393), 
          .COUT(n12394), .S0(d_out_d_11__N_1886[7]), .S1(d_out_d_11__N_1886[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_613_11.INIT0 = 16'h9696;
    defparam add_613_11.INIT1 = 16'h5999;
    defparam add_613_11.INJECT1_0 = "NO";
    defparam add_613_11.INJECT1_1 = "NO";
    CCU2D add_613_9 (.A0(d_out_d_11__N_1876[17]), .B0(d_out_d_11__N_1884[17]), 
          .C0(d_out_d_11__N_1884[4]), .D0(GND_net), .A1(d_out_d_11__N_1874[17]), 
          .B1(d_out_d_11__N_1884[17]), .C1(d_out_d_11__N_1884[5]), .D1(GND_net), 
          .CIN(n12392), .COUT(n12393), .S0(d_out_d_11__N_1886[5]), .S1(d_out_d_11__N_1886[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_613_9.INIT0 = 16'h9696;
    defparam add_613_9.INIT1 = 16'h9696;
    defparam add_613_9.INJECT1_0 = "NO";
    defparam add_613_9.INJECT1_1 = "NO";
    CCU2D add_613_7 (.A0(d_out_d_11__N_1880[17]), .B0(d_out_d_11__N_1884[17]), 
          .C0(d_out_d_11__N_1884[2]), .D0(GND_net), .A1(d_out_d_11__N_1878[17]), 
          .B1(d_out_d_11__N_1884[17]), .C1(d_out_d_11__N_1884[3]), .D1(GND_net), 
          .CIN(n12391), .COUT(n12392), .S0(d_out_d_11__N_1886[3]), .S1(d_out_d_11__N_1886[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_613_7.INIT0 = 16'h9696;
    defparam add_613_7.INIT1 = 16'h9696;
    defparam add_613_7.INJECT1_0 = "NO";
    defparam add_613_7.INJECT1_1 = "NO";
    CCU2D add_613_5 (.A0(d_out_d_11__N_1884[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1882[17]), .B1(d_out_d_11__N_1884[17]), 
          .C1(d_out_d_11__N_1884[1]), .D1(GND_net), .CIN(n12390), .COUT(n12391), 
          .S0(d_out_d_11__N_1886[1]), .S1(d_out_d_11__N_1886[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_613_5.INIT0 = 16'h5aaa;
    defparam add_613_5.INIT1 = 16'h9696;
    defparam add_613_5.INJECT1_0 = "NO";
    defparam add_613_5.INJECT1_1 = "NO";
    CCU2D add_613_3 (.A0(ISquare[8]), .B0(d_out_d_11__N_1884[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12389), .COUT(n12390), .S1(d_out_d_11__N_1886[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_613_3.INIT0 = 16'h5666;
    defparam add_613_3.INIT1 = 16'h5555;
    defparam add_613_3.INJECT1_0 = "NO";
    defparam add_613_3.INJECT1_1 = "NO";
    CCU2D add_613_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1884[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n12389));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_613_1.INIT0 = 16'hF000;
    defparam add_613_1.INIT1 = 16'h0aaa;
    defparam add_613_1.INJECT1_0 = "NO";
    defparam add_613_1.INJECT1_1 = "NO";
    CCU2D add_653_19 (.A0(d_out_d_11__N_1882[14]), .B0(d_out_d_11__N_1882[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1882[15]), .B1(d_out_d_11__N_1882[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12383), .S0(d_out_d_11__N_1884[15]), 
          .S1(d_out_d_11__N_1884[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_653_19.INIT0 = 16'h5999;
    defparam add_653_19.INIT1 = 16'h5999;
    defparam add_653_19.INJECT1_0 = "NO";
    defparam add_653_19.INJECT1_1 = "NO";
    CCU2D add_653_17 (.A0(d_out_d_11__N_1882[12]), .B0(d_out_d_11__N_1882[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1882[13]), .B1(d_out_d_11__N_1882[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12382), .COUT(n12383), .S0(d_out_d_11__N_1884[13]), 
          .S1(d_out_d_11__N_1884[14]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_653_17.INIT0 = 16'h5999;
    defparam add_653_17.INIT1 = 16'h5999;
    defparam add_653_17.INJECT1_0 = "NO";
    defparam add_653_17.INJECT1_1 = "NO";
    CCU2D add_653_15 (.A0(d_out_d_11__N_1882[10]), .B0(d_out_d_11__N_1882[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1882[11]), .B1(d_out_d_11__N_1882[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12381), .COUT(n12382), .S0(d_out_d_11__N_1884[11]), 
          .S1(d_out_d_11__N_1884[12]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_653_15.INIT0 = 16'h5999;
    defparam add_653_15.INIT1 = 16'h5999;
    defparam add_653_15.INJECT1_0 = "NO";
    defparam add_653_15.INJECT1_1 = "NO";
    CCU2D add_653_13 (.A0(ISquare[31]), .B0(d_out_d_11__N_1882[17]), .C0(d_out_d_11__N_1882[8]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1882[17]), 
          .C1(d_out_d_11__N_1882[9]), .D1(GND_net), .CIN(n12380), .COUT(n12381), 
          .S0(d_out_d_11__N_1884[9]), .S1(d_out_d_11__N_1884[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_653_13.INIT0 = 16'h6969;
    defparam add_653_13.INIT1 = 16'h6969;
    defparam add_653_13.INJECT1_0 = "NO";
    defparam add_653_13.INJECT1_1 = "NO";
    CCU2D add_653_11 (.A0(d_out_d_11__N_1882[6]), .B0(d_out_d_11__N_1882[17]), 
          .C0(GND_net), .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1882[17]), 
          .C1(d_out_d_11__N_1882[7]), .D1(GND_net), .CIN(n12379), .COUT(n12380), 
          .S0(d_out_d_11__N_1884[7]), .S1(d_out_d_11__N_1884[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_653_11.INIT0 = 16'h5999;
    defparam add_653_11.INIT1 = 16'h6969;
    defparam add_653_11.INJECT1_0 = "NO";
    defparam add_653_11.INJECT1_1 = "NO";
    CCU2D add_653_9 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1882[17]), 
          .C0(d_out_d_11__N_1882[4]), .D0(GND_net), .A1(d_out_d_11__N_1872[17]), 
          .B1(d_out_d_11__N_1882[17]), .C1(d_out_d_11__N_1882[5]), .D1(GND_net), 
          .CIN(n12378), .COUT(n12379), .S0(d_out_d_11__N_1884[5]), .S1(d_out_d_11__N_1884[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_653_9.INIT0 = 16'h9696;
    defparam add_653_9.INIT1 = 16'h9696;
    defparam add_653_9.INJECT1_0 = "NO";
    defparam add_653_9.INJECT1_1 = "NO";
    CCU2D add_653_7 (.A0(d_out_d_11__N_1878[17]), .B0(d_out_d_11__N_1882[17]), 
          .C0(d_out_d_11__N_1882[2]), .D0(GND_net), .A1(d_out_d_11__N_1876[17]), 
          .B1(d_out_d_11__N_1882[17]), .C1(d_out_d_11__N_1882[3]), .D1(GND_net), 
          .CIN(n12377), .COUT(n12378), .S0(d_out_d_11__N_1884[3]), .S1(d_out_d_11__N_1884[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_653_7.INIT0 = 16'h9696;
    defparam add_653_7.INIT1 = 16'h9696;
    defparam add_653_7.INJECT1_0 = "NO";
    defparam add_653_7.INJECT1_1 = "NO";
    CCU2D add_653_5 (.A0(d_out_d_11__N_1882[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1880[17]), .B1(d_out_d_11__N_1882[17]), 
          .C1(d_out_d_11__N_1882[1]), .D1(GND_net), .CIN(n12376), .COUT(n12377), 
          .S0(d_out_d_11__N_1884[1]), .S1(d_out_d_11__N_1884[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_653_5.INIT0 = 16'h5aaa;
    defparam add_653_5.INIT1 = 16'h9696;
    defparam add_653_5.INJECT1_0 = "NO";
    defparam add_653_5.INJECT1_1 = "NO";
    CCU2D add_653_3 (.A0(ISquare[10]), .B0(d_out_d_11__N_1882[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12375), .COUT(n12376), .S1(d_out_d_11__N_1884[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_653_3.INIT0 = 16'h5666;
    defparam add_653_3.INIT1 = 16'h5555;
    defparam add_653_3.INJECT1_0 = "NO";
    defparam add_653_3.INJECT1_1 = "NO";
    CCU2D add_653_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1882[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n12375));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_653_1.INIT0 = 16'hF000;
    defparam add_653_1.INIT1 = 16'h0aaa;
    defparam add_653_1.INJECT1_0 = "NO";
    defparam add_653_1.INJECT1_1 = "NO";
    CCU2D add_533_19 (.A0(d_out_d_11__N_1890[14]), .B0(d_out_d_11__N_1890[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1890[15]), .B1(d_out_d_11__N_1890[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12369), .S0(d_out_d_11__N_1892[15]), 
          .S1(d_out_d_11__N_1892[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_533_19.INIT0 = 16'h5999;
    defparam add_533_19.INIT1 = 16'h5999;
    defparam add_533_19.INJECT1_0 = "NO";
    defparam add_533_19.INJECT1_1 = "NO";
    CCU2D add_533_17 (.A0(ISquare[31]), .B0(d_out_d_11__N_1890[17]), .C0(d_out_d_11__N_1890[12]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1890[17]), 
          .C1(d_out_d_11__N_1890[13]), .D1(GND_net), .CIN(n12368), .COUT(n12369), 
          .S0(d_out_d_11__N_1892[13]), .S1(d_out_d_11__N_1892[14]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_533_17.INIT0 = 16'h6969;
    defparam add_533_17.INIT1 = 16'h6969;
    defparam add_533_17.INJECT1_0 = "NO";
    defparam add_533_17.INJECT1_1 = "NO";
    CCU2D add_533_15 (.A0(d_out_d_11__N_1890[10]), .B0(d_out_d_11__N_1890[17]), 
          .C0(GND_net), .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1890[17]), 
          .C1(d_out_d_11__N_1890[11]), .D1(GND_net), .CIN(n12367), .COUT(n12368), 
          .S0(d_out_d_11__N_1892[11]), .S1(d_out_d_11__N_1892[12]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_533_15.INIT0 = 16'h5999;
    defparam add_533_15.INIT1 = 16'h6969;
    defparam add_533_15.INJECT1_0 = "NO";
    defparam add_533_15.INJECT1_1 = "NO";
    CCU2D add_533_13 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(d_out_d_11__N_1890[8]), .D0(GND_net), .A1(d_out_d_11__N_1872[17]), 
          .B1(d_out_d_11__N_1890[17]), .C1(d_out_d_11__N_1890[9]), .D1(GND_net), 
          .CIN(n12366), .COUT(n12367), .S0(d_out_d_11__N_1892[9]), .S1(d_out_d_11__N_1892[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_533_13.INIT0 = 16'h9696;
    defparam add_533_13.INIT1 = 16'h9696;
    defparam add_533_13.INJECT1_0 = "NO";
    defparam add_533_13.INJECT1_1 = "NO";
    CCU2D add_533_11 (.A0(d_out_d_11__N_1878[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(d_out_d_11__N_1890[6]), .D0(GND_net), .A1(d_out_d_11__N_1876[17]), 
          .B1(d_out_d_11__N_1890[17]), .C1(d_out_d_11__N_1890[7]), .D1(GND_net), 
          .CIN(n12365), .COUT(n12366), .S0(d_out_d_11__N_1892[7]), .S1(d_out_d_11__N_1892[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_533_11.INIT0 = 16'h9696;
    defparam add_533_11.INIT1 = 16'h9696;
    defparam add_533_11.INJECT1_0 = "NO";
    defparam add_533_11.INJECT1_1 = "NO";
    CCU2D add_533_9 (.A0(d_out_d_11__N_1882[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(d_out_d_11__N_1890[4]), .D0(GND_net), .A1(d_out_d_11__N_1880[17]), 
          .B1(d_out_d_11__N_1890[17]), .C1(d_out_d_11__N_1890[5]), .D1(GND_net), 
          .CIN(n12364), .COUT(n12365), .S0(d_out_d_11__N_1892[5]), .S1(d_out_d_11__N_1892[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_533_9.INIT0 = 16'h9696;
    defparam add_533_9.INIT1 = 16'h9696;
    defparam add_533_9.INJECT1_0 = "NO";
    defparam add_533_9.INJECT1_1 = "NO";
    CCU2D add_533_7 (.A0(d_out_d_11__N_1886[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(d_out_d_11__N_1890[2]), .D0(GND_net), .A1(d_out_d_11__N_1884[17]), 
          .B1(d_out_d_11__N_1890[17]), .C1(d_out_d_11__N_1890[3]), .D1(GND_net), 
          .CIN(n12363), .COUT(n12364), .S0(d_out_d_11__N_1892[3]), .S1(d_out_d_11__N_1892[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_533_7.INIT0 = 16'h9696;
    defparam add_533_7.INIT1 = 16'h9696;
    defparam add_533_7.INJECT1_0 = "NO";
    defparam add_533_7.INJECT1_1 = "NO";
    CCU2D add_533_5 (.A0(d_out_d_11__N_1890[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1888[17]), .B1(d_out_d_11__N_1890[17]), 
          .C1(d_out_d_11__N_1890[1]), .D1(GND_net), .CIN(n12362), .COUT(n12363), 
          .S0(d_out_d_11__N_1892[1]), .S1(d_out_d_11__N_1892[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_533_5.INIT0 = 16'h5aaa;
    defparam add_533_5.INIT1 = 16'h9696;
    defparam add_533_5.INJECT1_0 = "NO";
    defparam add_533_5.INJECT1_1 = "NO";
    CCU2D add_533_3 (.A0(ISquare[2]), .B0(d_out_d_11__N_1890[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12361), .COUT(n12362), .S1(d_out_d_11__N_1892[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_533_3.INIT0 = 16'h5666;
    defparam add_533_3.INIT1 = 16'h5555;
    defparam add_533_3.INJECT1_0 = "NO";
    defparam add_533_3.INJECT1_1 = "NO";
    CCU2D add_533_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1890[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n12361));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_533_1.INIT0 = 16'hF000;
    defparam add_533_1.INIT1 = 16'h0aaa;
    defparam add_533_1.INJECT1_0 = "NO";
    defparam add_533_1.INJECT1_1 = "NO";
    CCU2D add_553_19 (.A0(d_out_d_11__N_1888[14]), .B0(d_out_d_11__N_1888[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1888[15]), .B1(d_out_d_11__N_1888[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12355), .S0(d_out_d_11__N_1890[15]), 
          .S1(d_out_d_11__N_1890[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_553_19.INIT0 = 16'h5999;
    defparam add_553_19.INIT1 = 16'h5999;
    defparam add_553_19.INJECT1_0 = "NO";
    defparam add_553_19.INJECT1_1 = "NO";
    CCU2D add_553_17 (.A0(ISquare[31]), .B0(d_out_d_11__N_1888[17]), .C0(d_out_d_11__N_1888[12]), 
          .D0(GND_net), .A1(d_out_d_11__N_1888[13]), .B1(d_out_d_11__N_1888[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12354), .COUT(n12355), .S0(d_out_d_11__N_1890[13]), 
          .S1(d_out_d_11__N_1890[14]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_553_17.INIT0 = 16'h6969;
    defparam add_553_17.INIT1 = 16'h5999;
    defparam add_553_17.INJECT1_0 = "NO";
    defparam add_553_17.INJECT1_1 = "NO";
    CCU2D add_553_15 (.A0(ISquare[31]), .B0(d_out_d_11__N_1888[17]), .C0(d_out_d_11__N_1888[10]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1888[17]), 
          .C1(d_out_d_11__N_1888[11]), .D1(GND_net), .CIN(n12353), .COUT(n12354), 
          .S0(d_out_d_11__N_1890[11]), .S1(d_out_d_11__N_1890[12]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_553_15.INIT0 = 16'h6969;
    defparam add_553_15.INIT1 = 16'h6969;
    defparam add_553_15.INJECT1_0 = "NO";
    defparam add_553_15.INJECT1_1 = "NO";
    CCU2D add_553_13 (.A0(d_out_d_11__N_1872[17]), .B0(d_out_d_11__N_1888[17]), 
          .C0(d_out_d_11__N_1888[8]), .D0(GND_net), .A1(d_out_d_11__N_1888[9]), 
          .B1(d_out_d_11__N_1888[17]), .C1(GND_net), .D1(GND_net), .CIN(n12352), 
          .COUT(n12353), .S0(d_out_d_11__N_1890[9]), .S1(d_out_d_11__N_1890[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_553_13.INIT0 = 16'h9696;
    defparam add_553_13.INIT1 = 16'h5999;
    defparam add_553_13.INJECT1_0 = "NO";
    defparam add_553_13.INJECT1_1 = "NO";
    LUT4 d_out_d_11__I_1_1_lut (.A(d_out_d_11__N_1874[17]), .Z(d_out_d_11__N_1873)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_1_1_lut.init = 16'h5555;
    CCU2D add_553_11 (.A0(d_out_d_11__N_1876[17]), .B0(d_out_d_11__N_1888[17]), 
          .C0(d_out_d_11__N_1888[6]), .D0(GND_net), .A1(d_out_d_11__N_1874[17]), 
          .B1(d_out_d_11__N_1888[17]), .C1(d_out_d_11__N_1888[7]), .D1(GND_net), 
          .CIN(n12351), .COUT(n12352), .S0(d_out_d_11__N_1890[7]), .S1(d_out_d_11__N_1890[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_553_11.INIT0 = 16'h9696;
    defparam add_553_11.INIT1 = 16'h9696;
    defparam add_553_11.INJECT1_0 = "NO";
    defparam add_553_11.INJECT1_1 = "NO";
    CCU2D add_553_9 (.A0(d_out_d_11__N_1880[17]), .B0(d_out_d_11__N_1888[17]), 
          .C0(d_out_d_11__N_1888[4]), .D0(GND_net), .A1(d_out_d_11__N_1878[17]), 
          .B1(d_out_d_11__N_1888[17]), .C1(d_out_d_11__N_1888[5]), .D1(GND_net), 
          .CIN(n12350), .COUT(n12351), .S0(d_out_d_11__N_1890[5]), .S1(d_out_d_11__N_1890[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_553_9.INIT0 = 16'h9696;
    defparam add_553_9.INIT1 = 16'h9696;
    defparam add_553_9.INJECT1_0 = "NO";
    defparam add_553_9.INJECT1_1 = "NO";
    CCU2D add_553_7 (.A0(d_out_d_11__N_1884[17]), .B0(d_out_d_11__N_1888[17]), 
          .C0(d_out_d_11__N_1888[2]), .D0(GND_net), .A1(d_out_d_11__N_1882[17]), 
          .B1(d_out_d_11__N_1888[17]), .C1(d_out_d_11__N_1888[3]), .D1(GND_net), 
          .CIN(n12349), .COUT(n12350), .S0(d_out_d_11__N_1890[3]), .S1(d_out_d_11__N_1890[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_553_7.INIT0 = 16'h9696;
    defparam add_553_7.INIT1 = 16'h9696;
    defparam add_553_7.INJECT1_0 = "NO";
    defparam add_553_7.INJECT1_1 = "NO";
    CCU2D add_553_5 (.A0(d_out_d_11__N_1888[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1886[17]), .B1(d_out_d_11__N_1888[17]), 
          .C1(d_out_d_11__N_1888[1]), .D1(GND_net), .CIN(n12348), .COUT(n12349), 
          .S0(d_out_d_11__N_1890[1]), .S1(d_out_d_11__N_1890[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_553_5.INIT0 = 16'h5aaa;
    defparam add_553_5.INIT1 = 16'h9696;
    defparam add_553_5.INJECT1_0 = "NO";
    defparam add_553_5.INJECT1_1 = "NO";
    CCU2D add_553_3 (.A0(ISquare[4]), .B0(d_out_d_11__N_1888[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12347), .COUT(n12348), .S1(d_out_d_11__N_1890[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_553_3.INIT0 = 16'h5666;
    defparam add_553_3.INIT1 = 16'h5555;
    defparam add_553_3.INJECT1_0 = "NO";
    defparam add_553_3.INJECT1_1 = "NO";
    CCU2D add_553_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1888[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n12347));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_553_1.INIT0 = 16'hF000;
    defparam add_553_1.INIT1 = 16'h0aaa;
    defparam add_553_1.INJECT1_0 = "NO";
    defparam add_553_1.INJECT1_1 = "NO";
    CCU2D add_433_15 (.A0(d_out_d_11__N_1876[17]), .B0(d_out_d_11__N_1875), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1876[17]), .B1(d_out_d_11__N_1875), 
          .C1(GND_net), .D1(GND_net), .CIN(n12341), .S0(d_out_d_11__N_1878[11]), 
          .S1(d_out_d_11__N_1878[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_433_15.INIT0 = 16'h5666;
    defparam add_433_15.INIT1 = 16'h5666;
    defparam add_433_15.INJECT1_0 = "NO";
    defparam add_433_15.INJECT1_1 = "NO";
    CCU2D add_433_13 (.A0(d_out_d_11__N_1876[8]), .B0(d_out_d_11__N_1876[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1876[9]), .B1(d_out_d_11__N_1876[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12340), .COUT(n12341), .S0(d_out_d_11__N_1878[9]), 
          .S1(d_out_d_11__N_1878[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_433_13.INIT0 = 16'h5999;
    defparam add_433_13.INIT1 = 16'h5999;
    defparam add_433_13.INJECT1_0 = "NO";
    defparam add_433_13.INJECT1_1 = "NO";
    CCU2D add_433_11 (.A0(ISquare[31]), .B0(d_out_d_11__N_1876[17]), .C0(d_out_d_11__N_1876[6]), 
          .D0(GND_net), .A1(d_out_d_11__N_1876[7]), .B1(d_out_d_11__N_1876[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12339), .COUT(n12340), .S0(d_out_d_11__N_1878[7]), 
          .S1(d_out_d_11__N_1878[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_433_11.INIT0 = 16'h6969;
    defparam add_433_11.INIT1 = 16'h5999;
    defparam add_433_11.INJECT1_0 = "NO";
    defparam add_433_11.INJECT1_1 = "NO";
    CCU2D add_433_9 (.A0(ISquare[31]), .B0(d_out_d_11__N_1876[17]), .C0(d_out_d_11__N_1876[4]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1876[17]), 
          .C1(d_out_d_11__N_1876[5]), .D1(GND_net), .CIN(n12338), .COUT(n12339), 
          .S0(d_out_d_11__N_1878[5]), .S1(d_out_d_11__N_1878[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_433_9.INIT0 = 16'h6969;
    defparam add_433_9.INIT1 = 16'h6969;
    defparam add_433_9.INJECT1_0 = "NO";
    defparam add_433_9.INJECT1_1 = "NO";
    CCU2D add_433_7 (.A0(d_out_d_11__N_1872[17]), .B0(d_out_d_11__N_1876[17]), 
          .C0(d_out_d_11__N_1876[2]), .D0(GND_net), .A1(d_out_d_11__N_1876[3]), 
          .B1(d_out_d_11__N_1876[17]), .C1(GND_net), .D1(GND_net), .CIN(n12337), 
          .COUT(n12338), .S0(d_out_d_11__N_1878[3]), .S1(d_out_d_11__N_1878[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_433_7.INIT0 = 16'h9696;
    defparam add_433_7.INIT1 = 16'h5999;
    defparam add_433_7.INJECT1_0 = "NO";
    defparam add_433_7.INJECT1_1 = "NO";
    CCU2D add_433_5 (.A0(d_out_d_11__N_1876[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1874[17]), .B1(d_out_d_11__N_1876[17]), 
          .C1(d_out_d_11__N_1876[1]), .D1(GND_net), .CIN(n12336), .COUT(n12337), 
          .S0(d_out_d_11__N_1878[1]), .S1(d_out_d_11__N_1878[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_433_5.INIT0 = 16'h5aaa;
    defparam add_433_5.INIT1 = 16'h9696;
    defparam add_433_5.INJECT1_0 = "NO";
    defparam add_433_5.INJECT1_1 = "NO";
    CCU2D add_433_3 (.A0(ISquare[16]), .B0(d_out_d_11__N_1876[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12335), .COUT(n12336), .S1(d_out_d_11__N_1878[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_433_3.INIT0 = 16'h5666;
    defparam add_433_3.INIT1 = 16'h5555;
    defparam add_433_3.INJECT1_0 = "NO";
    defparam add_433_3.INJECT1_1 = "NO";
    CCU2D add_433_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1876[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n12335));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_433_1.INIT0 = 16'hF000;
    defparam add_433_1.INIT1 = 16'h0aaa;
    defparam add_433_1.INJECT1_0 = "NO";
    defparam add_433_1.INJECT1_1 = "NO";
    LUT4 d_out_d_11__I_0_1_lut (.A(d_out_d_11__N_1872[17]), .Z(d_out_d_11__N_1871)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_0_1_lut.init = 16'h5555;
    LUT4 i4984_2_lut (.A(ISquare[23]), .B(ISquare[22]), .Z(n12447)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i4984_2_lut.init = 16'h9999;
    LUT4 d_out_d_11__I_9_1_lut (.A(d_out_d_11__N_1890[17]), .Z(d_out_d_11__N_1889)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_9_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_8_1_lut (.A(d_out_d_11__N_1888[17]), .Z(d_out_d_11__N_1887)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_8_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_7_1_lut (.A(d_out_d_11__N_1886[17]), .Z(d_out_d_11__N_1885)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_7_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_6_1_lut (.A(d_out_d_11__N_1884[17]), .Z(d_out_d_11__N_1883)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_6_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_5_1_lut (.A(d_out_d_11__N_1882[17]), .Z(d_out_d_11__N_1881)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_5_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_4_1_lut (.A(d_out_d_11__N_1880[17]), .Z(d_out_d_11__N_1879)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_4_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_3_1_lut (.A(d_out_d_11__N_1878[17]), .Z(d_out_d_11__N_1877)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_3_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_2_1_lut (.A(d_out_d_11__N_1876[17]), .Z(d_out_d_11__N_1875)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_2_1_lut.init = 16'h5555;
    LUT4 i1328_1_lut (.A(ISquare[31]), .Z(n209)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1328_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_10_1_lut (.A(d_out_d_11__N_1892[17]), .Z(d_out_d_11__N_1891)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_10_1_lut.init = 16'h5555;
    Multiplier Multiplier2 (.CIC1_out_clkSin(CIC1_out_clkSin), .VCC_net(VCC_net), 
            .GND_net(GND_net), .MultDataC({MultDataC}), .MultResult2({MultResult2})) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    Multiplier_U0 Multiplier1 (.CIC1_out_clkSin(CIC1_out_clkSin), .VCC_net(VCC_net), 
            .GND_net(GND_net), .MultDataB({MultDataB}), .MultResult1({MultResult1})) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    
endmodule
//
// Verilog Description of module Multiplier
//

module Multiplier (CIC1_out_clkSin, VCC_net, GND_net, MultDataC, MultResult2) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input CIC1_out_clkSin;
    input VCC_net;
    input GND_net;
    input [11:0]MultDataC;
    output [23:0]MultResult2;
    
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(82[6:21])
    
    wire Multiplier_0_mult_0_5_n1, regb_b_1, rega_a_11, Multiplier_0_pp_1_2, 
        regb_b_2, regb_b_0, Multiplier_0_mult_2_5_n1, regb_b_3, Multiplier_0_pp_2_4, 
        regb_b_4, Multiplier_0_mult_4_5_n1, regb_b_5, Multiplier_0_pp_3_6, 
        regb_b_6, Multiplier_0_mult_6_5_n1, regb_b_7, Multiplier_0_pp_4_8, 
        regb_b_8, Multiplier_0_mult_8_5_n1, regb_b_9, Multiplier_0_pp_5_10, 
        regb_b_10, Multiplier_0_mult_10_0_n0, regb_b_11, Multiplier_0_mult_10_1_n1, 
        rega_a_3, rega_a_2, Multiplier_0_mult_10_1_n0, Multiplier_0_mult_10_2_n1, 
        rega_a_5, rega_a_4, Multiplier_0_mult_10_2_n0, Multiplier_0_mult_10_3_n1, 
        rega_a_7, rega_a_6, Multiplier_0_mult_10_3_n0, Multiplier_0_mult_10_4_n1, 
        rega_a_9, rega_a_8, Multiplier_0_mult_10_4_n0, Multiplier_0_mult_10_5_n2, 
        rega_a_10, Multiplier_0_mult_10_5_n0, rega_a_1, rego_o_0, rego_o_1, 
        rego_o_2, rego_o_3, rego_o_4, rego_o_5, rego_o_6, rego_o_7, 
        rego_o_8, rego_o_9, rego_o_10, rego_o_11, rego_o_12, rego_o_13, 
        rego_o_14, rego_o_15, rego_o_16, rego_o_17, rego_o_18, rego_o_19, 
        rego_o_20, rego_o_21, rego_o_22, rego_o_23, Multiplier_0_pp_0_0, 
        Multiplier_0_pp_0_1, s_Multiplier_0_0_2, s_Multiplier_0_0_3, s_Multiplier_0_0_4, 
        f_s_Multiplier_0_0_4, s_Multiplier_0_0_5, f_s_Multiplier_0_0_5, 
        s_Multiplier_0_0_6, f_s_Multiplier_0_0_6, s_Multiplier_0_0_7, 
        f_s_Multiplier_0_0_7, s_Multiplier_0_0_8, f_s_Multiplier_0_0_8, 
        s_Multiplier_0_0_9, f_s_Multiplier_0_0_9, s_Multiplier_0_0_10, 
        f_s_Multiplier_0_0_10, s_Multiplier_0_0_11, f_s_Multiplier_0_0_11, 
        s_Multiplier_0_0_12, f_s_Multiplier_0_0_12, s_Multiplier_0_0_13, 
        f_s_Multiplier_0_0_13, s_Multiplier_0_0_14, f_s_Multiplier_0_0_14, 
        s_Multiplier_0_0_15, f_s_Multiplier_0_0_15, s_Multiplier_0_0_16, 
        f_s_Multiplier_0_0_16, s_Multiplier_0_0_17, f_s_Multiplier_0_0_17, 
        f_Multiplier_0_pp_2_4, f_Multiplier_0_pp_2_5, Multiplier_0_pp_2_5, 
        s_Multiplier_0_1_6, f_s_Multiplier_0_1_6, s_Multiplier_0_1_7, 
        f_s_Multiplier_0_1_7, s_Multiplier_0_1_8, f_s_Multiplier_0_1_8, 
        s_Multiplier_0_1_9, f_s_Multiplier_0_1_9, s_Multiplier_0_1_10, 
        f_s_Multiplier_0_1_10, s_Multiplier_0_1_11, f_s_Multiplier_0_1_11, 
        s_Multiplier_0_1_12, f_s_Multiplier_0_1_12, s_Multiplier_0_1_13, 
        f_s_Multiplier_0_1_13, s_Multiplier_0_1_14, f_s_Multiplier_0_1_14, 
        s_Multiplier_0_1_15, f_s_Multiplier_0_1_15, s_Multiplier_0_1_16, 
        f_s_Multiplier_0_1_16, s_Multiplier_0_1_17, f_s_Multiplier_0_1_17, 
        s_Multiplier_0_1_18, f_s_Multiplier_0_1_18, s_Multiplier_0_1_19, 
        f_s_Multiplier_0_1_19, s_Multiplier_0_1_20, f_s_Multiplier_0_1_20, 
        s_Multiplier_0_1_21, f_s_Multiplier_0_1_21, f_Multiplier_0_pp_4_8, 
        f_Multiplier_0_pp_4_9, Multiplier_0_pp_4_9, s_Multiplier_0_2_10, 
        f_s_Multiplier_0_2_10, s_Multiplier_0_2_11, f_s_Multiplier_0_2_11, 
        s_Multiplier_0_2_12, f_s_Multiplier_0_2_12, s_Multiplier_0_2_13, 
        f_s_Multiplier_0_2_13, s_Multiplier_0_2_14, f_s_Multiplier_0_2_14, 
        s_Multiplier_0_2_15, f_s_Multiplier_0_2_15, s_Multiplier_0_2_16, 
        f_s_Multiplier_0_2_16, s_Multiplier_0_2_17, f_s_Multiplier_0_2_17, 
        s_Multiplier_0_2_18, f_s_Multiplier_0_2_18, s_Multiplier_0_2_19, 
        f_s_Multiplier_0_2_19, s_Multiplier_0_2_20, f_s_Multiplier_0_2_20, 
        s_Multiplier_0_2_21, f_s_Multiplier_0_2_21, s_Multiplier_0_2_22, 
        f_s_Multiplier_0_2_22, s_Multiplier_0_2_23, f_s_Multiplier_0_2_23, 
        Multiplier_0_cin_lr_0, Multiplier_0_pp_0_13, mfco, Multiplier_0_cin_lr_2, 
        Multiplier_0_pp_1_15, mfco_1, Multiplier_0_cin_lr_4, Multiplier_0_pp_2_17, 
        mfco_2, Multiplier_0_cin_lr_6, Multiplier_0_pp_3_19, mfco_3, 
        Multiplier_0_cin_lr_8, Multiplier_0_pp_4_21, mfco_4, Multiplier_0_cin_lr_10, 
        Multiplier_0_pp_5_23, mfco_5, co_Multiplier_0_0_1, Multiplier_0_pp_0_2, 
        co_Multiplier_0_0_2, Multiplier_0_pp_0_4, Multiplier_0_pp_0_3, 
        Multiplier_0_pp_1_4, Multiplier_0_pp_1_3, co_Multiplier_0_0_3, 
        Multiplier_0_pp_0_6, Multiplier_0_pp_0_5, Multiplier_0_pp_1_6, 
        Multiplier_0_pp_1_5, co_Multiplier_0_0_4, Multiplier_0_pp_0_8, 
        Multiplier_0_pp_0_7, Multiplier_0_pp_1_8, Multiplier_0_pp_1_7, 
        co_Multiplier_0_0_5, Multiplier_0_pp_0_10, Multiplier_0_pp_0_9, 
        Multiplier_0_pp_1_10, Multiplier_0_pp_1_9, co_Multiplier_0_0_6, 
        Multiplier_0_pp_0_12, Multiplier_0_pp_0_11, Multiplier_0_pp_1_12, 
        Multiplier_0_pp_1_11, co_Multiplier_0_0_7, Multiplier_0_pp_1_14, 
        Multiplier_0_pp_1_13, co_Multiplier_0_0_8, co_Multiplier_0_1_1, 
        Multiplier_0_pp_2_6, co_Multiplier_0_1_2, Multiplier_0_pp_2_8, 
        Multiplier_0_pp_2_7, Multiplier_0_pp_3_8, Multiplier_0_pp_3_7, 
        co_Multiplier_0_1_3, Multiplier_0_pp_2_10, Multiplier_0_pp_2_9, 
        Multiplier_0_pp_3_10, Multiplier_0_pp_3_9, co_Multiplier_0_1_4, 
        Multiplier_0_pp_2_12, Multiplier_0_pp_2_11, Multiplier_0_pp_3_12, 
        Multiplier_0_pp_3_11, co_Multiplier_0_1_5, Multiplier_0_pp_2_14, 
        Multiplier_0_pp_2_13, Multiplier_0_pp_3_14, Multiplier_0_pp_3_13, 
        co_Multiplier_0_1_6, Multiplier_0_pp_2_16, Multiplier_0_pp_2_15, 
        Multiplier_0_pp_3_16, Multiplier_0_pp_3_15, co_Multiplier_0_1_7, 
        Multiplier_0_pp_3_18, Multiplier_0_pp_3_17, co_Multiplier_0_1_8, 
        co_Multiplier_0_2_1, Multiplier_0_pp_4_10, co_Multiplier_0_2_2, 
        Multiplier_0_pp_4_12, Multiplier_0_pp_4_11, Multiplier_0_pp_5_12, 
        Multiplier_0_pp_5_11, co_Multiplier_0_2_3, Multiplier_0_pp_4_14, 
        Multiplier_0_pp_4_13, Multiplier_0_pp_5_14, Multiplier_0_pp_5_13, 
        co_Multiplier_0_2_4, Multiplier_0_pp_4_16, Multiplier_0_pp_4_15, 
        Multiplier_0_pp_5_16, Multiplier_0_pp_5_15, co_Multiplier_0_2_5, 
        Multiplier_0_pp_4_18, Multiplier_0_pp_4_17, Multiplier_0_pp_5_18, 
        Multiplier_0_pp_5_17, co_Multiplier_0_2_6, Multiplier_0_pp_4_20, 
        Multiplier_0_pp_4_19, Multiplier_0_pp_5_20, Multiplier_0_pp_5_19, 
        co_Multiplier_0_2_7, Multiplier_0_pp_5_22, Multiplier_0_pp_5_21, 
        co_Multiplier_0_3_1, co_Multiplier_0_3_2, co_Multiplier_0_3_3, 
        s_Multiplier_0_3_8, co_Multiplier_0_3_4, s_Multiplier_0_3_9, s_Multiplier_0_3_10, 
        co_Multiplier_0_3_5, s_Multiplier_0_3_11, s_Multiplier_0_3_12, 
        co_Multiplier_0_3_6, s_Multiplier_0_3_13, s_Multiplier_0_3_14, 
        co_Multiplier_0_3_7, s_Multiplier_0_3_15, s_Multiplier_0_3_16, 
        co_Multiplier_0_3_8, s_Multiplier_0_3_17, s_Multiplier_0_3_18, 
        co_Multiplier_0_3_9, s_Multiplier_0_3_19, s_Multiplier_0_3_20, 
        co_Multiplier_0_3_10, s_Multiplier_0_3_21, s_Multiplier_0_3_22, 
        s_Multiplier_0_3_23, co_t_Multiplier_0_4_1, co_t_Multiplier_0_4_2, 
        co_t_Multiplier_0_4_3, co_t_Multiplier_0_4_4, co_t_Multiplier_0_4_5, 
        co_t_Multiplier_0_4_6, co_t_Multiplier_0_4_7, co_t_Multiplier_0_4_8, 
        mco, mco_1, mco_2, mco_3, mco_4, Multiplier_0_mult_0_5_n2, 
        mco_5, mco_6, mco_7, mco_8, mco_9, Multiplier_0_mult_2_5_n2, 
        mco_10, mco_11, mco_12, mco_13, mco_14, Multiplier_0_mult_4_5_n2, 
        mco_15, mco_16, mco_17, mco_18, mco_19, Multiplier_0_mult_6_5_n2, 
        mco_20, mco_21, mco_22, mco_23, mco_24, Multiplier_0_mult_8_5_n2, 
        Multiplier_0_mult_10_0_n1, mco_25, mco_26, mco_27, mco_28, 
        mco_29;
    
    ND2 ND2_t25 (.A(rega_a_11), .B(regb_b_1), .Z(Multiplier_0_mult_0_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    AND2 AND2_t24 (.A(regb_b_0), .B(regb_b_2), .Z(Multiplier_0_pp_1_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(382[10:72])
    ND2 ND2_t22 (.A(rega_a_11), .B(regb_b_3), .Z(Multiplier_0_mult_2_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    AND2 AND2_t21 (.A(regb_b_0), .B(regb_b_4), .Z(Multiplier_0_pp_2_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(388[10:72])
    ND2 ND2_t19 (.A(rega_a_11), .B(regb_b_5), .Z(Multiplier_0_mult_4_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    AND2 AND2_t18 (.A(regb_b_0), .B(regb_b_6), .Z(Multiplier_0_pp_3_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(394[10:72])
    ND2 ND2_t16 (.A(rega_a_11), .B(regb_b_7), .Z(Multiplier_0_mult_6_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    AND2 AND2_t15 (.A(regb_b_0), .B(regb_b_8), .Z(Multiplier_0_pp_4_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(400[10:72])
    ND2 ND2_t13 (.A(rega_a_11), .B(regb_b_9), .Z(Multiplier_0_mult_8_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    AND2 AND2_t12 (.A(regb_b_0), .B(regb_b_10), .Z(Multiplier_0_pp_5_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(406[10:74])
    ND2 ND2_t10 (.A(regb_b_0), .B(regb_b_11), .Z(Multiplier_0_mult_10_0_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t9 (.A(rega_a_3), .B(regb_b_11), .Z(Multiplier_0_mult_10_1_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t8 (.A(rega_a_2), .B(regb_b_11), .Z(Multiplier_0_mult_10_1_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t7 (.A(rega_a_5), .B(regb_b_11), .Z(Multiplier_0_mult_10_2_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t6 (.A(rega_a_4), .B(regb_b_11), .Z(Multiplier_0_mult_10_2_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t5 (.A(rega_a_7), .B(regb_b_11), .Z(Multiplier_0_mult_10_3_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t4 (.A(rega_a_6), .B(regb_b_11), .Z(Multiplier_0_mult_10_3_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t3 (.A(rega_a_9), .B(regb_b_11), .Z(Multiplier_0_mult_10_4_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t2 (.A(rega_a_8), .B(regb_b_11), .Z(Multiplier_0_mult_10_4_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t1 (.A(rega_a_11), .B(regb_b_10), .Z(Multiplier_0_mult_10_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t0 (.A(rega_a_10), .B(regb_b_11), .Z(Multiplier_0_mult_10_5_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FD1P3DX FF_98 (.D(MultDataC[1]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(435[13:82])
    defparam FF_98.GSR = "ENABLED";
    FD1P3DX FF_97 (.D(MultDataC[2]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(438[13:82])
    defparam FF_97.GSR = "ENABLED";
    FD1P3DX FF_96 (.D(MultDataC[3]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(441[13:82])
    defparam FF_96.GSR = "ENABLED";
    FD1P3DX FF_95 (.D(MultDataC[4]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(444[13:82])
    defparam FF_95.GSR = "ENABLED";
    FD1P3DX FF_94 (.D(MultDataC[5]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(447[13:82])
    defparam FF_94.GSR = "ENABLED";
    FD1P3DX FF_93 (.D(MultDataC[6]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(450[13:82])
    defparam FF_93.GSR = "ENABLED";
    FD1P3DX FF_92 (.D(MultDataC[7]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(453[13:82])
    defparam FF_92.GSR = "ENABLED";
    FD1P3DX FF_91 (.D(MultDataC[8]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(456[13:82])
    defparam FF_91.GSR = "ENABLED";
    FD1P3DX FF_90 (.D(MultDataC[9]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(459[13:82])
    defparam FF_90.GSR = "ENABLED";
    FD1P3DX FF_89 (.D(MultDataC[10]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(462[13:84])
    defparam FF_89.GSR = "ENABLED";
    FD1P3DX FF_88 (.D(MultDataC[11]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(465[13:84])
    defparam FF_88.GSR = "ENABLED";
    FD1P3DX FF_87 (.D(MultDataC[0]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_0)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(468[13:82])
    defparam FF_87.GSR = "ENABLED";
    FD1P3DX FF_86 (.D(MultDataC[1]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(471[13:82])
    defparam FF_86.GSR = "ENABLED";
    FD1P3DX FF_85 (.D(MultDataC[2]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(474[13:82])
    defparam FF_85.GSR = "ENABLED";
    FD1P3DX FF_84 (.D(MultDataC[3]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(477[13:82])
    defparam FF_84.GSR = "ENABLED";
    FD1P3DX FF_83 (.D(MultDataC[4]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(480[13:82])
    defparam FF_83.GSR = "ENABLED";
    FD1P3DX FF_82 (.D(MultDataC[5]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(483[13:82])
    defparam FF_82.GSR = "ENABLED";
    FD1P3DX FF_81 (.D(MultDataC[6]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(486[13:82])
    defparam FF_81.GSR = "ENABLED";
    FD1P3DX FF_80 (.D(MultDataC[7]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(489[13:82])
    defparam FF_80.GSR = "ENABLED";
    FD1P3DX FF_79 (.D(MultDataC[8]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(492[13:82])
    defparam FF_79.GSR = "ENABLED";
    FD1P3DX FF_78 (.D(MultDataC[9]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(495[13:82])
    defparam FF_78.GSR = "ENABLED";
    FD1P3DX FF_77 (.D(MultDataC[10]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(498[13:84])
    defparam FF_77.GSR = "ENABLED";
    FD1P3DX FF_76 (.D(MultDataC[11]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(501[13:84])
    defparam FF_76.GSR = "ENABLED";
    FD1P3DX FF_75 (.D(rego_o_0), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[0])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(504[13:83])
    defparam FF_75.GSR = "ENABLED";
    FD1P3DX FF_74 (.D(rego_o_1), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[1])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(507[13:83])
    defparam FF_74.GSR = "ENABLED";
    FD1P3DX FF_73 (.D(rego_o_2), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[2])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(510[13:83])
    defparam FF_73.GSR = "ENABLED";
    FD1P3DX FF_72 (.D(rego_o_3), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[3])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(513[13:83])
    defparam FF_72.GSR = "ENABLED";
    FD1P3DX FF_71 (.D(rego_o_4), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[4])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(516[13:83])
    defparam FF_71.GSR = "ENABLED";
    FD1P3DX FF_70 (.D(rego_o_5), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[5])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(519[13:83])
    defparam FF_70.GSR = "ENABLED";
    FD1P3DX FF_69 (.D(rego_o_6), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[6])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(522[13:83])
    defparam FF_69.GSR = "ENABLED";
    FD1P3DX FF_68 (.D(rego_o_7), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[7])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(525[13:83])
    defparam FF_68.GSR = "ENABLED";
    FD1P3DX FF_67 (.D(rego_o_8), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[8])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(528[13:83])
    defparam FF_67.GSR = "ENABLED";
    FD1P3DX FF_66 (.D(rego_o_9), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[9])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(531[13:83])
    defparam FF_66.GSR = "ENABLED";
    FD1P3DX FF_65 (.D(rego_o_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[10])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(534[13:85])
    defparam FF_65.GSR = "ENABLED";
    FD1P3DX FF_64 (.D(rego_o_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[11])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(537[13:85])
    defparam FF_64.GSR = "ENABLED";
    FD1P3DX FF_63 (.D(rego_o_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[12])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(540[13:85])
    defparam FF_63.GSR = "ENABLED";
    FD1P3DX FF_62 (.D(rego_o_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[13])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(543[13:85])
    defparam FF_62.GSR = "ENABLED";
    FD1P3DX FF_61 (.D(rego_o_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[14])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(546[13:85])
    defparam FF_61.GSR = "ENABLED";
    FD1P3DX FF_60 (.D(rego_o_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[15])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(549[13:85])
    defparam FF_60.GSR = "ENABLED";
    FD1P3DX FF_59 (.D(rego_o_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[16])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(552[13:85])
    defparam FF_59.GSR = "ENABLED";
    FD1P3DX FF_58 (.D(rego_o_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[17])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(555[13:85])
    defparam FF_58.GSR = "ENABLED";
    FD1P3DX FF_57 (.D(rego_o_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[18])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(558[13:85])
    defparam FF_57.GSR = "ENABLED";
    FD1P3DX FF_56 (.D(rego_o_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[19])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(561[13:85])
    defparam FF_56.GSR = "ENABLED";
    FD1P3DX FF_55 (.D(rego_o_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[20])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(564[13:85])
    defparam FF_55.GSR = "ENABLED";
    FD1P3DX FF_54 (.D(rego_o_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[21])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(567[13:85])
    defparam FF_54.GSR = "ENABLED";
    FD1P3DX FF_53 (.D(rego_o_22), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[22])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(570[13:85])
    defparam FF_53.GSR = "ENABLED";
    FD1P3DX FF_52 (.D(rego_o_23), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[23])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(573[13:85])
    defparam FF_52.GSR = "ENABLED";
    FD1P3DX FF_51 (.D(Multiplier_0_pp_0_0), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_0)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(576[13] 577[35])
    defparam FF_51.GSR = "ENABLED";
    FD1P3DX FF_50 (.D(Multiplier_0_pp_0_1), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(580[13] 581[35])
    defparam FF_50.GSR = "ENABLED";
    FD1P3DX FF_49 (.D(s_Multiplier_0_0_2), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(584[13] 585[34])
    defparam FF_49.GSR = "ENABLED";
    FD1P3DX FF_48 (.D(s_Multiplier_0_0_3), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(588[13] 589[34])
    defparam FF_48.GSR = "ENABLED";
    FD1P3DX FF_47 (.D(s_Multiplier_0_0_4), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(592[13] 593[34])
    defparam FF_47.GSR = "ENABLED";
    FD1P3DX FF_46 (.D(s_Multiplier_0_0_5), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(596[13] 597[34])
    defparam FF_46.GSR = "ENABLED";
    FD1P3DX FF_45 (.D(s_Multiplier_0_0_6), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(600[13] 601[34])
    defparam FF_45.GSR = "ENABLED";
    FD1P3DX FF_44 (.D(s_Multiplier_0_0_7), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(604[13] 605[34])
    defparam FF_44.GSR = "ENABLED";
    FD1P3DX FF_43 (.D(s_Multiplier_0_0_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(608[13] 609[34])
    defparam FF_43.GSR = "ENABLED";
    FD1P3DX FF_42 (.D(s_Multiplier_0_0_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(612[13] 613[34])
    defparam FF_42.GSR = "ENABLED";
    FD1P3DX FF_41 (.D(s_Multiplier_0_0_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(616[13] 617[35])
    defparam FF_41.GSR = "ENABLED";
    FD1P3DX FF_40 (.D(s_Multiplier_0_0_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(620[13] 621[35])
    defparam FF_40.GSR = "ENABLED";
    FD1P3DX FF_39 (.D(s_Multiplier_0_0_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(624[13] 625[35])
    defparam FF_39.GSR = "ENABLED";
    FD1P3DX FF_38 (.D(s_Multiplier_0_0_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(628[13] 629[35])
    defparam FF_38.GSR = "ENABLED";
    FD1P3DX FF_37 (.D(s_Multiplier_0_0_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(632[13] 633[35])
    defparam FF_37.GSR = "ENABLED";
    FD1P3DX FF_36 (.D(s_Multiplier_0_0_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(636[13] 637[35])
    defparam FF_36.GSR = "ENABLED";
    FD1P3DX FF_35 (.D(s_Multiplier_0_0_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(640[13] 641[35])
    defparam FF_35.GSR = "ENABLED";
    FD1P3DX FF_34 (.D(s_Multiplier_0_0_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(644[13] 645[35])
    defparam FF_34.GSR = "ENABLED";
    FD1P3DX FF_33 (.D(Multiplier_0_pp_2_4), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_2_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(648[13] 649[35])
    defparam FF_33.GSR = "ENABLED";
    FD1P3DX FF_32 (.D(Multiplier_0_pp_2_5), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_2_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(652[13] 653[35])
    defparam FF_32.GSR = "ENABLED";
    FD1P3DX FF_31 (.D(s_Multiplier_0_1_6), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(656[13] 657[34])
    defparam FF_31.GSR = "ENABLED";
    FD1P3DX FF_30 (.D(s_Multiplier_0_1_7), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(660[13] 661[34])
    defparam FF_30.GSR = "ENABLED";
    FD1P3DX FF_29 (.D(s_Multiplier_0_1_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(664[13] 665[34])
    defparam FF_29.GSR = "ENABLED";
    FD1P3DX FF_28 (.D(s_Multiplier_0_1_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(668[13] 669[34])
    defparam FF_28.GSR = "ENABLED";
    FD1P3DX FF_27 (.D(s_Multiplier_0_1_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(672[13] 673[35])
    defparam FF_27.GSR = "ENABLED";
    FD1P3DX FF_26 (.D(s_Multiplier_0_1_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(676[13] 677[35])
    defparam FF_26.GSR = "ENABLED";
    FD1P3DX FF_25 (.D(s_Multiplier_0_1_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(680[13] 681[35])
    defparam FF_25.GSR = "ENABLED";
    FD1P3DX FF_24 (.D(s_Multiplier_0_1_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(684[13] 685[35])
    defparam FF_24.GSR = "ENABLED";
    FD1P3DX FF_23 (.D(s_Multiplier_0_1_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(688[13] 689[35])
    defparam FF_23.GSR = "ENABLED";
    FD1P3DX FF_22 (.D(s_Multiplier_0_1_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(692[13] 693[35])
    defparam FF_22.GSR = "ENABLED";
    FD1P3DX FF_21 (.D(s_Multiplier_0_1_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(696[13] 697[35])
    defparam FF_21.GSR = "ENABLED";
    FD1P3DX FF_20 (.D(s_Multiplier_0_1_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(700[13] 701[35])
    defparam FF_20.GSR = "ENABLED";
    FD1P3DX FF_19 (.D(s_Multiplier_0_1_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(704[13] 705[35])
    defparam FF_19.GSR = "ENABLED";
    FD1P3DX FF_18 (.D(s_Multiplier_0_1_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(708[13] 709[35])
    defparam FF_18.GSR = "ENABLED";
    FD1P3DX FF_17 (.D(s_Multiplier_0_1_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(712[13] 713[35])
    defparam FF_17.GSR = "ENABLED";
    FD1P3DX FF_16 (.D(s_Multiplier_0_1_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(716[13] 717[35])
    defparam FF_16.GSR = "ENABLED";
    FD1P3DX FF_15 (.D(Multiplier_0_pp_4_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_4_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(720[13] 721[35])
    defparam FF_15.GSR = "ENABLED";
    FD1P3DX FF_14 (.D(Multiplier_0_pp_4_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_4_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(724[13] 725[35])
    defparam FF_14.GSR = "ENABLED";
    FD1P3DX FF_13 (.D(s_Multiplier_0_2_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(728[13] 729[35])
    defparam FF_13.GSR = "ENABLED";
    FD1P3DX FF_12 (.D(s_Multiplier_0_2_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(732[13] 733[35])
    defparam FF_12.GSR = "ENABLED";
    FD1P3DX FF_11 (.D(s_Multiplier_0_2_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(736[13] 737[35])
    defparam FF_11.GSR = "ENABLED";
    FD1P3DX FF_10 (.D(s_Multiplier_0_2_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(740[13] 741[35])
    defparam FF_10.GSR = "ENABLED";
    FD1P3DX FF_9 (.D(s_Multiplier_0_2_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(744[13] 745[35])
    defparam FF_9.GSR = "ENABLED";
    FD1P3DX FF_8 (.D(s_Multiplier_0_2_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(748[13] 749[35])
    defparam FF_8.GSR = "ENABLED";
    FD1P3DX FF_7 (.D(s_Multiplier_0_2_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(752[13] 753[35])
    defparam FF_7.GSR = "ENABLED";
    FD1P3DX FF_6 (.D(s_Multiplier_0_2_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(756[13] 757[35])
    defparam FF_6.GSR = "ENABLED";
    FD1P3DX FF_5 (.D(s_Multiplier_0_2_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(760[13] 761[35])
    defparam FF_5.GSR = "ENABLED";
    FD1P3DX FF_4 (.D(s_Multiplier_0_2_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(764[13] 765[35])
    defparam FF_4.GSR = "ENABLED";
    FD1P3DX FF_3 (.D(s_Multiplier_0_2_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(768[13] 769[35])
    defparam FF_3.GSR = "ENABLED";
    FD1P3DX FF_2 (.D(s_Multiplier_0_2_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(772[13] 773[35])
    defparam FF_2.GSR = "ENABLED";
    FD1P3DX FF_1 (.D(s_Multiplier_0_2_22), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_22)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(776[13] 777[35])
    defparam FF_1.GSR = "ENABLED";
    FD1P3DX FF_0 (.D(s_Multiplier_0_2_23), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_23)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(780[13] 781[35])
    defparam FF_0.GSR = "ENABLED";
    FADD2B Multiplier_0_cin_lr_add_0 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_Cadd_0_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco), .S0(Multiplier_0_pp_0_13)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_cin_lr_add_2 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_Cadd_2_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_1), .S0(Multiplier_0_pp_1_15)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_cin_lr_add_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_Cadd_4_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_2), .S0(Multiplier_0_pp_2_17)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_cin_lr_add_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_Cadd_6_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_3), .S0(Multiplier_0_pp_3_19)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_cin_lr_add_8 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_Cadd_8_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_4), .S0(Multiplier_0_pp_4_21)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_cin_lr_add_10 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_Cadd_10_6 (.A0(VCC_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_5), .S0(Multiplier_0_pp_5_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_Multiplier_0_0_1 (.A0(GND_net), .A1(Multiplier_0_pp_0_2), 
           .B0(GND_net), .B1(Multiplier_0_pp_1_2), .CI(GND_net), .COUT(co_Multiplier_0_0_1), 
           .S1(s_Multiplier_0_0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_0_2 (.A0(Multiplier_0_pp_0_3), .A1(Multiplier_0_pp_0_4), 
           .B0(Multiplier_0_pp_1_3), .B1(Multiplier_0_pp_1_4), .CI(co_Multiplier_0_0_1), 
           .COUT(co_Multiplier_0_0_2), .S0(s_Multiplier_0_0_3), .S1(s_Multiplier_0_0_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_0_3 (.A0(Multiplier_0_pp_0_5), .A1(Multiplier_0_pp_0_6), 
           .B0(Multiplier_0_pp_1_5), .B1(Multiplier_0_pp_1_6), .CI(co_Multiplier_0_0_2), 
           .COUT(co_Multiplier_0_0_3), .S0(s_Multiplier_0_0_5), .S1(s_Multiplier_0_0_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_0_4 (.A0(Multiplier_0_pp_0_7), .A1(Multiplier_0_pp_0_8), 
           .B0(Multiplier_0_pp_1_7), .B1(Multiplier_0_pp_1_8), .CI(co_Multiplier_0_0_3), 
           .COUT(co_Multiplier_0_0_4), .S0(s_Multiplier_0_0_7), .S1(s_Multiplier_0_0_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_0_5 (.A0(Multiplier_0_pp_0_9), .A1(Multiplier_0_pp_0_10), 
           .B0(Multiplier_0_pp_1_9), .B1(Multiplier_0_pp_1_10), .CI(co_Multiplier_0_0_4), 
           .COUT(co_Multiplier_0_0_5), .S0(s_Multiplier_0_0_9), .S1(s_Multiplier_0_0_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_0_6 (.A0(Multiplier_0_pp_0_11), .A1(Multiplier_0_pp_0_12), 
           .B0(Multiplier_0_pp_1_11), .B1(Multiplier_0_pp_1_12), .CI(co_Multiplier_0_0_5), 
           .COUT(co_Multiplier_0_0_6), .S0(s_Multiplier_0_0_11), .S1(s_Multiplier_0_0_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_0_7 (.A0(Multiplier_0_pp_0_13), .A1(GND_net), 
           .B0(Multiplier_0_pp_1_13), .B1(Multiplier_0_pp_1_14), .CI(co_Multiplier_0_0_6), 
           .COUT(co_Multiplier_0_0_7), .S0(s_Multiplier_0_0_13), .S1(s_Multiplier_0_0_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_0_8 (.A0(GND_net), .A1(GND_net), .B0(Multiplier_0_pp_1_15), 
           .B1(GND_net), .CI(co_Multiplier_0_0_7), .COUT(co_Multiplier_0_0_8), 
           .S0(s_Multiplier_0_0_15), .S1(s_Multiplier_0_0_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_Multiplier_0_0_9 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_Multiplier_0_0_8), .S0(s_Multiplier_0_0_17)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_Multiplier_0_1_1 (.A0(GND_net), .A1(Multiplier_0_pp_2_6), 
           .B0(GND_net), .B1(Multiplier_0_pp_3_6), .CI(GND_net), .COUT(co_Multiplier_0_1_1), 
           .S1(s_Multiplier_0_1_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_1_2 (.A0(Multiplier_0_pp_2_7), .A1(Multiplier_0_pp_2_8), 
           .B0(Multiplier_0_pp_3_7), .B1(Multiplier_0_pp_3_8), .CI(co_Multiplier_0_1_1), 
           .COUT(co_Multiplier_0_1_2), .S0(s_Multiplier_0_1_7), .S1(s_Multiplier_0_1_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_1_3 (.A0(Multiplier_0_pp_2_9), .A1(Multiplier_0_pp_2_10), 
           .B0(Multiplier_0_pp_3_9), .B1(Multiplier_0_pp_3_10), .CI(co_Multiplier_0_1_2), 
           .COUT(co_Multiplier_0_1_3), .S0(s_Multiplier_0_1_9), .S1(s_Multiplier_0_1_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_1_4 (.A0(Multiplier_0_pp_2_11), .A1(Multiplier_0_pp_2_12), 
           .B0(Multiplier_0_pp_3_11), .B1(Multiplier_0_pp_3_12), .CI(co_Multiplier_0_1_3), 
           .COUT(co_Multiplier_0_1_4), .S0(s_Multiplier_0_1_11), .S1(s_Multiplier_0_1_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_1_5 (.A0(Multiplier_0_pp_2_13), .A1(Multiplier_0_pp_2_14), 
           .B0(Multiplier_0_pp_3_13), .B1(Multiplier_0_pp_3_14), .CI(co_Multiplier_0_1_4), 
           .COUT(co_Multiplier_0_1_5), .S0(s_Multiplier_0_1_13), .S1(s_Multiplier_0_1_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_1_6 (.A0(Multiplier_0_pp_2_15), .A1(Multiplier_0_pp_2_16), 
           .B0(Multiplier_0_pp_3_15), .B1(Multiplier_0_pp_3_16), .CI(co_Multiplier_0_1_5), 
           .COUT(co_Multiplier_0_1_6), .S0(s_Multiplier_0_1_15), .S1(s_Multiplier_0_1_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_1_7 (.A0(Multiplier_0_pp_2_17), .A1(GND_net), 
           .B0(Multiplier_0_pp_3_17), .B1(Multiplier_0_pp_3_18), .CI(co_Multiplier_0_1_6), 
           .COUT(co_Multiplier_0_1_7), .S0(s_Multiplier_0_1_17), .S1(s_Multiplier_0_1_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_1_8 (.A0(GND_net), .A1(GND_net), .B0(Multiplier_0_pp_3_19), 
           .B1(GND_net), .CI(co_Multiplier_0_1_7), .COUT(co_Multiplier_0_1_8), 
           .S0(s_Multiplier_0_1_19), .S1(s_Multiplier_0_1_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_Multiplier_0_1_9 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_Multiplier_0_1_8), .S0(s_Multiplier_0_1_21)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_Multiplier_0_2_1 (.A0(GND_net), .A1(Multiplier_0_pp_4_10), 
           .B0(GND_net), .B1(Multiplier_0_pp_5_10), .CI(GND_net), .COUT(co_Multiplier_0_2_1), 
           .S1(s_Multiplier_0_2_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_2_2 (.A0(Multiplier_0_pp_4_11), .A1(Multiplier_0_pp_4_12), 
           .B0(Multiplier_0_pp_5_11), .B1(Multiplier_0_pp_5_12), .CI(co_Multiplier_0_2_1), 
           .COUT(co_Multiplier_0_2_2), .S0(s_Multiplier_0_2_11), .S1(s_Multiplier_0_2_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_2_3 (.A0(Multiplier_0_pp_4_13), .A1(Multiplier_0_pp_4_14), 
           .B0(Multiplier_0_pp_5_13), .B1(Multiplier_0_pp_5_14), .CI(co_Multiplier_0_2_2), 
           .COUT(co_Multiplier_0_2_3), .S0(s_Multiplier_0_2_13), .S1(s_Multiplier_0_2_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_2_4 (.A0(Multiplier_0_pp_4_15), .A1(Multiplier_0_pp_4_16), 
           .B0(Multiplier_0_pp_5_15), .B1(Multiplier_0_pp_5_16), .CI(co_Multiplier_0_2_3), 
           .COUT(co_Multiplier_0_2_4), .S0(s_Multiplier_0_2_15), .S1(s_Multiplier_0_2_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_2_5 (.A0(Multiplier_0_pp_4_17), .A1(Multiplier_0_pp_4_18), 
           .B0(Multiplier_0_pp_5_17), .B1(Multiplier_0_pp_5_18), .CI(co_Multiplier_0_2_4), 
           .COUT(co_Multiplier_0_2_5), .S0(s_Multiplier_0_2_17), .S1(s_Multiplier_0_2_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_2_6 (.A0(Multiplier_0_pp_4_19), .A1(Multiplier_0_pp_4_20), 
           .B0(Multiplier_0_pp_5_19), .B1(Multiplier_0_pp_5_20), .CI(co_Multiplier_0_2_5), 
           .COUT(co_Multiplier_0_2_6), .S0(s_Multiplier_0_2_19), .S1(s_Multiplier_0_2_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_2_7 (.A0(Multiplier_0_pp_4_21), .A1(GND_net), 
           .B0(Multiplier_0_pp_5_21), .B1(Multiplier_0_pp_5_22), .CI(co_Multiplier_0_2_6), 
           .COUT(co_Multiplier_0_2_7), .S0(s_Multiplier_0_2_21), .S1(s_Multiplier_0_2_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_2_8 (.A0(GND_net), .A1(GND_net), .B0(Multiplier_0_pp_5_23), 
           .B1(GND_net), .CI(co_Multiplier_0_2_7), .S0(s_Multiplier_0_2_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_Multiplier_0_3_1 (.A0(GND_net), .A1(f_s_Multiplier_0_0_4), 
           .B0(GND_net), .B1(f_Multiplier_0_pp_2_4), .CI(GND_net), .COUT(co_Multiplier_0_3_1), 
           .S1(rego_o_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_2 (.A0(f_s_Multiplier_0_0_5), .A1(f_s_Multiplier_0_0_6), 
           .B0(f_Multiplier_0_pp_2_5), .B1(f_s_Multiplier_0_1_6), .CI(co_Multiplier_0_3_1), 
           .COUT(co_Multiplier_0_3_2), .S0(rego_o_5), .S1(rego_o_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_3 (.A0(f_s_Multiplier_0_0_7), .A1(f_s_Multiplier_0_0_8), 
           .B0(f_s_Multiplier_0_1_7), .B1(f_s_Multiplier_0_1_8), .CI(co_Multiplier_0_3_2), 
           .COUT(co_Multiplier_0_3_3), .S0(rego_o_7), .S1(s_Multiplier_0_3_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_4 (.A0(f_s_Multiplier_0_0_9), .A1(f_s_Multiplier_0_0_10), 
           .B0(f_s_Multiplier_0_1_9), .B1(f_s_Multiplier_0_1_10), .CI(co_Multiplier_0_3_3), 
           .COUT(co_Multiplier_0_3_4), .S0(s_Multiplier_0_3_9), .S1(s_Multiplier_0_3_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_5 (.A0(f_s_Multiplier_0_0_11), .A1(f_s_Multiplier_0_0_12), 
           .B0(f_s_Multiplier_0_1_11), .B1(f_s_Multiplier_0_1_12), .CI(co_Multiplier_0_3_4), 
           .COUT(co_Multiplier_0_3_5), .S0(s_Multiplier_0_3_11), .S1(s_Multiplier_0_3_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_6 (.A0(f_s_Multiplier_0_0_13), .A1(f_s_Multiplier_0_0_14), 
           .B0(f_s_Multiplier_0_1_13), .B1(f_s_Multiplier_0_1_14), .CI(co_Multiplier_0_3_5), 
           .COUT(co_Multiplier_0_3_6), .S0(s_Multiplier_0_3_13), .S1(s_Multiplier_0_3_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_7 (.A0(f_s_Multiplier_0_0_15), .A1(f_s_Multiplier_0_0_16), 
           .B0(f_s_Multiplier_0_1_15), .B1(f_s_Multiplier_0_1_16), .CI(co_Multiplier_0_3_6), 
           .COUT(co_Multiplier_0_3_7), .S0(s_Multiplier_0_3_15), .S1(s_Multiplier_0_3_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_8 (.A0(f_s_Multiplier_0_0_17), .A1(GND_net), 
           .B0(f_s_Multiplier_0_1_17), .B1(f_s_Multiplier_0_1_18), .CI(co_Multiplier_0_3_7), 
           .COUT(co_Multiplier_0_3_8), .S0(s_Multiplier_0_3_17), .S1(s_Multiplier_0_3_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_9 (.A0(GND_net), .A1(GND_net), .B0(f_s_Multiplier_0_1_19), 
           .B1(f_s_Multiplier_0_1_20), .CI(co_Multiplier_0_3_8), .COUT(co_Multiplier_0_3_9), 
           .S0(s_Multiplier_0_3_19), .S1(s_Multiplier_0_3_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_10 (.A0(GND_net), .A1(GND_net), .B0(f_s_Multiplier_0_1_21), 
           .B1(GND_net), .CI(co_Multiplier_0_3_9), .COUT(co_Multiplier_0_3_10), 
           .S0(s_Multiplier_0_3_21), .S1(s_Multiplier_0_3_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_Multiplier_0_3_11 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_Multiplier_0_3_10), .S0(s_Multiplier_0_3_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_t_Multiplier_0_4_1 (.A0(GND_net), .A1(s_Multiplier_0_3_8), 
           .B0(GND_net), .B1(f_Multiplier_0_pp_4_8), .CI(GND_net), .COUT(co_t_Multiplier_0_4_1), 
           .S1(rego_o_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_2 (.A0(s_Multiplier_0_3_9), .A1(s_Multiplier_0_3_10), 
           .B0(f_Multiplier_0_pp_4_9), .B1(f_s_Multiplier_0_2_10), .CI(co_t_Multiplier_0_4_1), 
           .COUT(co_t_Multiplier_0_4_2), .S0(rego_o_9), .S1(rego_o_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_3 (.A0(s_Multiplier_0_3_11), .A1(s_Multiplier_0_3_12), 
           .B0(f_s_Multiplier_0_2_11), .B1(f_s_Multiplier_0_2_12), .CI(co_t_Multiplier_0_4_2), 
           .COUT(co_t_Multiplier_0_4_3), .S0(rego_o_11), .S1(rego_o_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_4 (.A0(s_Multiplier_0_3_13), .A1(s_Multiplier_0_3_14), 
           .B0(f_s_Multiplier_0_2_13), .B1(f_s_Multiplier_0_2_14), .CI(co_t_Multiplier_0_4_3), 
           .COUT(co_t_Multiplier_0_4_4), .S0(rego_o_13), .S1(rego_o_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_5 (.A0(s_Multiplier_0_3_15), .A1(s_Multiplier_0_3_16), 
           .B0(f_s_Multiplier_0_2_15), .B1(f_s_Multiplier_0_2_16), .CI(co_t_Multiplier_0_4_4), 
           .COUT(co_t_Multiplier_0_4_5), .S0(rego_o_15), .S1(rego_o_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_6 (.A0(s_Multiplier_0_3_17), .A1(s_Multiplier_0_3_18), 
           .B0(f_s_Multiplier_0_2_17), .B1(f_s_Multiplier_0_2_18), .CI(co_t_Multiplier_0_4_5), 
           .COUT(co_t_Multiplier_0_4_6), .S0(rego_o_17), .S1(rego_o_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_7 (.A0(s_Multiplier_0_3_19), .A1(s_Multiplier_0_3_20), 
           .B0(f_s_Multiplier_0_2_19), .B1(f_s_Multiplier_0_2_20), .CI(co_t_Multiplier_0_4_6), 
           .COUT(co_t_Multiplier_0_4_7), .S0(rego_o_19), .S1(rego_o_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_8 (.A0(s_Multiplier_0_3_21), .A1(s_Multiplier_0_3_22), 
           .B0(f_s_Multiplier_0_2_21), .B1(f_s_Multiplier_0_2_22), .CI(co_t_Multiplier_0_4_7), 
           .COUT(co_t_Multiplier_0_4_8), .S0(rego_o_21), .S1(rego_o_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_9 (.A0(s_Multiplier_0_3_23), .A1(GND_net), 
           .B0(f_s_Multiplier_0_2_23), .B1(GND_net), .CI(co_t_Multiplier_0_4_8), 
           .S0(rego_o_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_0_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(Multiplier_0_cin_lr_0), .CO(mco), .P0(Multiplier_0_pp_0_1), 
          .P1(Multiplier_0_pp_0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_0_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco), .CO(mco_1), .P0(Multiplier_0_pp_0_3), 
          .P1(Multiplier_0_pp_0_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_0_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco_1), .CO(mco_2), .P0(Multiplier_0_pp_0_5), 
          .P1(Multiplier_0_pp_0_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_0_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco_2), .CO(mco_3), .P0(Multiplier_0_pp_0_7), 
          .P1(Multiplier_0_pp_0_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_0_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco_3), .CO(mco_4), .P0(Multiplier_0_pp_0_9), 
          .P1(Multiplier_0_pp_0_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_0_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_0_5_n2), 
          .A2(Multiplier_0_mult_0_5_n1), .A3(VCC_net), .B0(regb_b_1), 
          .B1(VCC_net), .B2(VCC_net), .B3(VCC_net), .CI(mco_4), .CO(mfco), 
          .P0(Multiplier_0_pp_0_11), .P1(Multiplier_0_pp_0_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_2_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(Multiplier_0_cin_lr_2), .CO(mco_5), .P0(Multiplier_0_pp_1_3), 
          .P1(Multiplier_0_pp_1_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_2_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_5), .CO(mco_6), .P0(Multiplier_0_pp_1_5), 
          .P1(Multiplier_0_pp_1_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_2_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_6), .CO(mco_7), .P0(Multiplier_0_pp_1_7), 
          .P1(Multiplier_0_pp_1_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_2_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_7), .CO(mco_8), .P0(Multiplier_0_pp_1_9), 
          .P1(Multiplier_0_pp_1_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_2_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_8), .CO(mco_9), .P0(Multiplier_0_pp_1_11), 
          .P1(Multiplier_0_pp_1_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_2_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_2_5_n2), 
          .A2(Multiplier_0_mult_2_5_n1), .A3(GND_net), .B0(regb_b_3), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_2), .CI(mco_9), .CO(mfco_1), 
          .P0(Multiplier_0_pp_1_13), .P1(Multiplier_0_pp_1_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_4_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(Multiplier_0_cin_lr_4), .CO(mco_10), .P0(Multiplier_0_pp_2_5), 
          .P1(Multiplier_0_pp_2_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_4_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_10), .CO(mco_11), .P0(Multiplier_0_pp_2_7), 
          .P1(Multiplier_0_pp_2_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_4_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_11), .CO(mco_12), .P0(Multiplier_0_pp_2_9), 
          .P1(Multiplier_0_pp_2_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_4_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_12), .CO(mco_13), .P0(Multiplier_0_pp_2_11), 
          .P1(Multiplier_0_pp_2_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_4_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_13), .CO(mco_14), .P0(Multiplier_0_pp_2_13), 
          .P1(Multiplier_0_pp_2_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_4_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_4_5_n2), 
          .A2(Multiplier_0_mult_4_5_n1), .A3(GND_net), .B0(regb_b_5), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_4), .CI(mco_14), .CO(mfco_2), 
          .P0(Multiplier_0_pp_2_15), .P1(Multiplier_0_pp_2_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_6_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(Multiplier_0_cin_lr_6), .CO(mco_15), .P0(Multiplier_0_pp_3_7), 
          .P1(Multiplier_0_pp_3_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_6_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_15), .CO(mco_16), .P0(Multiplier_0_pp_3_9), 
          .P1(Multiplier_0_pp_3_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_6_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_16), .CO(mco_17), .P0(Multiplier_0_pp_3_11), 
          .P1(Multiplier_0_pp_3_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_6_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_17), .CO(mco_18), .P0(Multiplier_0_pp_3_13), 
          .P1(Multiplier_0_pp_3_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_6_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_18), .CO(mco_19), .P0(Multiplier_0_pp_3_15), 
          .P1(Multiplier_0_pp_3_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_6_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_6_5_n2), 
          .A2(Multiplier_0_mult_6_5_n1), .A3(GND_net), .B0(regb_b_7), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_6), .CI(mco_19), .CO(mfco_3), 
          .P0(Multiplier_0_pp_3_17), .P1(Multiplier_0_pp_3_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_8_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(Multiplier_0_cin_lr_8), .CO(mco_20), .P0(Multiplier_0_pp_4_9), 
          .P1(Multiplier_0_pp_4_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_8_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_20), .CO(mco_21), .P0(Multiplier_0_pp_4_11), 
          .P1(Multiplier_0_pp_4_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_8_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_21), .CO(mco_22), .P0(Multiplier_0_pp_4_13), 
          .P1(Multiplier_0_pp_4_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_8_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_22), .CO(mco_23), .P0(Multiplier_0_pp_4_15), 
          .P1(Multiplier_0_pp_4_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_8_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_23), .CO(mco_24), .P0(Multiplier_0_pp_4_17), 
          .P1(Multiplier_0_pp_4_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_8_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_8_5_n2), 
          .A2(Multiplier_0_mult_8_5_n1), .A3(GND_net), .B0(regb_b_9), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_8), .CI(mco_24), .CO(mfco_4), 
          .P0(Multiplier_0_pp_4_19), .P1(Multiplier_0_pp_4_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_10_0 (.A0(Multiplier_0_mult_10_0_n0), .A1(rega_a_1), 
          .A2(Multiplier_0_mult_10_0_n1), .A3(rega_a_2), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(Multiplier_0_cin_lr_10), 
          .CO(mco_25), .P0(Multiplier_0_pp_5_11), .P1(Multiplier_0_pp_5_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_10_1 (.A0(Multiplier_0_mult_10_1_n0), .A1(rega_a_3), 
          .A2(Multiplier_0_mult_10_1_n1), .A3(rega_a_4), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_25), 
          .CO(mco_26), .P0(Multiplier_0_pp_5_13), .P1(Multiplier_0_pp_5_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_10_2 (.A0(Multiplier_0_mult_10_2_n0), .A1(rega_a_5), 
          .A2(Multiplier_0_mult_10_2_n1), .A3(rega_a_6), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_26), 
          .CO(mco_27), .P0(Multiplier_0_pp_5_15), .P1(Multiplier_0_pp_5_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_10_3 (.A0(Multiplier_0_mult_10_3_n0), .A1(rega_a_7), 
          .A2(Multiplier_0_mult_10_3_n1), .A3(rega_a_8), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_27), 
          .CO(mco_28), .P0(Multiplier_0_pp_5_17), .P1(Multiplier_0_pp_5_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_10_4 (.A0(Multiplier_0_mult_10_4_n0), .A1(rega_a_9), 
          .A2(Multiplier_0_mult_10_4_n1), .A3(rega_a_10), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_28), 
          .CO(mco_29), .P0(Multiplier_0_pp_5_19), .P1(Multiplier_0_pp_5_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_10_5 (.A0(Multiplier_0_mult_10_5_n0), .A1(Multiplier_0_mult_10_5_n2), 
          .A2(rega_a_11), .A3(GND_net), .B0(VCC_net), .B1(VCC_net), 
          .B2(regb_b_11), .B3(regb_b_10), .CI(mco_29), .CO(mfco_5), 
          .P0(Multiplier_0_pp_5_21), .P1(Multiplier_0_pp_5_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    AND2 AND2_t27 (.A(regb_b_0), .B(regb_b_0), .Z(Multiplier_0_pp_0_0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(376[10:72])
    ND2 ND2_t26 (.A(rega_a_11), .B(regb_b_0), .Z(Multiplier_0_mult_0_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t23 (.A(rega_a_11), .B(regb_b_2), .Z(Multiplier_0_mult_2_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t20 (.A(rega_a_11), .B(regb_b_4), .Z(Multiplier_0_mult_4_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t17 (.A(rega_a_11), .B(regb_b_6), .Z(Multiplier_0_mult_6_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t14 (.A(rega_a_11), .B(regb_b_8), .Z(Multiplier_0_mult_8_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t11 (.A(rega_a_1), .B(regb_b_11), .Z(Multiplier_0_mult_10_0_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    
endmodule
//
// Verilog Description of module Multiplier_U0
//

module Multiplier_U0 (CIC1_out_clkSin, VCC_net, GND_net, MultDataB, 
            MultResult1) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input CIC1_out_clkSin;
    input VCC_net;
    input GND_net;
    input [11:0]MultDataB;
    output [23:0]MultResult1;
    
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(82[6:21])
    
    wire Multiplier_0_mult_0_5_n1, regb_b_1, rega_a_11, Multiplier_0_pp_1_2, 
        regb_b_2, regb_b_0, Multiplier_0_mult_2_5_n1, regb_b_3, Multiplier_0_pp_2_4, 
        regb_b_4, Multiplier_0_mult_4_5_n1, regb_b_5, Multiplier_0_pp_3_6, 
        regb_b_6, Multiplier_0_mult_6_5_n1, regb_b_7, Multiplier_0_pp_4_8, 
        regb_b_8, Multiplier_0_mult_8_5_n1, regb_b_9, Multiplier_0_pp_5_10, 
        regb_b_10, Multiplier_0_mult_10_0_n0, regb_b_11, Multiplier_0_mult_10_1_n1, 
        rega_a_3, rega_a_2, Multiplier_0_mult_10_1_n0, Multiplier_0_mult_10_2_n1, 
        rega_a_5, rega_a_4, Multiplier_0_mult_10_2_n0, Multiplier_0_mult_10_3_n1, 
        rega_a_7, rega_a_6, Multiplier_0_mult_10_3_n0, Multiplier_0_mult_10_4_n1, 
        rega_a_9, rega_a_8, Multiplier_0_mult_10_4_n0, Multiplier_0_mult_10_5_n2, 
        rega_a_10, Multiplier_0_mult_10_5_n0, rega_a_1, rego_o_0, rego_o_1, 
        rego_o_2, rego_o_3, rego_o_4, rego_o_5, rego_o_6, rego_o_7, 
        rego_o_8, rego_o_9, rego_o_10, rego_o_11, rego_o_12, rego_o_13, 
        rego_o_14, rego_o_15, rego_o_16, rego_o_17, rego_o_18, rego_o_19, 
        rego_o_20, rego_o_21, rego_o_22, rego_o_23, Multiplier_0_pp_0_0, 
        Multiplier_0_pp_0_1, s_Multiplier_0_0_2, s_Multiplier_0_0_3, s_Multiplier_0_0_4, 
        f_s_Multiplier_0_0_4, s_Multiplier_0_0_5, f_s_Multiplier_0_0_5, 
        s_Multiplier_0_0_6, f_s_Multiplier_0_0_6, s_Multiplier_0_0_7, 
        f_s_Multiplier_0_0_7, s_Multiplier_0_0_8, f_s_Multiplier_0_0_8, 
        s_Multiplier_0_0_9, f_s_Multiplier_0_0_9, s_Multiplier_0_0_10, 
        f_s_Multiplier_0_0_10, s_Multiplier_0_0_11, f_s_Multiplier_0_0_11, 
        s_Multiplier_0_0_12, f_s_Multiplier_0_0_12, s_Multiplier_0_0_13, 
        f_s_Multiplier_0_0_13, s_Multiplier_0_0_14, f_s_Multiplier_0_0_14, 
        s_Multiplier_0_0_15, f_s_Multiplier_0_0_15, s_Multiplier_0_0_16, 
        f_s_Multiplier_0_0_16, s_Multiplier_0_0_17, f_s_Multiplier_0_0_17, 
        f_Multiplier_0_pp_2_4, f_Multiplier_0_pp_2_5, Multiplier_0_pp_2_5, 
        s_Multiplier_0_1_6, f_s_Multiplier_0_1_6, s_Multiplier_0_1_7, 
        f_s_Multiplier_0_1_7, s_Multiplier_0_1_8, f_s_Multiplier_0_1_8, 
        s_Multiplier_0_1_9, f_s_Multiplier_0_1_9, s_Multiplier_0_1_10, 
        f_s_Multiplier_0_1_10, s_Multiplier_0_1_11, f_s_Multiplier_0_1_11, 
        s_Multiplier_0_1_12, f_s_Multiplier_0_1_12, s_Multiplier_0_1_13, 
        f_s_Multiplier_0_1_13, s_Multiplier_0_1_14, f_s_Multiplier_0_1_14, 
        s_Multiplier_0_1_15, f_s_Multiplier_0_1_15, s_Multiplier_0_1_16, 
        f_s_Multiplier_0_1_16, s_Multiplier_0_1_17, f_s_Multiplier_0_1_17, 
        s_Multiplier_0_1_18, f_s_Multiplier_0_1_18, s_Multiplier_0_1_19, 
        f_s_Multiplier_0_1_19, s_Multiplier_0_1_20, f_s_Multiplier_0_1_20, 
        s_Multiplier_0_1_21, f_s_Multiplier_0_1_21, f_Multiplier_0_pp_4_8, 
        f_Multiplier_0_pp_4_9, Multiplier_0_pp_4_9, s_Multiplier_0_2_10, 
        f_s_Multiplier_0_2_10, s_Multiplier_0_2_11, f_s_Multiplier_0_2_11, 
        s_Multiplier_0_2_12, f_s_Multiplier_0_2_12, s_Multiplier_0_2_13, 
        f_s_Multiplier_0_2_13, s_Multiplier_0_2_14, f_s_Multiplier_0_2_14, 
        s_Multiplier_0_2_15, f_s_Multiplier_0_2_15, s_Multiplier_0_2_16, 
        f_s_Multiplier_0_2_16, s_Multiplier_0_2_17, f_s_Multiplier_0_2_17, 
        s_Multiplier_0_2_18, f_s_Multiplier_0_2_18, s_Multiplier_0_2_19, 
        f_s_Multiplier_0_2_19, s_Multiplier_0_2_20, f_s_Multiplier_0_2_20, 
        s_Multiplier_0_2_21, f_s_Multiplier_0_2_21, s_Multiplier_0_2_22, 
        f_s_Multiplier_0_2_22, s_Multiplier_0_2_23, f_s_Multiplier_0_2_23, 
        Multiplier_0_cin_lr_0, Multiplier_0_pp_0_13, mfco, Multiplier_0_cin_lr_2, 
        Multiplier_0_pp_1_15, mfco_1, Multiplier_0_cin_lr_4, Multiplier_0_pp_2_17, 
        mfco_2, Multiplier_0_cin_lr_6, Multiplier_0_pp_3_19, mfco_3, 
        Multiplier_0_cin_lr_8, Multiplier_0_pp_4_21, mfco_4, Multiplier_0_cin_lr_10, 
        Multiplier_0_pp_5_23, mfco_5, co_Multiplier_0_0_1, Multiplier_0_pp_0_2, 
        co_Multiplier_0_0_2, Multiplier_0_pp_0_4, Multiplier_0_pp_0_3, 
        Multiplier_0_pp_1_4, Multiplier_0_pp_1_3, co_Multiplier_0_0_3, 
        Multiplier_0_pp_0_6, Multiplier_0_pp_0_5, Multiplier_0_pp_1_6, 
        Multiplier_0_pp_1_5, co_Multiplier_0_0_4, Multiplier_0_pp_0_8, 
        Multiplier_0_pp_0_7, Multiplier_0_pp_1_8, Multiplier_0_pp_1_7, 
        co_Multiplier_0_0_5, Multiplier_0_pp_0_10, Multiplier_0_pp_0_9, 
        Multiplier_0_pp_1_10, Multiplier_0_pp_1_9, co_Multiplier_0_0_6, 
        Multiplier_0_pp_0_12, Multiplier_0_pp_0_11, Multiplier_0_pp_1_12, 
        Multiplier_0_pp_1_11, co_Multiplier_0_0_7, Multiplier_0_pp_1_14, 
        Multiplier_0_pp_1_13, co_Multiplier_0_0_8, co_Multiplier_0_1_1, 
        Multiplier_0_pp_2_6, co_Multiplier_0_1_2, Multiplier_0_pp_2_8, 
        Multiplier_0_pp_2_7, Multiplier_0_pp_3_8, Multiplier_0_pp_3_7, 
        co_Multiplier_0_1_3, Multiplier_0_pp_2_10, Multiplier_0_pp_2_9, 
        Multiplier_0_pp_3_10, Multiplier_0_pp_3_9, co_Multiplier_0_1_4, 
        Multiplier_0_pp_2_12, Multiplier_0_pp_2_11, Multiplier_0_pp_3_12, 
        Multiplier_0_pp_3_11, co_Multiplier_0_1_5, Multiplier_0_pp_2_14, 
        Multiplier_0_pp_2_13, Multiplier_0_pp_3_14, Multiplier_0_pp_3_13, 
        co_Multiplier_0_1_6, Multiplier_0_pp_2_16, Multiplier_0_pp_2_15, 
        Multiplier_0_pp_3_16, Multiplier_0_pp_3_15, co_Multiplier_0_1_7, 
        Multiplier_0_pp_3_18, Multiplier_0_pp_3_17, co_Multiplier_0_1_8, 
        co_Multiplier_0_2_1, Multiplier_0_pp_4_10, co_Multiplier_0_2_2, 
        Multiplier_0_pp_4_12, Multiplier_0_pp_4_11, Multiplier_0_pp_5_12, 
        Multiplier_0_pp_5_11, co_Multiplier_0_2_3, Multiplier_0_pp_4_14, 
        Multiplier_0_pp_4_13, Multiplier_0_pp_5_14, Multiplier_0_pp_5_13, 
        co_Multiplier_0_2_4, Multiplier_0_pp_4_16, Multiplier_0_pp_4_15, 
        Multiplier_0_pp_5_16, Multiplier_0_pp_5_15, co_Multiplier_0_2_5, 
        Multiplier_0_pp_4_18, Multiplier_0_pp_4_17, Multiplier_0_pp_5_18, 
        Multiplier_0_pp_5_17, co_Multiplier_0_2_6, Multiplier_0_pp_4_20, 
        Multiplier_0_pp_4_19, Multiplier_0_pp_5_20, Multiplier_0_pp_5_19, 
        co_Multiplier_0_2_7, Multiplier_0_pp_5_22, Multiplier_0_pp_5_21, 
        co_Multiplier_0_3_1, co_Multiplier_0_3_2, co_Multiplier_0_3_3, 
        s_Multiplier_0_3_8, co_Multiplier_0_3_4, s_Multiplier_0_3_9, s_Multiplier_0_3_10, 
        co_Multiplier_0_3_5, s_Multiplier_0_3_11, s_Multiplier_0_3_12, 
        co_Multiplier_0_3_6, s_Multiplier_0_3_13, s_Multiplier_0_3_14, 
        co_Multiplier_0_3_7, s_Multiplier_0_3_15, s_Multiplier_0_3_16, 
        co_Multiplier_0_3_8, s_Multiplier_0_3_17, s_Multiplier_0_3_18, 
        co_Multiplier_0_3_9, s_Multiplier_0_3_19, s_Multiplier_0_3_20, 
        co_Multiplier_0_3_10, s_Multiplier_0_3_21, s_Multiplier_0_3_22, 
        s_Multiplier_0_3_23, co_t_Multiplier_0_4_1, co_t_Multiplier_0_4_2, 
        co_t_Multiplier_0_4_3, co_t_Multiplier_0_4_4, co_t_Multiplier_0_4_5, 
        co_t_Multiplier_0_4_6, co_t_Multiplier_0_4_7, co_t_Multiplier_0_4_8, 
        mco, mco_1, mco_2, mco_3, mco_4, Multiplier_0_mult_0_5_n2, 
        mco_5, mco_6, mco_7, mco_8, mco_9, Multiplier_0_mult_2_5_n2, 
        mco_10, mco_11, mco_12, mco_13, mco_14, Multiplier_0_mult_4_5_n2, 
        mco_15, mco_16, mco_17, mco_18, mco_19, Multiplier_0_mult_6_5_n2, 
        mco_20, mco_21, mco_22, mco_23, mco_24, Multiplier_0_mult_8_5_n2, 
        Multiplier_0_mult_10_0_n1, mco_25, mco_26, mco_27, mco_28, 
        mco_29;
    
    ND2 ND2_t25 (.A(rega_a_11), .B(regb_b_1), .Z(Multiplier_0_mult_0_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    AND2 AND2_t24 (.A(regb_b_0), .B(regb_b_2), .Z(Multiplier_0_pp_1_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(382[10:72])
    ND2 ND2_t22 (.A(rega_a_11), .B(regb_b_3), .Z(Multiplier_0_mult_2_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    AND2 AND2_t21 (.A(regb_b_0), .B(regb_b_4), .Z(Multiplier_0_pp_2_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(388[10:72])
    ND2 ND2_t19 (.A(rega_a_11), .B(regb_b_5), .Z(Multiplier_0_mult_4_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    AND2 AND2_t18 (.A(regb_b_0), .B(regb_b_6), .Z(Multiplier_0_pp_3_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(394[10:72])
    ND2 ND2_t16 (.A(rega_a_11), .B(regb_b_7), .Z(Multiplier_0_mult_6_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    AND2 AND2_t15 (.A(regb_b_0), .B(regb_b_8), .Z(Multiplier_0_pp_4_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(400[10:72])
    ND2 ND2_t13 (.A(rega_a_11), .B(regb_b_9), .Z(Multiplier_0_mult_8_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    AND2 AND2_t12 (.A(regb_b_0), .B(regb_b_10), .Z(Multiplier_0_pp_5_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(406[10:74])
    ND2 ND2_t10 (.A(regb_b_0), .B(regb_b_11), .Z(Multiplier_0_mult_10_0_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t9 (.A(rega_a_3), .B(regb_b_11), .Z(Multiplier_0_mult_10_1_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t8 (.A(rega_a_2), .B(regb_b_11), .Z(Multiplier_0_mult_10_1_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t7 (.A(rega_a_5), .B(regb_b_11), .Z(Multiplier_0_mult_10_2_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t6 (.A(rega_a_4), .B(regb_b_11), .Z(Multiplier_0_mult_10_2_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t5 (.A(rega_a_7), .B(regb_b_11), .Z(Multiplier_0_mult_10_3_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t4 (.A(rega_a_6), .B(regb_b_11), .Z(Multiplier_0_mult_10_3_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t3 (.A(rega_a_9), .B(regb_b_11), .Z(Multiplier_0_mult_10_4_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t2 (.A(rega_a_8), .B(regb_b_11), .Z(Multiplier_0_mult_10_4_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t1 (.A(rega_a_11), .B(regb_b_10), .Z(Multiplier_0_mult_10_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t0 (.A(rega_a_10), .B(regb_b_11), .Z(Multiplier_0_mult_10_5_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FD1P3DX FF_98 (.D(MultDataB[1]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(435[13:82])
    defparam FF_98.GSR = "ENABLED";
    FD1P3DX FF_97 (.D(MultDataB[2]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(438[13:82])
    defparam FF_97.GSR = "ENABLED";
    FD1P3DX FF_96 (.D(MultDataB[3]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(441[13:82])
    defparam FF_96.GSR = "ENABLED";
    FD1P3DX FF_95 (.D(MultDataB[4]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(444[13:82])
    defparam FF_95.GSR = "ENABLED";
    FD1P3DX FF_94 (.D(MultDataB[5]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(447[13:82])
    defparam FF_94.GSR = "ENABLED";
    FD1P3DX FF_93 (.D(MultDataB[6]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(450[13:82])
    defparam FF_93.GSR = "ENABLED";
    FD1P3DX FF_92 (.D(MultDataB[7]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(453[13:82])
    defparam FF_92.GSR = "ENABLED";
    FD1P3DX FF_91 (.D(MultDataB[8]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(456[13:82])
    defparam FF_91.GSR = "ENABLED";
    FD1P3DX FF_90 (.D(MultDataB[9]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(459[13:82])
    defparam FF_90.GSR = "ENABLED";
    FD1P3DX FF_89 (.D(MultDataB[10]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(462[13:84])
    defparam FF_89.GSR = "ENABLED";
    FD1P3DX FF_88 (.D(MultDataB[11]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(465[13:84])
    defparam FF_88.GSR = "ENABLED";
    FD1P3DX FF_87 (.D(MultDataB[0]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_0)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(468[13:82])
    defparam FF_87.GSR = "ENABLED";
    FD1P3DX FF_86 (.D(MultDataB[1]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(471[13:82])
    defparam FF_86.GSR = "ENABLED";
    FD1P3DX FF_85 (.D(MultDataB[2]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(474[13:82])
    defparam FF_85.GSR = "ENABLED";
    FD1P3DX FF_84 (.D(MultDataB[3]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(477[13:82])
    defparam FF_84.GSR = "ENABLED";
    FD1P3DX FF_83 (.D(MultDataB[4]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(480[13:82])
    defparam FF_83.GSR = "ENABLED";
    FD1P3DX FF_82 (.D(MultDataB[5]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(483[13:82])
    defparam FF_82.GSR = "ENABLED";
    FD1P3DX FF_81 (.D(MultDataB[6]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(486[13:82])
    defparam FF_81.GSR = "ENABLED";
    FD1P3DX FF_80 (.D(MultDataB[7]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(489[13:82])
    defparam FF_80.GSR = "ENABLED";
    FD1P3DX FF_79 (.D(MultDataB[8]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(492[13:82])
    defparam FF_79.GSR = "ENABLED";
    FD1P3DX FF_78 (.D(MultDataB[9]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(495[13:82])
    defparam FF_78.GSR = "ENABLED";
    FD1P3DX FF_77 (.D(MultDataB[10]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(498[13:84])
    defparam FF_77.GSR = "ENABLED";
    FD1P3DX FF_76 (.D(MultDataB[11]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(501[13:84])
    defparam FF_76.GSR = "ENABLED";
    FD1P3DX FF_75 (.D(rego_o_0), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[0])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(504[13:83])
    defparam FF_75.GSR = "ENABLED";
    FD1P3DX FF_74 (.D(rego_o_1), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[1])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(507[13:83])
    defparam FF_74.GSR = "ENABLED";
    FD1P3DX FF_73 (.D(rego_o_2), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[2])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(510[13:83])
    defparam FF_73.GSR = "ENABLED";
    FD1P3DX FF_72 (.D(rego_o_3), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[3])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(513[13:83])
    defparam FF_72.GSR = "ENABLED";
    FD1P3DX FF_71 (.D(rego_o_4), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[4])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(516[13:83])
    defparam FF_71.GSR = "ENABLED";
    FD1P3DX FF_70 (.D(rego_o_5), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[5])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(519[13:83])
    defparam FF_70.GSR = "ENABLED";
    FD1P3DX FF_69 (.D(rego_o_6), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[6])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(522[13:83])
    defparam FF_69.GSR = "ENABLED";
    FD1P3DX FF_68 (.D(rego_o_7), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[7])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(525[13:83])
    defparam FF_68.GSR = "ENABLED";
    FD1P3DX FF_67 (.D(rego_o_8), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[8])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(528[13:83])
    defparam FF_67.GSR = "ENABLED";
    FD1P3DX FF_66 (.D(rego_o_9), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[9])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(531[13:83])
    defparam FF_66.GSR = "ENABLED";
    FD1P3DX FF_65 (.D(rego_o_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[10])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(534[13:85])
    defparam FF_65.GSR = "ENABLED";
    FD1P3DX FF_64 (.D(rego_o_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[11])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(537[13:85])
    defparam FF_64.GSR = "ENABLED";
    FD1P3DX FF_63 (.D(rego_o_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[12])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(540[13:85])
    defparam FF_63.GSR = "ENABLED";
    FD1P3DX FF_62 (.D(rego_o_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[13])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(543[13:85])
    defparam FF_62.GSR = "ENABLED";
    FD1P3DX FF_61 (.D(rego_o_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[14])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(546[13:85])
    defparam FF_61.GSR = "ENABLED";
    FD1P3DX FF_60 (.D(rego_o_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[15])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(549[13:85])
    defparam FF_60.GSR = "ENABLED";
    FD1P3DX FF_59 (.D(rego_o_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[16])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(552[13:85])
    defparam FF_59.GSR = "ENABLED";
    FD1P3DX FF_58 (.D(rego_o_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[17])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(555[13:85])
    defparam FF_58.GSR = "ENABLED";
    FD1P3DX FF_57 (.D(rego_o_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[18])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(558[13:85])
    defparam FF_57.GSR = "ENABLED";
    FD1P3DX FF_56 (.D(rego_o_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[19])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(561[13:85])
    defparam FF_56.GSR = "ENABLED";
    FD1P3DX FF_55 (.D(rego_o_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[20])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(564[13:85])
    defparam FF_55.GSR = "ENABLED";
    FD1P3DX FF_54 (.D(rego_o_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[21])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(567[13:85])
    defparam FF_54.GSR = "ENABLED";
    FD1P3DX FF_53 (.D(rego_o_22), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[22])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(570[13:85])
    defparam FF_53.GSR = "ENABLED";
    FD1P3DX FF_52 (.D(rego_o_23), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[23])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(573[13:85])
    defparam FF_52.GSR = "ENABLED";
    FD1P3DX FF_51 (.D(Multiplier_0_pp_0_0), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_0)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(576[13] 577[35])
    defparam FF_51.GSR = "ENABLED";
    FD1P3DX FF_50 (.D(Multiplier_0_pp_0_1), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(580[13] 581[35])
    defparam FF_50.GSR = "ENABLED";
    FD1P3DX FF_49 (.D(s_Multiplier_0_0_2), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(584[13] 585[34])
    defparam FF_49.GSR = "ENABLED";
    FD1P3DX FF_48 (.D(s_Multiplier_0_0_3), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(588[13] 589[34])
    defparam FF_48.GSR = "ENABLED";
    FD1P3DX FF_47 (.D(s_Multiplier_0_0_4), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(592[13] 593[34])
    defparam FF_47.GSR = "ENABLED";
    FD1P3DX FF_46 (.D(s_Multiplier_0_0_5), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(596[13] 597[34])
    defparam FF_46.GSR = "ENABLED";
    FD1P3DX FF_45 (.D(s_Multiplier_0_0_6), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(600[13] 601[34])
    defparam FF_45.GSR = "ENABLED";
    FD1P3DX FF_44 (.D(s_Multiplier_0_0_7), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(604[13] 605[34])
    defparam FF_44.GSR = "ENABLED";
    FD1P3DX FF_43 (.D(s_Multiplier_0_0_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(608[13] 609[34])
    defparam FF_43.GSR = "ENABLED";
    FD1P3DX FF_42 (.D(s_Multiplier_0_0_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(612[13] 613[34])
    defparam FF_42.GSR = "ENABLED";
    FD1P3DX FF_41 (.D(s_Multiplier_0_0_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(616[13] 617[35])
    defparam FF_41.GSR = "ENABLED";
    FD1P3DX FF_40 (.D(s_Multiplier_0_0_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(620[13] 621[35])
    defparam FF_40.GSR = "ENABLED";
    FD1P3DX FF_39 (.D(s_Multiplier_0_0_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(624[13] 625[35])
    defparam FF_39.GSR = "ENABLED";
    FD1P3DX FF_38 (.D(s_Multiplier_0_0_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(628[13] 629[35])
    defparam FF_38.GSR = "ENABLED";
    FD1P3DX FF_37 (.D(s_Multiplier_0_0_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(632[13] 633[35])
    defparam FF_37.GSR = "ENABLED";
    FD1P3DX FF_36 (.D(s_Multiplier_0_0_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(636[13] 637[35])
    defparam FF_36.GSR = "ENABLED";
    FD1P3DX FF_35 (.D(s_Multiplier_0_0_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(640[13] 641[35])
    defparam FF_35.GSR = "ENABLED";
    FD1P3DX FF_34 (.D(s_Multiplier_0_0_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(644[13] 645[35])
    defparam FF_34.GSR = "ENABLED";
    FD1P3DX FF_33 (.D(Multiplier_0_pp_2_4), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_2_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(648[13] 649[35])
    defparam FF_33.GSR = "ENABLED";
    FD1P3DX FF_32 (.D(Multiplier_0_pp_2_5), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_2_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(652[13] 653[35])
    defparam FF_32.GSR = "ENABLED";
    FD1P3DX FF_31 (.D(s_Multiplier_0_1_6), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(656[13] 657[34])
    defparam FF_31.GSR = "ENABLED";
    FD1P3DX FF_30 (.D(s_Multiplier_0_1_7), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(660[13] 661[34])
    defparam FF_30.GSR = "ENABLED";
    FD1P3DX FF_29 (.D(s_Multiplier_0_1_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(664[13] 665[34])
    defparam FF_29.GSR = "ENABLED";
    FD1P3DX FF_28 (.D(s_Multiplier_0_1_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(668[13] 669[34])
    defparam FF_28.GSR = "ENABLED";
    FD1P3DX FF_27 (.D(s_Multiplier_0_1_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(672[13] 673[35])
    defparam FF_27.GSR = "ENABLED";
    FD1P3DX FF_26 (.D(s_Multiplier_0_1_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(676[13] 677[35])
    defparam FF_26.GSR = "ENABLED";
    FD1P3DX FF_25 (.D(s_Multiplier_0_1_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(680[13] 681[35])
    defparam FF_25.GSR = "ENABLED";
    FD1P3DX FF_24 (.D(s_Multiplier_0_1_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(684[13] 685[35])
    defparam FF_24.GSR = "ENABLED";
    FD1P3DX FF_23 (.D(s_Multiplier_0_1_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(688[13] 689[35])
    defparam FF_23.GSR = "ENABLED";
    FD1P3DX FF_22 (.D(s_Multiplier_0_1_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(692[13] 693[35])
    defparam FF_22.GSR = "ENABLED";
    FD1P3DX FF_21 (.D(s_Multiplier_0_1_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(696[13] 697[35])
    defparam FF_21.GSR = "ENABLED";
    FD1P3DX FF_20 (.D(s_Multiplier_0_1_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(700[13] 701[35])
    defparam FF_20.GSR = "ENABLED";
    FD1P3DX FF_19 (.D(s_Multiplier_0_1_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(704[13] 705[35])
    defparam FF_19.GSR = "ENABLED";
    FD1P3DX FF_18 (.D(s_Multiplier_0_1_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(708[13] 709[35])
    defparam FF_18.GSR = "ENABLED";
    FD1P3DX FF_17 (.D(s_Multiplier_0_1_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(712[13] 713[35])
    defparam FF_17.GSR = "ENABLED";
    FD1P3DX FF_16 (.D(s_Multiplier_0_1_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(716[13] 717[35])
    defparam FF_16.GSR = "ENABLED";
    FD1P3DX FF_15 (.D(Multiplier_0_pp_4_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_4_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(720[13] 721[35])
    defparam FF_15.GSR = "ENABLED";
    FD1P3DX FF_14 (.D(Multiplier_0_pp_4_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_4_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(724[13] 725[35])
    defparam FF_14.GSR = "ENABLED";
    FD1P3DX FF_13 (.D(s_Multiplier_0_2_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(728[13] 729[35])
    defparam FF_13.GSR = "ENABLED";
    FD1P3DX FF_12 (.D(s_Multiplier_0_2_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(732[13] 733[35])
    defparam FF_12.GSR = "ENABLED";
    FD1P3DX FF_11 (.D(s_Multiplier_0_2_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(736[13] 737[35])
    defparam FF_11.GSR = "ENABLED";
    FD1P3DX FF_10 (.D(s_Multiplier_0_2_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(740[13] 741[35])
    defparam FF_10.GSR = "ENABLED";
    FD1P3DX FF_9 (.D(s_Multiplier_0_2_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(744[13] 745[35])
    defparam FF_9.GSR = "ENABLED";
    FD1P3DX FF_8 (.D(s_Multiplier_0_2_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(748[13] 749[35])
    defparam FF_8.GSR = "ENABLED";
    FD1P3DX FF_7 (.D(s_Multiplier_0_2_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(752[13] 753[35])
    defparam FF_7.GSR = "ENABLED";
    FD1P3DX FF_6 (.D(s_Multiplier_0_2_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(756[13] 757[35])
    defparam FF_6.GSR = "ENABLED";
    FD1P3DX FF_5 (.D(s_Multiplier_0_2_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(760[13] 761[35])
    defparam FF_5.GSR = "ENABLED";
    FD1P3DX FF_4 (.D(s_Multiplier_0_2_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(764[13] 765[35])
    defparam FF_4.GSR = "ENABLED";
    FD1P3DX FF_3 (.D(s_Multiplier_0_2_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(768[13] 769[35])
    defparam FF_3.GSR = "ENABLED";
    FD1P3DX FF_2 (.D(s_Multiplier_0_2_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(772[13] 773[35])
    defparam FF_2.GSR = "ENABLED";
    FD1P3DX FF_1 (.D(s_Multiplier_0_2_22), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_22)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(776[13] 777[35])
    defparam FF_1.GSR = "ENABLED";
    FD1P3DX FF_0 (.D(s_Multiplier_0_2_23), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_23)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(780[13] 781[35])
    defparam FF_0.GSR = "ENABLED";
    FADD2B Multiplier_0_cin_lr_add_0 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_Cadd_0_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco), .S0(Multiplier_0_pp_0_13)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_cin_lr_add_2 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_Cadd_2_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_1), .S0(Multiplier_0_pp_1_15)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_cin_lr_add_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_Cadd_4_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_2), .S0(Multiplier_0_pp_2_17)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_cin_lr_add_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_Cadd_6_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_3), .S0(Multiplier_0_pp_3_19)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_cin_lr_add_8 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_Cadd_8_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_4), .S0(Multiplier_0_pp_4_21)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_cin_lr_add_10 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_Cadd_10_6 (.A0(VCC_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_5), .S0(Multiplier_0_pp_5_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_Multiplier_0_0_1 (.A0(GND_net), .A1(Multiplier_0_pp_0_2), 
           .B0(GND_net), .B1(Multiplier_0_pp_1_2), .CI(GND_net), .COUT(co_Multiplier_0_0_1), 
           .S1(s_Multiplier_0_0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_0_2 (.A0(Multiplier_0_pp_0_3), .A1(Multiplier_0_pp_0_4), 
           .B0(Multiplier_0_pp_1_3), .B1(Multiplier_0_pp_1_4), .CI(co_Multiplier_0_0_1), 
           .COUT(co_Multiplier_0_0_2), .S0(s_Multiplier_0_0_3), .S1(s_Multiplier_0_0_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_0_3 (.A0(Multiplier_0_pp_0_5), .A1(Multiplier_0_pp_0_6), 
           .B0(Multiplier_0_pp_1_5), .B1(Multiplier_0_pp_1_6), .CI(co_Multiplier_0_0_2), 
           .COUT(co_Multiplier_0_0_3), .S0(s_Multiplier_0_0_5), .S1(s_Multiplier_0_0_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_0_4 (.A0(Multiplier_0_pp_0_7), .A1(Multiplier_0_pp_0_8), 
           .B0(Multiplier_0_pp_1_7), .B1(Multiplier_0_pp_1_8), .CI(co_Multiplier_0_0_3), 
           .COUT(co_Multiplier_0_0_4), .S0(s_Multiplier_0_0_7), .S1(s_Multiplier_0_0_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_0_5 (.A0(Multiplier_0_pp_0_9), .A1(Multiplier_0_pp_0_10), 
           .B0(Multiplier_0_pp_1_9), .B1(Multiplier_0_pp_1_10), .CI(co_Multiplier_0_0_4), 
           .COUT(co_Multiplier_0_0_5), .S0(s_Multiplier_0_0_9), .S1(s_Multiplier_0_0_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_0_6 (.A0(Multiplier_0_pp_0_11), .A1(Multiplier_0_pp_0_12), 
           .B0(Multiplier_0_pp_1_11), .B1(Multiplier_0_pp_1_12), .CI(co_Multiplier_0_0_5), 
           .COUT(co_Multiplier_0_0_6), .S0(s_Multiplier_0_0_11), .S1(s_Multiplier_0_0_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_0_7 (.A0(Multiplier_0_pp_0_13), .A1(GND_net), 
           .B0(Multiplier_0_pp_1_13), .B1(Multiplier_0_pp_1_14), .CI(co_Multiplier_0_0_6), 
           .COUT(co_Multiplier_0_0_7), .S0(s_Multiplier_0_0_13), .S1(s_Multiplier_0_0_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_0_8 (.A0(GND_net), .A1(GND_net), .B0(Multiplier_0_pp_1_15), 
           .B1(GND_net), .CI(co_Multiplier_0_0_7), .COUT(co_Multiplier_0_0_8), 
           .S0(s_Multiplier_0_0_15), .S1(s_Multiplier_0_0_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_Multiplier_0_0_9 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_Multiplier_0_0_8), .S0(s_Multiplier_0_0_17)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_Multiplier_0_1_1 (.A0(GND_net), .A1(Multiplier_0_pp_2_6), 
           .B0(GND_net), .B1(Multiplier_0_pp_3_6), .CI(GND_net), .COUT(co_Multiplier_0_1_1), 
           .S1(s_Multiplier_0_1_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_1_2 (.A0(Multiplier_0_pp_2_7), .A1(Multiplier_0_pp_2_8), 
           .B0(Multiplier_0_pp_3_7), .B1(Multiplier_0_pp_3_8), .CI(co_Multiplier_0_1_1), 
           .COUT(co_Multiplier_0_1_2), .S0(s_Multiplier_0_1_7), .S1(s_Multiplier_0_1_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_1_3 (.A0(Multiplier_0_pp_2_9), .A1(Multiplier_0_pp_2_10), 
           .B0(Multiplier_0_pp_3_9), .B1(Multiplier_0_pp_3_10), .CI(co_Multiplier_0_1_2), 
           .COUT(co_Multiplier_0_1_3), .S0(s_Multiplier_0_1_9), .S1(s_Multiplier_0_1_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_1_4 (.A0(Multiplier_0_pp_2_11), .A1(Multiplier_0_pp_2_12), 
           .B0(Multiplier_0_pp_3_11), .B1(Multiplier_0_pp_3_12), .CI(co_Multiplier_0_1_3), 
           .COUT(co_Multiplier_0_1_4), .S0(s_Multiplier_0_1_11), .S1(s_Multiplier_0_1_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_1_5 (.A0(Multiplier_0_pp_2_13), .A1(Multiplier_0_pp_2_14), 
           .B0(Multiplier_0_pp_3_13), .B1(Multiplier_0_pp_3_14), .CI(co_Multiplier_0_1_4), 
           .COUT(co_Multiplier_0_1_5), .S0(s_Multiplier_0_1_13), .S1(s_Multiplier_0_1_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_1_6 (.A0(Multiplier_0_pp_2_15), .A1(Multiplier_0_pp_2_16), 
           .B0(Multiplier_0_pp_3_15), .B1(Multiplier_0_pp_3_16), .CI(co_Multiplier_0_1_5), 
           .COUT(co_Multiplier_0_1_6), .S0(s_Multiplier_0_1_15), .S1(s_Multiplier_0_1_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_1_7 (.A0(Multiplier_0_pp_2_17), .A1(GND_net), 
           .B0(Multiplier_0_pp_3_17), .B1(Multiplier_0_pp_3_18), .CI(co_Multiplier_0_1_6), 
           .COUT(co_Multiplier_0_1_7), .S0(s_Multiplier_0_1_17), .S1(s_Multiplier_0_1_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_1_8 (.A0(GND_net), .A1(GND_net), .B0(Multiplier_0_pp_3_19), 
           .B1(GND_net), .CI(co_Multiplier_0_1_7), .COUT(co_Multiplier_0_1_8), 
           .S0(s_Multiplier_0_1_19), .S1(s_Multiplier_0_1_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_Multiplier_0_1_9 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_Multiplier_0_1_8), .S0(s_Multiplier_0_1_21)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_Multiplier_0_2_1 (.A0(GND_net), .A1(Multiplier_0_pp_4_10), 
           .B0(GND_net), .B1(Multiplier_0_pp_5_10), .CI(GND_net), .COUT(co_Multiplier_0_2_1), 
           .S1(s_Multiplier_0_2_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_2_2 (.A0(Multiplier_0_pp_4_11), .A1(Multiplier_0_pp_4_12), 
           .B0(Multiplier_0_pp_5_11), .B1(Multiplier_0_pp_5_12), .CI(co_Multiplier_0_2_1), 
           .COUT(co_Multiplier_0_2_2), .S0(s_Multiplier_0_2_11), .S1(s_Multiplier_0_2_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_2_3 (.A0(Multiplier_0_pp_4_13), .A1(Multiplier_0_pp_4_14), 
           .B0(Multiplier_0_pp_5_13), .B1(Multiplier_0_pp_5_14), .CI(co_Multiplier_0_2_2), 
           .COUT(co_Multiplier_0_2_3), .S0(s_Multiplier_0_2_13), .S1(s_Multiplier_0_2_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_2_4 (.A0(Multiplier_0_pp_4_15), .A1(Multiplier_0_pp_4_16), 
           .B0(Multiplier_0_pp_5_15), .B1(Multiplier_0_pp_5_16), .CI(co_Multiplier_0_2_3), 
           .COUT(co_Multiplier_0_2_4), .S0(s_Multiplier_0_2_15), .S1(s_Multiplier_0_2_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_2_5 (.A0(Multiplier_0_pp_4_17), .A1(Multiplier_0_pp_4_18), 
           .B0(Multiplier_0_pp_5_17), .B1(Multiplier_0_pp_5_18), .CI(co_Multiplier_0_2_4), 
           .COUT(co_Multiplier_0_2_5), .S0(s_Multiplier_0_2_17), .S1(s_Multiplier_0_2_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_2_6 (.A0(Multiplier_0_pp_4_19), .A1(Multiplier_0_pp_4_20), 
           .B0(Multiplier_0_pp_5_19), .B1(Multiplier_0_pp_5_20), .CI(co_Multiplier_0_2_5), 
           .COUT(co_Multiplier_0_2_6), .S0(s_Multiplier_0_2_19), .S1(s_Multiplier_0_2_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_2_7 (.A0(Multiplier_0_pp_4_21), .A1(GND_net), 
           .B0(Multiplier_0_pp_5_21), .B1(Multiplier_0_pp_5_22), .CI(co_Multiplier_0_2_6), 
           .COUT(co_Multiplier_0_2_7), .S0(s_Multiplier_0_2_21), .S1(s_Multiplier_0_2_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_2_8 (.A0(GND_net), .A1(GND_net), .B0(Multiplier_0_pp_5_23), 
           .B1(GND_net), .CI(co_Multiplier_0_2_7), .S0(s_Multiplier_0_2_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_Multiplier_0_3_1 (.A0(GND_net), .A1(f_s_Multiplier_0_0_4), 
           .B0(GND_net), .B1(f_Multiplier_0_pp_2_4), .CI(GND_net), .COUT(co_Multiplier_0_3_1), 
           .S1(rego_o_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_2 (.A0(f_s_Multiplier_0_0_5), .A1(f_s_Multiplier_0_0_6), 
           .B0(f_Multiplier_0_pp_2_5), .B1(f_s_Multiplier_0_1_6), .CI(co_Multiplier_0_3_1), 
           .COUT(co_Multiplier_0_3_2), .S0(rego_o_5), .S1(rego_o_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_3 (.A0(f_s_Multiplier_0_0_7), .A1(f_s_Multiplier_0_0_8), 
           .B0(f_s_Multiplier_0_1_7), .B1(f_s_Multiplier_0_1_8), .CI(co_Multiplier_0_3_2), 
           .COUT(co_Multiplier_0_3_3), .S0(rego_o_7), .S1(s_Multiplier_0_3_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_4 (.A0(f_s_Multiplier_0_0_9), .A1(f_s_Multiplier_0_0_10), 
           .B0(f_s_Multiplier_0_1_9), .B1(f_s_Multiplier_0_1_10), .CI(co_Multiplier_0_3_3), 
           .COUT(co_Multiplier_0_3_4), .S0(s_Multiplier_0_3_9), .S1(s_Multiplier_0_3_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_5 (.A0(f_s_Multiplier_0_0_11), .A1(f_s_Multiplier_0_0_12), 
           .B0(f_s_Multiplier_0_1_11), .B1(f_s_Multiplier_0_1_12), .CI(co_Multiplier_0_3_4), 
           .COUT(co_Multiplier_0_3_5), .S0(s_Multiplier_0_3_11), .S1(s_Multiplier_0_3_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_6 (.A0(f_s_Multiplier_0_0_13), .A1(f_s_Multiplier_0_0_14), 
           .B0(f_s_Multiplier_0_1_13), .B1(f_s_Multiplier_0_1_14), .CI(co_Multiplier_0_3_5), 
           .COUT(co_Multiplier_0_3_6), .S0(s_Multiplier_0_3_13), .S1(s_Multiplier_0_3_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_7 (.A0(f_s_Multiplier_0_0_15), .A1(f_s_Multiplier_0_0_16), 
           .B0(f_s_Multiplier_0_1_15), .B1(f_s_Multiplier_0_1_16), .CI(co_Multiplier_0_3_6), 
           .COUT(co_Multiplier_0_3_7), .S0(s_Multiplier_0_3_15), .S1(s_Multiplier_0_3_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_8 (.A0(f_s_Multiplier_0_0_17), .A1(GND_net), 
           .B0(f_s_Multiplier_0_1_17), .B1(f_s_Multiplier_0_1_18), .CI(co_Multiplier_0_3_7), 
           .COUT(co_Multiplier_0_3_8), .S0(s_Multiplier_0_3_17), .S1(s_Multiplier_0_3_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_9 (.A0(GND_net), .A1(GND_net), .B0(f_s_Multiplier_0_1_19), 
           .B1(f_s_Multiplier_0_1_20), .CI(co_Multiplier_0_3_8), .COUT(co_Multiplier_0_3_9), 
           .S0(s_Multiplier_0_3_19), .S1(s_Multiplier_0_3_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_10 (.A0(GND_net), .A1(GND_net), .B0(f_s_Multiplier_0_1_21), 
           .B1(GND_net), .CI(co_Multiplier_0_3_9), .COUT(co_Multiplier_0_3_10), 
           .S0(s_Multiplier_0_3_21), .S1(s_Multiplier_0_3_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_Multiplier_0_3_11 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_Multiplier_0_3_10), .S0(s_Multiplier_0_3_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_t_Multiplier_0_4_1 (.A0(GND_net), .A1(s_Multiplier_0_3_8), 
           .B0(GND_net), .B1(f_Multiplier_0_pp_4_8), .CI(GND_net), .COUT(co_t_Multiplier_0_4_1), 
           .S1(rego_o_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_2 (.A0(s_Multiplier_0_3_9), .A1(s_Multiplier_0_3_10), 
           .B0(f_Multiplier_0_pp_4_9), .B1(f_s_Multiplier_0_2_10), .CI(co_t_Multiplier_0_4_1), 
           .COUT(co_t_Multiplier_0_4_2), .S0(rego_o_9), .S1(rego_o_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_3 (.A0(s_Multiplier_0_3_11), .A1(s_Multiplier_0_3_12), 
           .B0(f_s_Multiplier_0_2_11), .B1(f_s_Multiplier_0_2_12), .CI(co_t_Multiplier_0_4_2), 
           .COUT(co_t_Multiplier_0_4_3), .S0(rego_o_11), .S1(rego_o_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_4 (.A0(s_Multiplier_0_3_13), .A1(s_Multiplier_0_3_14), 
           .B0(f_s_Multiplier_0_2_13), .B1(f_s_Multiplier_0_2_14), .CI(co_t_Multiplier_0_4_3), 
           .COUT(co_t_Multiplier_0_4_4), .S0(rego_o_13), .S1(rego_o_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_5 (.A0(s_Multiplier_0_3_15), .A1(s_Multiplier_0_3_16), 
           .B0(f_s_Multiplier_0_2_15), .B1(f_s_Multiplier_0_2_16), .CI(co_t_Multiplier_0_4_4), 
           .COUT(co_t_Multiplier_0_4_5), .S0(rego_o_15), .S1(rego_o_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_6 (.A0(s_Multiplier_0_3_17), .A1(s_Multiplier_0_3_18), 
           .B0(f_s_Multiplier_0_2_17), .B1(f_s_Multiplier_0_2_18), .CI(co_t_Multiplier_0_4_5), 
           .COUT(co_t_Multiplier_0_4_6), .S0(rego_o_17), .S1(rego_o_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_7 (.A0(s_Multiplier_0_3_19), .A1(s_Multiplier_0_3_20), 
           .B0(f_s_Multiplier_0_2_19), .B1(f_s_Multiplier_0_2_20), .CI(co_t_Multiplier_0_4_6), 
           .COUT(co_t_Multiplier_0_4_7), .S0(rego_o_19), .S1(rego_o_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_8 (.A0(s_Multiplier_0_3_21), .A1(s_Multiplier_0_3_22), 
           .B0(f_s_Multiplier_0_2_21), .B1(f_s_Multiplier_0_2_22), .CI(co_t_Multiplier_0_4_7), 
           .COUT(co_t_Multiplier_0_4_8), .S0(rego_o_21), .S1(rego_o_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_9 (.A0(s_Multiplier_0_3_23), .A1(GND_net), 
           .B0(f_s_Multiplier_0_2_23), .B1(GND_net), .CI(co_t_Multiplier_0_4_8), 
           .S0(rego_o_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_0_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(Multiplier_0_cin_lr_0), .CO(mco), .P0(Multiplier_0_pp_0_1), 
          .P1(Multiplier_0_pp_0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_0_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco), .CO(mco_1), .P0(Multiplier_0_pp_0_3), 
          .P1(Multiplier_0_pp_0_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_0_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco_1), .CO(mco_2), .P0(Multiplier_0_pp_0_5), 
          .P1(Multiplier_0_pp_0_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_0_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco_2), .CO(mco_3), .P0(Multiplier_0_pp_0_7), 
          .P1(Multiplier_0_pp_0_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_0_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco_3), .CO(mco_4), .P0(Multiplier_0_pp_0_9), 
          .P1(Multiplier_0_pp_0_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_0_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_0_5_n2), 
          .A2(Multiplier_0_mult_0_5_n1), .A3(VCC_net), .B0(regb_b_1), 
          .B1(VCC_net), .B2(VCC_net), .B3(VCC_net), .CI(mco_4), .CO(mfco), 
          .P0(Multiplier_0_pp_0_11), .P1(Multiplier_0_pp_0_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_2_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(Multiplier_0_cin_lr_2), .CO(mco_5), .P0(Multiplier_0_pp_1_3), 
          .P1(Multiplier_0_pp_1_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_2_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_5), .CO(mco_6), .P0(Multiplier_0_pp_1_5), 
          .P1(Multiplier_0_pp_1_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_2_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_6), .CO(mco_7), .P0(Multiplier_0_pp_1_7), 
          .P1(Multiplier_0_pp_1_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_2_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_7), .CO(mco_8), .P0(Multiplier_0_pp_1_9), 
          .P1(Multiplier_0_pp_1_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_2_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_8), .CO(mco_9), .P0(Multiplier_0_pp_1_11), 
          .P1(Multiplier_0_pp_1_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_2_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_2_5_n2), 
          .A2(Multiplier_0_mult_2_5_n1), .A3(GND_net), .B0(regb_b_3), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_2), .CI(mco_9), .CO(mfco_1), 
          .P0(Multiplier_0_pp_1_13), .P1(Multiplier_0_pp_1_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_4_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(Multiplier_0_cin_lr_4), .CO(mco_10), .P0(Multiplier_0_pp_2_5), 
          .P1(Multiplier_0_pp_2_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_4_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_10), .CO(mco_11), .P0(Multiplier_0_pp_2_7), 
          .P1(Multiplier_0_pp_2_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_4_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_11), .CO(mco_12), .P0(Multiplier_0_pp_2_9), 
          .P1(Multiplier_0_pp_2_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_4_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_12), .CO(mco_13), .P0(Multiplier_0_pp_2_11), 
          .P1(Multiplier_0_pp_2_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_4_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_13), .CO(mco_14), .P0(Multiplier_0_pp_2_13), 
          .P1(Multiplier_0_pp_2_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_4_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_4_5_n2), 
          .A2(Multiplier_0_mult_4_5_n1), .A3(GND_net), .B0(regb_b_5), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_4), .CI(mco_14), .CO(mfco_2), 
          .P0(Multiplier_0_pp_2_15), .P1(Multiplier_0_pp_2_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_6_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(Multiplier_0_cin_lr_6), .CO(mco_15), .P0(Multiplier_0_pp_3_7), 
          .P1(Multiplier_0_pp_3_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_6_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_15), .CO(mco_16), .P0(Multiplier_0_pp_3_9), 
          .P1(Multiplier_0_pp_3_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_6_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_16), .CO(mco_17), .P0(Multiplier_0_pp_3_11), 
          .P1(Multiplier_0_pp_3_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_6_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_17), .CO(mco_18), .P0(Multiplier_0_pp_3_13), 
          .P1(Multiplier_0_pp_3_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_6_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_18), .CO(mco_19), .P0(Multiplier_0_pp_3_15), 
          .P1(Multiplier_0_pp_3_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_6_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_6_5_n2), 
          .A2(Multiplier_0_mult_6_5_n1), .A3(GND_net), .B0(regb_b_7), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_6), .CI(mco_19), .CO(mfco_3), 
          .P0(Multiplier_0_pp_3_17), .P1(Multiplier_0_pp_3_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_8_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(Multiplier_0_cin_lr_8), .CO(mco_20), .P0(Multiplier_0_pp_4_9), 
          .P1(Multiplier_0_pp_4_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_8_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_20), .CO(mco_21), .P0(Multiplier_0_pp_4_11), 
          .P1(Multiplier_0_pp_4_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_8_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_21), .CO(mco_22), .P0(Multiplier_0_pp_4_13), 
          .P1(Multiplier_0_pp_4_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_8_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_22), .CO(mco_23), .P0(Multiplier_0_pp_4_15), 
          .P1(Multiplier_0_pp_4_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_8_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_23), .CO(mco_24), .P0(Multiplier_0_pp_4_17), 
          .P1(Multiplier_0_pp_4_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_8_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_8_5_n2), 
          .A2(Multiplier_0_mult_8_5_n1), .A3(GND_net), .B0(regb_b_9), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_8), .CI(mco_24), .CO(mfco_4), 
          .P0(Multiplier_0_pp_4_19), .P1(Multiplier_0_pp_4_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_10_0 (.A0(Multiplier_0_mult_10_0_n0), .A1(rega_a_1), 
          .A2(Multiplier_0_mult_10_0_n1), .A3(rega_a_2), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(Multiplier_0_cin_lr_10), 
          .CO(mco_25), .P0(Multiplier_0_pp_5_11), .P1(Multiplier_0_pp_5_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_10_1 (.A0(Multiplier_0_mult_10_1_n0), .A1(rega_a_3), 
          .A2(Multiplier_0_mult_10_1_n1), .A3(rega_a_4), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_25), 
          .CO(mco_26), .P0(Multiplier_0_pp_5_13), .P1(Multiplier_0_pp_5_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_10_2 (.A0(Multiplier_0_mult_10_2_n0), .A1(rega_a_5), 
          .A2(Multiplier_0_mult_10_2_n1), .A3(rega_a_6), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_26), 
          .CO(mco_27), .P0(Multiplier_0_pp_5_15), .P1(Multiplier_0_pp_5_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_10_3 (.A0(Multiplier_0_mult_10_3_n0), .A1(rega_a_7), 
          .A2(Multiplier_0_mult_10_3_n1), .A3(rega_a_8), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_27), 
          .CO(mco_28), .P0(Multiplier_0_pp_5_17), .P1(Multiplier_0_pp_5_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_10_4 (.A0(Multiplier_0_mult_10_4_n0), .A1(rega_a_9), 
          .A2(Multiplier_0_mult_10_4_n1), .A3(rega_a_10), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_28), 
          .CO(mco_29), .P0(Multiplier_0_pp_5_19), .P1(Multiplier_0_pp_5_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_10_5 (.A0(Multiplier_0_mult_10_5_n0), .A1(Multiplier_0_mult_10_5_n2), 
          .A2(rega_a_11), .A3(GND_net), .B0(VCC_net), .B1(VCC_net), 
          .B2(regb_b_11), .B3(regb_b_10), .CI(mco_29), .CO(mfco_5), 
          .P0(Multiplier_0_pp_5_21), .P1(Multiplier_0_pp_5_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t26 (.A(rega_a_11), .B(regb_b_0), .Z(Multiplier_0_mult_0_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    AND2 AND2_t27 (.A(regb_b_0), .B(regb_b_0), .Z(Multiplier_0_pp_0_0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(376[10:72])
    ND2 ND2_t23 (.A(rega_a_11), .B(regb_b_2), .Z(Multiplier_0_mult_2_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t20 (.A(rega_a_11), .B(regb_b_4), .Z(Multiplier_0_mult_4_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t17 (.A(rega_a_11), .B(regb_b_6), .Z(Multiplier_0_mult_6_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t14 (.A(rega_a_11), .B(regb_b_8), .Z(Multiplier_0_mult_8_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t11 (.A(rega_a_1), .B(regb_b_11), .Z(Multiplier_0_mult_10_0_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=10, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    
endmodule
