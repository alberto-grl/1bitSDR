// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.11.2.446
// Netlist written on Sun Apr 05 20:40:24 2020
//
// Verilog Description of module top
//

module top (i_Rx_Serial, o_Tx_Serial, o_Rx_DV, o_Rx_Byte, MYLED, XIn, 
            XOut, RFIn, DiffOut, PWMOut, sinGen, sin_out, CIC_out_clkSin) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(38[8:11])
    input i_Rx_Serial;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(40[13:24])
    output o_Tx_Serial;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(42[11:22])
    output o_Rx_DV;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(43[13:20])
    output [7:0]o_Rx_Byte;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(44[16:25])
    output [7:0]MYLED;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(45[18:23])
    input XIn;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(46[8:11])
    output XOut;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(47[9:13])
    input RFIn;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(48[9:13])
    output DiffOut;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(49[9:16])
    output PWMOut;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[9:15])
    output sinGen;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(51[9:15])
    output sin_out;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(52[9:16])
    output CIC_out_clkSin;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(53[9:23])
    
    wire XIn_c /* synthesis is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(46[8:11])
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(55[8:15])
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(67[6:21])
    wire [7:0]UartClk_adj_2711 /* synthesis SET_AS_NETWORK=\uart_tx1/UartClk[2], is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(37[14:21])
    
    wire GND_net, VCC_net, i_Rx_Serial_c, o_Tx_Serial_c, o_Rx_Byte_c_7, 
        o_Rx_Byte_c_6, o_Rx_Byte_c_5, o_Rx_Byte_c_4, o_Rx_Byte_c_3, 
        o_Rx_Byte_c_2, n7319, o_Rx_Byte_c_0, MYLED_c_5, MYLED_c_4, 
        MYLED_c_3, MYLED_c_2, MYLED_c_1, MYLED_c_0, RFIn_c, DiffOut_c, 
        PWMOut_c, sinGen_c, n2244;
    wire [11:0]MixerOutSin;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(63[20:31])
    wire [11:0]MixerOutCos;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(64[20:31])
    wire [11:0]CIC1_outSin;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(66[20:31])
    wire [11:0]CIC1_outCos;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(69[20:31])
    wire [63:0]phase_accum;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(71[13:24])
    wire [12:0]LOSine;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(72[20:26])
    wire [12:0]LOCosine;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(73[20:28])
    wire [63:0]phase_inc_carrGen;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(75[19:36])
    wire [63:0]phase_inc_carrGen1;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(76[19:37])
    wire [11:0]DemodOut;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(79[20:28])
    wire [7:0]CICGain;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(81[11:18])
    
    wire n1003, n1002, n1001, n1000, n999, n998, n997, n996, 
        n995, n994, n993, n992, n991, n990, n989, n988, n987, 
        n986, n985, n984, n983, n982, n981, n980, n979, n978, 
        n977, n976, n975, n974, n973, n972, n971, n970, n969, 
        n968, n967, n966, n965, n964, n963, n962, n961, n960, 
        n959, n958, n957, n956, n955, n954, n953, n952, n951, 
        n950, n949, n948, n947, n946, n945, n943, n944, n13804, 
        n2335, n2331, n2330, n2316, n2314, n2310, n2309, n881, 
        n880, n882, n883, n884, n885, n886, n887, n888, n889, 
        n890, n891, n892, n893, n894, n895, n896, n897, n898, 
        n899, n900, n901, n902, n903, n904, n905, n906, n907, 
        n908, n909, n910, n911, n912, n913, n914, n915, n916, 
        n917, n918, n919, n920, n921, n922, n923, n924, n925, 
        n926, n927, n928, n929, n930, n931, n932, n933, n934, 
        n935, n936, n937, n938, n939, n940, n941, n2601, n2600, 
        n2728, n2727, n2301, n2249, n11611, n11610, n11609, n11608, 
        n11607, n11606, n11605, n13822, n11604, n11603, n11602, 
        n11601, n11600, n11599, n11598, n11597, n11596, n11595, 
        n11594, n11593, n11592, n11591, n11590, n11589, n11588, 
        n11587, n11586, n11585, n11584, n11583, n11582, n11581, 
        n11579, n11578, n11577, n11576, n11575, n11574, n11573, 
        n11572, n11571, n11570, n11569, n11568, n11567, n11566, 
        n11565, n11564, n11563, n11562, n11561, n11560, n11559, 
        n11558, n11557, n11556, n11555, n11554, n11553, n11552, 
        n11551, n11550, n2299, n2725;
    wire [71:0]d10_adj_2639;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(47[26:29])
    
    wire n2248, n2247, n2296, n2295, n2246, n2245;
    wire [71:0]d_out_11__N_1818_adj_2663;
    
    wire n9;
    wire [11:0]DataInReg_11__N_1855;
    
    wire n2724, n2243, n2242, n2241, n2240, n2239, n2238, n2237, 
        n2236, n2235, n2234, n9_adj_2616, n7, n2233, n2232, n2231, 
        n2230, n2229, n2228, n2227, n2226, n2225, n2224, n4, 
        n2223, n2222, n13061, n13818, n13817, n2221, n2220, n13815, 
        n2219, n2218, n2217, n2215, osc_clk_enable_1396, n2936, 
        n2935, n2934, n13812, n2933, n2932, n13811, n13810, n12896, 
        n2931, n2930, n2929, o_Rx_DV_c_0, n2928, n41, n14095, 
        osc_clk_enable_1458, n13753, n13806, n22, n6, n2897, n2896, 
        n2895, n2894, n2893, n2892, n2891, n2890, n2889, n2888, 
        n2887, n2886, n2885, n2884, n2883, n2881, n2277, n2276, 
        n2275, n2274, n2273, n2272, n2271, n2270, n2269, n2268, 
        n2267, n2266, n2265, n2264, n2263, n2262, n57, n2596, 
        n2595, n2594, n2591, n8980, n2586, n2581, n2580, n2579, 
        n2577, n2573, n2570, n2567, n2565, n2559, n2555, n8992, 
        n2552, n2551, n2550, n2548, n2723, n2722, n13816, n14101, 
        n2717, n2715, n2714, n2712, n2711, n2710, n2709, n2708, 
        n2707, n2704, n2702, n2701, n2700, n2699, n2698, n2696, 
        n13837, n2694, n2693, n2692, n2690, n2689, n2688, n2687, 
        n2683, n2682, n2681, n61, n62, n63, n64, n65, n66, 
        n67, n68, n70, n12946, n13805, n2880, n2879, n2882, 
        n2878, n8210, n2877, n2876, n2875, n2927, n2926, n2925, 
        n2924, n2261, n2260, n2259, n2258, n2257, n2256, n2255, 
        n2254, n2253, n2252, n2251, n2250, n2923, n2922, n2921, 
        n2920, n2919, n2918, n2917, n2916, n2915, n2914, n13803, 
        n2899, n2898, n13802, n13801, n2913, n13839, n12897, n13838, 
        n13836, n2912, n2911, n2910, n2909, n2908, n2907, n2906, 
        n2905, n2904, n2903, n2902, n2901, n2900, n13797, n8366, 
        n13796, osc_clk_enable_1457, n2731, n2732, n14098, n13792, 
        n2738, n2739, n13795, n2803, n13793, n13833, n13832, n13831, 
        n13791, n13788, n13785, n13824, n7695, n14097, n13823, 
        n13783, n9004, n13767, n8967, n13765, n12900, n12872, 
        n13151, n13763, n13776, n13775, n12219, n12218, n12217, 
        n12216, n12215, n12214, n12213, n14096, n12212, n12211, 
        n12210, n12209, n12208, n12207, n12206, n12205, n12204, 
        n12203, n12202, n12201, n12200, n12199, n12198, n12197, 
        n12196, n12195, n12194, n12193, n12192, n12191, n12190, 
        n13757, n12189, n14103, n14102, n14100, n14099, osc_clk_enable_1393, 
        n7986;
    
    VHI i2 (.Z(VCC_net));
    Mixer Mixer1 (.MixerOutCos({MixerOutCos}), .osc_clk(osc_clk), .MixerOutSin({MixerOutSin}), 
          .DiffOut_c(DiffOut_c), .RFIn_c(RFIn_c), .\LOCosine[2] (LOCosine[2]), 
          .\LOCosine[3] (LOCosine[3]), .\LOCosine[6] (LOCosine[6]), .\LOCosine[7] (LOCosine[7]), 
          .\LOCosine[8] (LOCosine[8]), .\LOCosine[9] (LOCosine[9]), .\LOCosine[10] (LOCosine[10]), 
          .\LOCosine[12] (LOCosine[12]), .GND_net(GND_net), .\LOCosine[11] (LOCosine[11]), 
          .\LOCosine[4] (LOCosine[4]), .\LOCosine[5] (LOCosine[5]), .\LOCosine[1] (LOCosine[1]), 
          .\LOSine[12] (LOSine[12]), .\LOSine[10] (LOSine[10]), .\LOSine[11] (LOSine[11]), 
          .\LOSine[8] (LOSine[8]), .\LOSine[9] (LOSine[9]), .\LOSine[6] (LOSine[6]), 
          .\LOSine[7] (LOSine[7]), .\LOSine[4] (LOSine[4]), .\LOSine[5] (LOSine[5]), 
          .\LOSine[2] (LOSine[2]), .\LOSine[3] (LOSine[3]), .\LOSine[1] (LOSine[1])) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(117[7] 125[2])
    LUT4 mux_378_i30_3_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(o_Rx_Byte_c_3), .D(n2579), .Z(n2710)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i30_3_lut_4_lut.init = 16'hfb0b;
    PUR PUR_INST (.PUR(VCC_net)) /* synthesis syn_instantiated=1 */ ;
    defparam PUR_INST.RST_PULSE = 1;
    FD1S3AX phase_inc_carrGen1_i0 (.D(phase_inc_carrGen[0]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[0]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i0.GSR = "ENABLED";
    PWM PWM1 (.osc_clk(osc_clk), .\DataInReg_11__N_1855[0] (DataInReg_11__N_1855[0]), 
        .PWMOut_c(PWMOut_c), .\DataInReg_11__N_1855[1] (DataInReg_11__N_1855[1]), 
        .\DataInReg_11__N_1855[2] (DataInReg_11__N_1855[2]), .\DataInReg_11__N_1855[3] (DataInReg_11__N_1855[3]), 
        .\DataInReg_11__N_1855[4] (DataInReg_11__N_1855[4]), .\DataInReg_11__N_1855[5] (DataInReg_11__N_1855[5]), 
        .\DataInReg_11__N_1855[6] (DataInReg_11__N_1855[6]), .\DataInReg_11__N_1855[7] (DataInReg_11__N_1855[7]), 
        .\DataInReg_11__N_1855[8] (DataInReg_11__N_1855[8]), .GND_net(GND_net), 
        .\DemodOut[9] (DemodOut[9])) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(146[5] 152[2])
    LUT4 mux_378_i12_4_lut (.A(o_Rx_Byte_c_0), .B(n2335), .C(o_Rx_Byte_c_3), 
         .D(o_Rx_Byte_c_2), .Z(n2728)) /* synthesis lut_function=(A (B (C (D)))+!A (B ((D)+!C)+!B !(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i12_4_lut.init = 16'hc505;
    LUT4 i2823_2_lut (.A(n932), .B(n7319), .Z(n2335)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i2823_2_lut.init = 16'hbbbb;
    FD1P3AX CICGain__i1 (.D(o_Rx_Byte_c_0), .SP(osc_clk_enable_1393), .CK(osc_clk), 
            .Q(CICGain[0]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam CICGain__i1.GSR = "ENABLED";
    LUT4 mux_378_i44_3_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(o_Rx_Byte_c_3), .D(n2565), .Z(n2696)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i44_3_lut_4_lut.init = 16'hfb0b;
    OB o_Rx_Byte_pad_6 (.I(o_Rx_Byte_c_6), .O(o_Rx_Byte[6]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(44[16:25])
    LUT4 mux_367_i8_4_lut (.A(n2732), .B(n999), .C(n2215), .D(n13757), 
         .Z(n2273)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i8_4_lut.init = 16'hc0ca;
    LUT4 mux_378_i28_3_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(o_Rx_Byte_c_3), .D(n2581), .Z(n2712)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i28_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_378_i23_3_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(o_Rx_Byte_c_3), .D(n2586), .Z(n2717)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i23_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_375_i8_3_lut (.A(n7319), .B(n936), .C(o_Rx_Byte_c_2), .Z(n2601)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_375_i8_3_lut.init = 16'hdada;
    LUT4 mux_378_i33_4_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(o_Rx_Byte_c_3), .D(n2314), .Z(n2707)) /* synthesis lut_function=(A (B ((D)+!C))+!A (B ((D)+!C)+!B !(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i33_4_lut_4_lut.init = 16'hcd0d;
    LUT4 mux_367_i9_4_lut (.A(n2731), .B(n998), .C(n2215), .D(n13757), 
         .Z(n2272)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i9_4_lut.init = 16'hcfca;
    LUT4 mux_378_i9_3_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), .C(o_Rx_Byte_c_3), 
         .D(n2600), .Z(n2731)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A ((D)+!C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i9_3_lut_4_lut.init = 16'hfd0d;
    LUT4 mux_375_i9_3_lut (.A(n7319), .B(n935), .C(o_Rx_Byte_c_2), .Z(n2600)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_375_i9_3_lut.init = 16'hdada;
    LUT4 mux_378_i42_3_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(o_Rx_Byte_c_3), .D(n2567), .Z(n2698)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i42_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_367_i5_4_lut (.A(n13791), .B(n1002), .C(n2215), .D(n13757), 
         .Z(n2276)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i5_4_lut.init = 16'hc0ca;
    LUT4 mux_378_i46_4_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(o_Rx_Byte_c_3), .D(n2301), .Z(n2694)) /* synthesis lut_function=(A ((C (D))+!B)+!A (B ((D)+!C)+!B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i46_4_lut_4_lut.init = 16'hf636;
    LUT4 mux_378_i8_3_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), .C(o_Rx_Byte_c_3), 
         .D(n2601), .Z(n2732)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i8_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_378_i36_3_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(o_Rx_Byte_c_3), .D(n2573), .Z(n2704)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i36_3_lut_4_lut.init = 16'hf606;
    OB o_Rx_Byte_pad_5 (.I(o_Rx_Byte_c_5), .O(o_Rx_Byte[5]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(44[16:25])
    LUT4 mux_378_i39_3_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(o_Rx_Byte_c_3), .D(n2570), .Z(n2701)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i39_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_378_i31_4_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(o_Rx_Byte_c_3), .D(n2316), .Z(n2709)) /* synthesis lut_function=(A ((C (D))+!B)+!A (B ((D)+!C)+!B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i31_4_lut_4_lut.init = 16'hf636;
    LUT4 mux_367_i10_4_lut (.A(n13797), .B(n997), .C(n2215), .D(n13757), 
         .Z(n2271)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i10_4_lut.init = 16'hc0ca;
    LUT4 mux_378_i48_4_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(o_Rx_Byte_c_3), .D(n2299), .Z(n2692)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (B ((D)+!C)+!B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i48_4_lut_4_lut.init = 16'hf434;
    LUT4 mux_367_i6_4_lut (.A(n13788), .B(n1001), .C(n2215), .D(n13757), 
         .Z(n2275)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i6_4_lut.init = 16'hc0ca;
    LUT4 i5907_3_lut (.A(n2215), .B(osc_clk_enable_1457), .C(n9004), .Z(osc_clk_enable_1396)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;
    defparam i5907_3_lut.init = 16'hc4c4;
    LUT4 mux_378_i22_4_lut_else_4_lut (.A(n922), .B(o_Rx_Byte_c_3), .C(o_Rx_Byte_c_2), 
         .D(n7319), .Z(n14098)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i22_4_lut_else_4_lut.init = 16'hbfff;
    OB o_Rx_Byte_pad_7 (.I(o_Rx_Byte_c_7), .O(o_Rx_Byte[7]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(44[16:25])
    OB o_Rx_DV_pad (.I(o_Rx_DV_c_0), .O(o_Rx_DV));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(43[13:20])
    OB o_Tx_Serial_pad (.I(o_Tx_Serial_c), .O(o_Tx_Serial));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(42[11:22])
    LUT4 mux_367_i53_4_lut (.A(n2687), .B(n954), .C(n2215), .D(n13757), 
         .Z(n2228)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i53_4_lut.init = 16'hc0ca;
    LUT4 i2745_4_lut (.A(o_Rx_Byte_c_2), .B(n13757), .C(n8967), .D(o_Rx_Byte_c_3), 
         .Z(n2803)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i2745_4_lut.init = 16'hfcee;
    \uart_tx(CLKS_PER_BIT=87)  uart_tx1 (.\UartClk[2] (UartClk_adj_2711[2]), 
            .o_Rx_Byte_c_0(o_Rx_Byte_c_0), .n12872(n12872), .n7319(n7319), 
            .o_Rx_Byte_c_4(o_Rx_Byte_c_4), .n2215(n2215), .o_Tx_Serial_c(o_Tx_Serial_c), 
            .o_Rx_DV_c_0(o_Rx_DV_c_0), .o_Rx_Byte_c_7(o_Rx_Byte_c_7), .o_Rx_Byte_c_2(o_Rx_Byte_c_2), 
            .osc_clk(osc_clk), .o_Rx_Byte_c_6(o_Rx_Byte_c_6), .o_Rx_Byte_c_5(o_Rx_Byte_c_5), 
            .o_Rx_Byte_c_3(o_Rx_Byte_c_3), .GND_net(GND_net), .n13765(n13765), 
            .n13753(n13753), .n13151(n13151)) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(184[32] 191[2])
    FD1S3AX phase_inc_carrGen1_i63 (.D(phase_inc_carrGen[63]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[63]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i63.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i62 (.D(phase_inc_carrGen[62]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[62]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i62.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i61 (.D(phase_inc_carrGen[61]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[61]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i61.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i60 (.D(phase_inc_carrGen[60]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[60]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i60.GSR = "ENABLED";
    LUT4 i2964_3_lut (.A(o_Rx_Byte_c_2), .B(n7319), .C(n941), .Z(n8967)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i2964_3_lut.init = 16'hc4c4;
    FD1S3AX phase_inc_carrGen1_i59 (.D(phase_inc_carrGen[59]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[59]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i59.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i58 (.D(phase_inc_carrGen[58]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[58]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i58.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i57 (.D(phase_inc_carrGen[57]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[57]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i57.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i56 (.D(phase_inc_carrGen[56]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[56]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i56.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i55 (.D(phase_inc_carrGen[55]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[55]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i55.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i54 (.D(phase_inc_carrGen[54]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[54]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i54.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i53 (.D(phase_inc_carrGen[53]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[53]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i53.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i52 (.D(phase_inc_carrGen[52]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[52]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i52.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i51 (.D(phase_inc_carrGen[51]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[51]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i51.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i50 (.D(phase_inc_carrGen[50]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[50]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i50.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i49 (.D(phase_inc_carrGen[49]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[49]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i49.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i48 (.D(phase_inc_carrGen[48]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[48]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i48.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i47 (.D(phase_inc_carrGen[47]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[47]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i47.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i46 (.D(phase_inc_carrGen[46]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[46]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i46.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i45 (.D(phase_inc_carrGen[45]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[45]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i45.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i44 (.D(phase_inc_carrGen[44]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[44]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i44.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i43 (.D(phase_inc_carrGen[43]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[43]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i43.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i42 (.D(phase_inc_carrGen[42]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[42]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i42.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i41 (.D(phase_inc_carrGen[41]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[41]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i41.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i40 (.D(phase_inc_carrGen[40]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[40]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i40.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i39 (.D(phase_inc_carrGen[39]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[39]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i39.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i38 (.D(phase_inc_carrGen[38]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[38]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i38.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i37 (.D(phase_inc_carrGen[37]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[37]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i37.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i36 (.D(phase_inc_carrGen[36]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[36]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i36.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i35 (.D(phase_inc_carrGen[35]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[35]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i35.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i34 (.D(phase_inc_carrGen[34]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[34]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i34.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i33 (.D(phase_inc_carrGen[33]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[33]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i33.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i32 (.D(phase_inc_carrGen[32]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[32]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i32.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i31 (.D(phase_inc_carrGen[31]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[31]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i31.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i30 (.D(phase_inc_carrGen[30]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[30]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i30.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i29 (.D(phase_inc_carrGen[29]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[29]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i29.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i28 (.D(phase_inc_carrGen[28]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[28]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i28.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i27 (.D(phase_inc_carrGen[27]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[27]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i27.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i26 (.D(phase_inc_carrGen[26]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[26]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i26.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i25 (.D(phase_inc_carrGen[25]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[25]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i25.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i24 (.D(phase_inc_carrGen[24]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[24]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i24.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i23 (.D(phase_inc_carrGen[23]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[23]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i23.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i22 (.D(phase_inc_carrGen[22]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[22]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i22.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i21 (.D(phase_inc_carrGen[21]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[21]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i21.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i20 (.D(phase_inc_carrGen[20]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[20]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i20.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i19 (.D(phase_inc_carrGen[19]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[19]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i19.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i18 (.D(phase_inc_carrGen[18]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[18]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i18.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i17 (.D(phase_inc_carrGen[17]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[17]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i17.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i16 (.D(phase_inc_carrGen[16]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[16]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i16.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i15 (.D(phase_inc_carrGen[15]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[15]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i15.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i14 (.D(phase_inc_carrGen[14]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[14]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i14.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i13 (.D(phase_inc_carrGen[13]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[13]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i13.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i12 (.D(phase_inc_carrGen[12]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[12]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i12.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i11 (.D(phase_inc_carrGen[11]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[11]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i11.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i10 (.D(phase_inc_carrGen[10]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[10]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i10.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i9 (.D(phase_inc_carrGen[9]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[9]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i9.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i8 (.D(phase_inc_carrGen[8]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[8]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i8.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i7 (.D(phase_inc_carrGen[7]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[7]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i7.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i6 (.D(phase_inc_carrGen[6]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[6]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i6.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i5 (.D(phase_inc_carrGen[5]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[5]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i5.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i4 (.D(phase_inc_carrGen[4]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[4]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i4.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i3 (.D(phase_inc_carrGen[3]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[3]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i3.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i2 (.D(phase_inc_carrGen[2]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[2]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i2.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i1 (.D(phase_inc_carrGen[1]), .CK(osc_clk), 
            .Q(phase_inc_carrGen1[1]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen1_i1.GSR = "ENABLED";
    OB o_Rx_Byte_pad_4 (.I(o_Rx_Byte_c_4), .O(o_Rx_Byte[4]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(44[16:25])
    OB o_Rx_Byte_pad_3 (.I(o_Rx_Byte_c_3), .O(o_Rx_Byte[3]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(44[16:25])
    OB o_Rx_Byte_pad_2 (.I(o_Rx_Byte_c_2), .O(o_Rx_Byte[2]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(44[16:25])
    OB o_Rx_Byte_pad_1 (.I(n7319), .O(o_Rx_Byte[1]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(44[16:25])
    OB o_Rx_Byte_pad_0 (.I(o_Rx_Byte_c_0), .O(o_Rx_Byte[0]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(44[16:25])
    OB MYLED_pad_7 (.I(GND_net), .O(MYLED[7]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(45[18:23])
    OB MYLED_pad_6 (.I(n7319), .O(MYLED[6]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(45[18:23])
    OB MYLED_pad_5 (.I(MYLED_c_5), .O(MYLED[5]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(45[18:23])
    OB MYLED_pad_4 (.I(MYLED_c_4), .O(MYLED[4]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(45[18:23])
    OB MYLED_pad_3 (.I(MYLED_c_3), .O(MYLED[3]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(45[18:23])
    OB MYLED_pad_2 (.I(MYLED_c_2), .O(MYLED[2]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(45[18:23])
    OB MYLED_pad_1 (.I(MYLED_c_1), .O(MYLED[1]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(45[18:23])
    OB MYLED_pad_0 (.I(MYLED_c_0), .O(MYLED[0]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(45[18:23])
    OB XOut_pad (.I(GND_net), .O(XOut));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(47[9:13])
    OB DiffOut_pad (.I(DiffOut_c), .O(DiffOut));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(49[9:16])
    OB PWMOut_pad (.I(PWMOut_c), .O(PWMOut));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(50[9:15])
    OB sinGen_pad (.I(sinGen_c), .O(sinGen));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(51[9:15])
    OB sin_out_pad (.I(GND_net), .O(sin_out));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(52[9:16])
    OB CIC_out_clkSin_pad (.I(GND_net), .O(CIC_out_clkSin));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(53[9:23])
    IB i_Rx_Serial_pad (.I(i_Rx_Serial), .O(i_Rx_Serial_c));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(40[13:24])
    IB XIn_pad (.I(XIn), .O(XIn_c));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(46[8:11])
    IB RFIn_pad (.I(RFIn), .O(RFIn_c));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(48[9:13])
    LUT4 mux_367_i4_4_lut (.A(n13785), .B(n1003), .C(n2215), .D(n13757), 
         .Z(n2277)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i4_4_lut.init = 16'hc0ca;
    LUT4 i5867_3_lut (.A(o_Rx_Byte_c_6), .B(n8210), .C(n41), .Z(osc_clk_enable_1457)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i5867_3_lut.init = 16'h2020;
    LUT4 i2800_4_lut (.A(n891), .B(o_Rx_Byte_c_3), .C(o_Rx_Byte_c_2), 
         .D(n7319), .Z(n2687)) /* synthesis lut_function=(A ((C)+!B)+!A !(B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i2800_4_lut.init = 16'hb3f3;
    LUT4 mux_378_i38_4_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(o_Rx_Byte_c_3), .D(n2309), .Z(n2702)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D))+!B !(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i38_4_lut_4_lut.init = 16'hcb0b;
    FD1P3AX CICGain__i2 (.D(n7319), .SP(osc_clk_enable_1393), .CK(osc_clk), 
            .Q(CICGain[1]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam CICGain__i2.GSR = "ENABLED";
    FD1P3JX phase_inc_carrGen_i0_i1 (.D(n2738), .SP(osc_clk_enable_1458), 
            .PD(n8366), .CK(osc_clk), .Q(phase_inc_carrGen[1]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i1.GSR = "ENABLED";
    LUT4 i5892_4_lut (.A(n22), .B(n8210), .C(o_Rx_Byte_c_4), .D(o_Rx_Byte_c_6), 
         .Z(n13061)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;
    defparam i5892_4_lut.init = 16'hfdff;
    LUT4 i33_4_lut (.A(o_Rx_Byte_c_3), .B(o_Rx_Byte_c_0), .C(o_Rx_Byte_c_2), 
         .D(n7319), .Z(n22)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A (B+((D)+!C)))) */ ;
    defparam i33_4_lut.init = 16'h2830;
    LUT4 mux_367_i7_4_lut (.A(n14097), .B(n1000), .C(n2215), .D(n13757), 
         .Z(n2274)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i7_4_lut.init = 16'hcfca;
    LUT4 mux_367_i54_4_lut (.A(n2555), .B(n953), .C(n2215), .D(n13753), 
         .Z(n2227)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i54_4_lut.init = 16'hcacf;
    LUT4 i2815_3_lut (.A(n890), .B(o_Rx_Byte_c_2), .C(n7319), .Z(n2555)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i2815_3_lut.init = 16'h8c8c;
    LUT4 mux_378_i34_4_lut_then_4_lut (.A(n910), .B(o_Rx_Byte_c_3), .C(o_Rx_Byte_c_2), 
         .D(n7319), .Z(n14102)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A !(B+(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i34_4_lut_then_4_lut.init = 16'h8303;
    LUT4 i5890_4_lut (.A(n12900), .B(n12896), .C(o_Rx_Byte_c_2), .D(n4), 
         .Z(n12897)) /* synthesis lut_function=(!(A (B)+!A !((C+!(D))+!B))) */ ;
    defparam i5890_4_lut.init = 16'h7377;
    LUT4 mux_378_i34_4_lut_else_4_lut (.A(n910), .B(o_Rx_Byte_c_3), .C(o_Rx_Byte_c_2), 
         .D(n7319), .Z(n14101)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A !(B+!(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i34_4_lut_else_4_lut.init = 16'hb030;
    LUT4 mux_367_i51_4_lut (.A(n2689), .B(n956), .C(n2215), .D(n13757), 
         .Z(n2230)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i51_4_lut.init = 16'hc0ca;
    LUT4 i2857_2_lut (.A(n893), .B(n7319), .Z(n2296)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i2857_2_lut.init = 16'h8888;
    LUT4 mux_367_i52_4_lut (.A(n2688), .B(n955), .C(n2215), .D(n13757), 
         .Z(n2229)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i52_4_lut.init = 16'hc0ca;
    LUT4 i2858_2_lut (.A(n892), .B(n7319), .Z(n2295)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i2858_2_lut.init = 16'hbbbb;
    LUT4 i5499_2_lut_3_lut (.A(o_Rx_Byte_c_3), .B(n13757), .C(n7319), 
         .Z(n12946)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i5499_2_lut_3_lut.init = 16'h2020;
    LUT4 mux_367_i49_4_lut (.A(n13839), .B(n958), .C(n2215), .D(n13757), 
         .Z(n2232)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i49_4_lut.init = 16'hcfca;
    LUT4 mux_378_i4_4_lut_else_4_lut (.A(o_Rx_Byte_c_2), .B(o_Rx_Byte_c_3), 
         .C(n7319), .D(o_Rx_Byte_c_0), .Z(n13783)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i4_4_lut_else_4_lut.init = 16'h6240;
    LUT4 mux_367_i50_4_lut (.A(n2690), .B(n957), .C(n2215), .D(n13757), 
         .Z(n2231)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i50_4_lut.init = 16'hc0ca;
    LUT4 mux_378_i50_3_lut (.A(o_Rx_Byte_c_0), .B(n2559), .C(o_Rx_Byte_c_3), 
         .Z(n2690)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i50_3_lut.init = 16'hc5c5;
    LUT4 mux_375_i50_3_lut (.A(n7319), .B(n894), .C(o_Rx_Byte_c_2), .Z(n2559)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_375_i50_3_lut.init = 16'hdada;
    LUT4 mux_367_i47_4_lut (.A(n2693), .B(n960), .C(n2215), .D(n13757), 
         .Z(n2234)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i47_4_lut.init = 16'hcfca;
    LUT4 mux_378_i47_4_lut (.A(o_Rx_Byte_c_2), .B(n897), .C(o_Rx_Byte_c_3), 
         .D(n7319), .Z(n2693)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A !(C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i47_4_lut.init = 16'h85a5;
    LUT4 mux_367_i48_4_lut (.A(n2692), .B(n959), .C(n2215), .D(n13757), 
         .Z(n2233)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i48_4_lut.init = 16'hc0ca;
    LUT4 i2854_2_lut (.A(n896), .B(n7319), .Z(n2299)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i2854_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_then_4_lut (.A(o_Rx_Byte_c_3), .B(o_Rx_Byte_c_0), .C(o_Rx_Byte_c_4), 
         .D(o_Rx_Byte_c_2), .Z(n13793)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C+!(D)))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(207[4] 232[10])
    defparam i1_4_lut_then_4_lut.init = 16'h021d;
    LUT4 i1_4_lut_else_4_lut (.A(o_Rx_Byte_c_3), .B(o_Rx_Byte_c_0), .C(o_Rx_Byte_c_4), 
         .D(o_Rx_Byte_c_2), .Z(n13792)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A (B (C)+!B !(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(207[4] 232[10])
    defparam i1_4_lut_else_4_lut.init = 16'h1f06;
    LUT4 mux_367_i45_4_lut (.A(n13836), .B(n962), .C(n2215), .D(n13757), 
         .Z(n2236)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i45_4_lut.init = 16'hc0ca;
    CCU2D add_702_63 (.A0(GND_net), .B0(n9004), .C0(n2218), .D0(phase_inc_carrGen[62]), 
          .A1(GND_net), .B1(n9004), .C1(n2217), .D1(phase_inc_carrGen[63]), 
          .CIN(n12219), .S0(n2876), .S1(n2875));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_63.INIT0 = 16'h569a;
    defparam add_702_63.INIT1 = 16'h569a;
    defparam add_702_63.INJECT1_0 = "NO";
    defparam add_702_63.INJECT1_1 = "NO";
    CCU2D add_702_61 (.A0(GND_net), .B0(n9004), .C0(n2220), .D0(phase_inc_carrGen[60]), 
          .A1(GND_net), .B1(n9004), .C1(n2219), .D1(phase_inc_carrGen[61]), 
          .CIN(n12218), .COUT(n12219), .S0(n2878), .S1(n2877));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_61.INIT0 = 16'h569a;
    defparam add_702_61.INIT1 = 16'h569a;
    defparam add_702_61.INJECT1_0 = "NO";
    defparam add_702_61.INJECT1_1 = "NO";
    LUT4 mux_378_i10_4_lut_then_4_lut (.A(o_Rx_Byte_c_2), .B(o_Rx_Byte_c_3), 
         .C(n7319), .D(o_Rx_Byte_c_0), .Z(n13796)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A (B (C)+!B (D))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i10_4_lut_then_4_lut.init = 16'hd1e2;
    CCU2D add_702_59 (.A0(GND_net), .B0(n9004), .C0(n2222), .D0(phase_inc_carrGen[58]), 
          .A1(GND_net), .B1(n9004), .C1(n2221), .D1(phase_inc_carrGen[59]), 
          .CIN(n12217), .COUT(n12218), .S0(n2880), .S1(n2879));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_59.INIT0 = 16'h569a;
    defparam add_702_59.INIT1 = 16'h569a;
    defparam add_702_59.INJECT1_0 = "NO";
    defparam add_702_59.INJECT1_1 = "NO";
    CCU2D add_702_57 (.A0(GND_net), .B0(n9004), .C0(n2224), .D0(phase_inc_carrGen[56]), 
          .A1(GND_net), .B1(n9004), .C1(n2223), .D1(phase_inc_carrGen[57]), 
          .CIN(n12216), .COUT(n12217), .S0(n2882), .S1(n2881));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_57.INIT0 = 16'h569a;
    defparam add_702_57.INIT1 = 16'h569a;
    defparam add_702_57.INJECT1_0 = "NO";
    defparam add_702_57.INJECT1_1 = "NO";
    CCU2D add_702_55 (.A0(GND_net), .B0(n9004), .C0(n2226), .D0(phase_inc_carrGen[54]), 
          .A1(GND_net), .B1(n9004), .C1(n2225), .D1(phase_inc_carrGen[55]), 
          .CIN(n12215), .COUT(n12216), .S0(n2884), .S1(n2883));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_55.INIT0 = 16'h569a;
    defparam add_702_55.INIT1 = 16'h569a;
    defparam add_702_55.INJECT1_0 = "NO";
    defparam add_702_55.INJECT1_1 = "NO";
    LUT4 mux_378_i10_4_lut_else_4_lut (.A(o_Rx_Byte_c_2), .B(o_Rx_Byte_c_3), 
         .C(n7319), .D(o_Rx_Byte_c_0), .Z(n13795)) /* synthesis lut_function=(!(A (B+(D))+!A !(B (C)+!B (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i10_4_lut_else_4_lut.init = 16'h5162;
    LUT4 mux_378_i58_3_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(o_Rx_Byte_c_3), .D(n2551), .Z(n2682)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i58_3_lut_4_lut.init = 16'hf202;
    CCU2D add_702_53 (.A0(GND_net), .B0(n9004), .C0(n2228), .D0(phase_inc_carrGen[52]), 
          .A1(GND_net), .B1(n9004), .C1(n2227), .D1(phase_inc_carrGen[53]), 
          .CIN(n12214), .COUT(n12215), .S0(n2886), .S1(n2885));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_53.INIT0 = 16'h569a;
    defparam add_702_53.INIT1 = 16'h569a;
    defparam add_702_53.INJECT1_0 = "NO";
    defparam add_702_53.INJECT1_1 = "NO";
    LUT4 mux_367_i46_4_lut (.A(n2694), .B(n961), .C(n2215), .D(n13757), 
         .Z(n2235)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i46_4_lut.init = 16'hc0ca;
    LUT4 mux_378_i32_3_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(o_Rx_Byte_c_3), .D(n2577), .Z(n2708)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i32_3_lut_4_lut.init = 16'hf202;
    LUT4 i2852_2_lut (.A(n898), .B(n7319), .Z(n2301)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i2852_2_lut.init = 16'h8888;
    CCU2D add_702_51 (.A0(o_Rx_Byte_c_4), .B0(n9004), .C0(n2230), .D0(phase_inc_carrGen[50]), 
          .A1(GND_net), .B1(n9004), .C1(n2229), .D1(phase_inc_carrGen[51]), 
          .CIN(n12213), .COUT(n12214), .S0(n2888), .S1(n2887));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_51.INIT0 = 16'hb874;
    defparam add_702_51.INIT1 = 16'h569a;
    defparam add_702_51.INJECT1_0 = "NO";
    defparam add_702_51.INJECT1_1 = "NO";
    CCU2D add_702_49 (.A0(o_Rx_Byte_c_4), .B0(n9004), .C0(n2232), .D0(phase_inc_carrGen[48]), 
          .A1(o_Rx_Byte_c_4), .B1(n9004), .C1(n2231), .D1(phase_inc_carrGen[49]), 
          .CIN(n12212), .COUT(n12213), .S0(n2890), .S1(n2889));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_49.INIT0 = 16'hb874;
    defparam add_702_49.INIT1 = 16'hb874;
    defparam add_702_49.INJECT1_0 = "NO";
    defparam add_702_49.INJECT1_1 = "NO";
    CCU2D add_702_47 (.A0(o_Rx_Byte_c_4), .B0(n9004), .C0(n2234), .D0(phase_inc_carrGen[46]), 
          .A1(GND_net), .B1(n9004), .C1(n2233), .D1(phase_inc_carrGen[47]), 
          .CIN(n12211), .COUT(n12212), .S0(n2892), .S1(n2891));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_47.INIT0 = 16'hb874;
    defparam add_702_47.INIT1 = 16'h569a;
    defparam add_702_47.INJECT1_0 = "NO";
    defparam add_702_47.INJECT1_1 = "NO";
    CCU2D add_702_45 (.A0(n9004), .B0(n9004), .C0(n2236), .D0(phase_inc_carrGen[44]), 
          .A1(GND_net), .B1(n9004), .C1(n2235), .D1(phase_inc_carrGen[45]), 
          .CIN(n12210), .COUT(n12211), .S0(n2894), .S1(n2893));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_45.INIT0 = 16'h569a;
    defparam add_702_45.INIT1 = 16'h569a;
    defparam add_702_45.INJECT1_0 = "NO";
    defparam add_702_45.INJECT1_1 = "NO";
    LUT4 mux_378_i57_3_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(o_Rx_Byte_c_3), .D(n2552), .Z(n2683)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i57_3_lut_4_lut.init = 16'hf101;
    LUT4 mux_378_i11_4_lut_then_4_lut (.A(n933), .B(o_Rx_Byte_c_3), .C(o_Rx_Byte_c_2), 
         .D(n7319), .Z(n13802)) /* synthesis lut_function=(A (B)+!A !((C (D))+!B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i11_4_lut_then_4_lut.init = 16'h8ccc;
    LUT4 mux_378_i11_4_lut_else_4_lut (.A(n933), .B(o_Rx_Byte_c_3), .C(o_Rx_Byte_c_2), 
         .D(n7319), .Z(n13801)) /* synthesis lut_function=(A (B+!(C))+!A !(B (C (D))+!B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i11_4_lut_else_4_lut.init = 16'h8fcf;
    LUT4 mux_378_i51_4_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(o_Rx_Byte_c_3), .D(n2296), .Z(n2689)) /* synthesis lut_function=(A (((D)+!C)+!B)+!A (B ((D)+!C)+!B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i51_4_lut_4_lut.init = 16'hfe3e;
    LUT4 i1_4_lut_then_4_lut_adj_60 (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(o_Rx_Byte_c_4), .D(o_Rx_Byte_c_3), .Z(n13805)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B (D)))) */ ;
    defparam i1_4_lut_then_4_lut_adj_60.init = 16'h0411;
    LUT4 mux_378_i18_3_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(o_Rx_Byte_c_3), .D(n2591), .Z(n2722)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i18_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i1_4_lut_else_4_lut_adj_61 (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_4), 
         .C(o_Rx_Byte_c_3), .Z(n13804)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_4_lut_else_4_lut_adj_61.init = 16'h1010;
    LUT4 mux_367_i43_4_lut (.A(n13833), .B(n964), .C(n2215), .D(n13757), 
         .Z(n2238)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i43_4_lut.init = 16'hcfca;
    LUT4 mux_378_i15_3_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(o_Rx_Byte_c_3), .D(n2594), .Z(n2725)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i15_3_lut_4_lut.init = 16'hf101;
    LUT4 i1_4_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), .C(o_Rx_Byte_c_3), 
         .D(n13765), .Z(n12900)) /* synthesis lut_function=(!(A (C+(D))+!A (B+((D)+!C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i1_4_lut_4_lut.init = 16'h001a;
    LUT4 mux_367_i44_4_lut (.A(n2696), .B(n963), .C(n2215), .D(n13757), 
         .Z(n2237)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i44_4_lut.init = 16'hc0ca;
    LUT4 mux_375_i44_3_lut (.A(n7319), .B(n900), .C(o_Rx_Byte_c_2), .Z(n2565)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_375_i44_3_lut.init = 16'hdada;
    LUT4 mux_378_i7_4_lut_then_4_lut (.A(n937), .B(o_Rx_Byte_c_3), .C(o_Rx_Byte_c_2), 
         .D(n7319), .Z(n14096)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A !(B+(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i7_4_lut_then_4_lut.init = 16'h8303;
    LUT4 mux_378_i59_3_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(o_Rx_Byte_c_3), .D(n2550), .Z(n2681)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i59_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_378_i52_4_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(o_Rx_Byte_c_3), .D(n2295), .Z(n2688)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B ((D)+!C)+!B !(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i52_4_lut_4_lut.init = 16'hc707;
    LUT4 i1_4_lut (.A(n7319), .B(o_Rx_Byte_c_3), .C(o_Rx_Byte_c_4), .D(o_Rx_Byte_c_0), 
         .Z(n4)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+(C+!(D))))) */ ;
    defparam i1_4_lut.init = 16'h0322;
    LUT4 mux_378_i20_4_lut_then_4_lut (.A(o_Rx_Byte_c_2), .B(o_Rx_Byte_c_3), 
         .C(n7319), .D(o_Rx_Byte_c_0), .Z(n13811)) /* synthesis lut_function=(A (B+!(D))+!A !(B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i20_4_lut_then_4_lut.init = 16'h9dbf;
    LUT4 mux_378_i29_3_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(o_Rx_Byte_c_3), .D(n2580), .Z(n2711)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i29_3_lut_4_lut.init = 16'hf707;
    SinCos SinCos1 (.osc_clk(osc_clk), .VCC_net(VCC_net), .GND_net(GND_net), 
           .\phase_accum[57] (phase_accum[57]), .\phase_accum[58] (phase_accum[58]), 
           .\phase_accum[59] (phase_accum[59]), .\phase_accum[60] (phase_accum[60]), 
           .\phase_accum[61] (phase_accum[61]), .\phase_accum[62] (phase_accum[62]), 
           .\phase_accum[63] (phase_accum[63]), .\LOSine[1] (LOSine[1]), 
           .\LOSine[2] (LOSine[2]), .\LOSine[3] (LOSine[3]), .\LOSine[4] (LOSine[4]), 
           .\LOSine[5] (LOSine[5]), .\LOSine[6] (LOSine[6]), .\LOSine[7] (LOSine[7]), 
           .\LOSine[8] (LOSine[8]), .\LOSine[9] (LOSine[9]), .\LOSine[10] (LOSine[10]), 
           .\LOSine[11] (LOSine[11]), .\LOSine[12] (LOSine[12]), .\LOCosine[1] (LOCosine[1]), 
           .\LOCosine[2] (LOCosine[2]), .\LOCosine[3] (LOCosine[3]), .\LOCosine[4] (LOCosine[4]), 
           .\LOCosine[5] (LOCosine[5]), .\LOCosine[6] (LOCosine[6]), .\LOCosine[7] (LOCosine[7]), 
           .\LOCosine[8] (LOCosine[8]), .\LOCosine[9] (LOCosine[9]), .\LOCosine[10] (LOCosine[10]), 
           .\LOCosine[11] (LOCosine[11]), .\LOCosine[12] (LOCosine[12]), 
           .\phase_accum[56] (phase_accum[56])) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    CCU2D add_702_43 (.A0(n9004), .B0(n9004), .C0(n2238), .D0(phase_inc_carrGen[42]), 
          .A1(o_Rx_Byte_c_4), .B1(n9004), .C1(n2237), .D1(phase_inc_carrGen[43]), 
          .CIN(n12209), .COUT(n12210), .S0(n2896), .S1(n2895));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_43.INIT0 = 16'h569a;
    defparam add_702_43.INIT1 = 16'hb874;
    defparam add_702_43.INJECT1_0 = "NO";
    defparam add_702_43.INJECT1_1 = "NO";
    CCU2D add_702_41 (.A0(o_Rx_Byte_c_4), .B0(n9004), .C0(n2240), .D0(phase_inc_carrGen[40]), 
          .A1(o_Rx_Byte_c_4), .B1(n9004), .C1(n2239), .D1(phase_inc_carrGen[41]), 
          .CIN(n12208), .COUT(n12209), .S0(n2898), .S1(n2897));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_41.INIT0 = 16'hb874;
    defparam add_702_41.INIT1 = 16'hb874;
    defparam add_702_41.INJECT1_0 = "NO";
    defparam add_702_41.INJECT1_1 = "NO";
    CCU2D add_702_39 (.A0(n9004), .B0(n9004), .C0(n2242), .D0(phase_inc_carrGen[38]), 
          .A1(o_Rx_Byte_c_4), .B1(n9004), .C1(n2241), .D1(phase_inc_carrGen[39]), 
          .CIN(n12207), .COUT(n12208), .S0(n2900), .S1(n2899));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_39.INIT0 = 16'h569a;
    defparam add_702_39.INIT1 = 16'h74b8;
    defparam add_702_39.INJECT1_0 = "NO";
    defparam add_702_39.INJECT1_1 = "NO";
    CCU2D add_702_37 (.A0(o_Rx_Byte_c_4), .B0(n9004), .C0(n2244), .D0(phase_inc_carrGen[36]), 
          .A1(n9004), .B1(n9004), .C1(n2243), .D1(phase_inc_carrGen[37]), 
          .CIN(n12206), .COUT(n12207), .S0(n2902), .S1(n2901));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_37.INIT0 = 16'h74b8;
    defparam add_702_37.INIT1 = 16'h569a;
    defparam add_702_37.INJECT1_0 = "NO";
    defparam add_702_37.INJECT1_1 = "NO";
    CCU2D add_702_35 (.A0(o_Rx_Byte_c_4), .B0(n9004), .C0(n2246), .D0(phase_inc_carrGen[34]), 
          .A1(n9004), .B1(n9004), .C1(n2245), .D1(phase_inc_carrGen[35]), 
          .CIN(n12205), .COUT(n12206), .S0(n2904), .S1(n2903));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_35.INIT0 = 16'hb874;
    defparam add_702_35.INIT1 = 16'h569a;
    defparam add_702_35.INJECT1_0 = "NO";
    defparam add_702_35.INJECT1_1 = "NO";
    CCU2D add_702_33 (.A0(o_Rx_Byte_c_4), .B0(n9004), .C0(n2248), .D0(phase_inc_carrGen[32]), 
          .A1(o_Rx_Byte_c_4), .B1(n9004), .C1(n2247), .D1(phase_inc_carrGen[33]), 
          .CIN(n12204), .COUT(n12205), .S0(n2906), .S1(n2905));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_33.INIT0 = 16'hb874;
    defparam add_702_33.INIT1 = 16'hb874;
    defparam add_702_33.INJECT1_0 = "NO";
    defparam add_702_33.INJECT1_1 = "NO";
    CCU2D add_702_31 (.A0(o_Rx_Byte_c_4), .B0(n9004), .C0(n2250), .D0(phase_inc_carrGen[30]), 
          .A1(n9004), .B1(n9004), .C1(n2249), .D1(phase_inc_carrGen[31]), 
          .CIN(n12203), .COUT(n12204), .S0(n2908), .S1(n2907));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_31.INIT0 = 16'hb874;
    defparam add_702_31.INIT1 = 16'h569a;
    defparam add_702_31.INJECT1_0 = "NO";
    defparam add_702_31.INJECT1_1 = "NO";
    CCU2D add_702_29 (.A0(n9004), .B0(n9004), .C0(n2252), .D0(phase_inc_carrGen[28]), 
          .A1(o_Rx_Byte_c_4), .B1(n9004), .C1(n2251), .D1(phase_inc_carrGen[29]), 
          .CIN(n12202), .COUT(n12203), .S0(n2910), .S1(n2909));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_29.INIT0 = 16'h569a;
    defparam add_702_29.INIT1 = 16'h74b8;
    defparam add_702_29.INJECT1_0 = "NO";
    defparam add_702_29.INJECT1_1 = "NO";
    CCU2D add_702_27 (.A0(o_Rx_Byte_c_4), .B0(n9004), .C0(n2254), .D0(phase_inc_carrGen[26]), 
          .A1(GND_net), .B1(n9004), .C1(n2253), .D1(phase_inc_carrGen[27]), 
          .CIN(n12201), .COUT(n12202), .S0(n2912), .S1(n2911));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_27.INIT0 = 16'h74b8;
    defparam add_702_27.INIT1 = 16'h569a;
    defparam add_702_27.INJECT1_0 = "NO";
    defparam add_702_27.INJECT1_1 = "NO";
    CCU2D add_702_25 (.A0(o_Rx_Byte_c_4), .B0(n9004), .C0(n2256), .D0(phase_inc_carrGen[24]), 
          .A1(o_Rx_Byte_c_4), .B1(n9004), .C1(n2255), .D1(phase_inc_carrGen[25]), 
          .CIN(n12200), .COUT(n12201), .S0(n2914), .S1(n2913));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_25.INIT0 = 16'h74b8;
    defparam add_702_25.INIT1 = 16'hb874;
    defparam add_702_25.INJECT1_0 = "NO";
    defparam add_702_25.INJECT1_1 = "NO";
    CCU2D add_702_23 (.A0(GND_net), .B0(n9004), .C0(n2258), .D0(phase_inc_carrGen[22]), 
          .A1(o_Rx_Byte_c_4), .B1(n9004), .C1(n2257), .D1(phase_inc_carrGen[23]), 
          .CIN(n12199), .COUT(n12200), .S0(n2916), .S1(n2915));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_23.INIT0 = 16'h569a;
    defparam add_702_23.INIT1 = 16'h74b8;
    defparam add_702_23.INJECT1_0 = "NO";
    defparam add_702_23.INJECT1_1 = "NO";
    CCU2D add_702_21 (.A0(o_Rx_Byte_c_4), .B0(n9004), .C0(n2260), .D0(phase_inc_carrGen[20]), 
          .A1(GND_net), .B1(n9004), .C1(n2259), .D1(phase_inc_carrGen[21]), 
          .CIN(n12198), .COUT(n12199), .S0(n2918), .S1(n2917));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_21.INIT0 = 16'hb874;
    defparam add_702_21.INIT1 = 16'h569a;
    defparam add_702_21.INJECT1_0 = "NO";
    defparam add_702_21.INJECT1_1 = "NO";
    CCU2D add_702_19 (.A0(o_Rx_Byte_c_4), .B0(n9004), .C0(n2262), .D0(phase_inc_carrGen[18]), 
          .A1(n9004), .B1(n9004), .C1(n2261), .D1(phase_inc_carrGen[19]), 
          .CIN(n12197), .COUT(n12198), .S0(n2920), .S1(n2919));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_19.INIT0 = 16'hb874;
    defparam add_702_19.INIT1 = 16'h569a;
    defparam add_702_19.INJECT1_0 = "NO";
    defparam add_702_19.INJECT1_1 = "NO";
    CCU2D add_702_17 (.A0(o_Rx_Byte_c_4), .B0(n9004), .C0(n2264), .D0(phase_inc_carrGen[16]), 
          .A1(o_Rx_Byte_c_4), .B1(n9004), .C1(n2263), .D1(phase_inc_carrGen[17]), 
          .CIN(n12196), .COUT(n12197), .S0(n2922), .S1(n2921));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_17.INIT0 = 16'hb874;
    defparam add_702_17.INIT1 = 16'hb874;
    defparam add_702_17.INJECT1_0 = "NO";
    defparam add_702_17.INJECT1_1 = "NO";
    CCU2D add_702_15 (.A0(n9004), .B0(n9004), .C0(n2266), .D0(phase_inc_carrGen[14]), 
          .A1(n9004), .B1(n9004), .C1(n2265), .D1(phase_inc_carrGen[15]), 
          .CIN(n12195), .COUT(n12196), .S0(n2924), .S1(n2923));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_15.INIT0 = 16'h569a;
    defparam add_702_15.INIT1 = 16'h569a;
    defparam add_702_15.INJECT1_0 = "NO";
    defparam add_702_15.INJECT1_1 = "NO";
    CCU2D add_702_13 (.A0(o_Rx_Byte_c_4), .B0(n9004), .C0(n2268), .D0(phase_inc_carrGen[12]), 
          .A1(n9004), .B1(n9004), .C1(n2267), .D1(phase_inc_carrGen[13]), 
          .CIN(n12194), .COUT(n12195), .S0(n2926), .S1(n2925));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_13.INIT0 = 16'hb874;
    defparam add_702_13.INIT1 = 16'h569a;
    defparam add_702_13.INJECT1_0 = "NO";
    defparam add_702_13.INJECT1_1 = "NO";
    CCU2D add_702_11 (.A0(GND_net), .B0(n9004), .C0(n2270), .D0(phase_inc_carrGen[10]), 
          .A1(GND_net), .B1(n9004), .C1(n2269), .D1(phase_inc_carrGen[11]), 
          .CIN(n12193), .COUT(n12194), .S0(n2928), .S1(n2927));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_11.INIT0 = 16'h569a;
    defparam add_702_11.INIT1 = 16'h569a;
    defparam add_702_11.INJECT1_0 = "NO";
    defparam add_702_11.INJECT1_1 = "NO";
    CCU2D add_702_9 (.A0(o_Rx_Byte_c_4), .B0(n9004), .C0(n2272), .D0(phase_inc_carrGen[8]), 
          .A1(n9004), .B1(n9004), .C1(n2271), .D1(phase_inc_carrGen[9]), 
          .CIN(n12192), .COUT(n12193), .S0(n2930), .S1(n2929));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_9.INIT0 = 16'h74b8;
    defparam add_702_9.INIT1 = 16'h569a;
    defparam add_702_9.INJECT1_0 = "NO";
    defparam add_702_9.INJECT1_1 = "NO";
    CCU2D add_702_7 (.A0(n9004), .B0(n9004), .C0(n2274), .D0(phase_inc_carrGen[6]), 
          .A1(o_Rx_Byte_c_4), .B1(n9004), .C1(n2273), .D1(phase_inc_carrGen[7]), 
          .CIN(n12191), .COUT(n12192), .S0(n2932), .S1(n2931));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_7.INIT0 = 16'h569a;
    defparam add_702_7.INIT1 = 16'hb874;
    defparam add_702_7.INJECT1_0 = "NO";
    defparam add_702_7.INJECT1_1 = "NO";
    CCU2D add_702_5 (.A0(GND_net), .B0(n9004), .C0(n2276), .D0(phase_inc_carrGen[4]), 
          .A1(n9004), .B1(n9004), .C1(n2275), .D1(phase_inc_carrGen[5]), 
          .CIN(n12190), .COUT(n12191), .S0(n2934), .S1(n2933));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_5.INIT0 = 16'h569a;
    defparam add_702_5.INIT1 = 16'h569a;
    defparam add_702_5.INJECT1_0 = "NO";
    defparam add_702_5.INJECT1_1 = "NO";
    CCU2D add_702_3 (.A0(o_Rx_Byte_c_4), .B0(n9004), .C0(n2803), .D0(phase_inc_carrGen[2]), 
          .A1(o_Rx_Byte_c_4), .B1(n9004), .C1(n2277), .D1(phase_inc_carrGen[3]), 
          .CIN(n12189), .COUT(n12190), .S0(n2936), .S1(n2935));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_3.INIT0 = 16'hb874;
    defparam add_702_3.INIT1 = 16'h74b8;
    defparam add_702_3.INJECT1_0 = "NO";
    defparam add_702_3.INJECT1_1 = "NO";
    CCU2D add_702_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n13061), .B1(n12897), .C1(GND_net), .D1(GND_net), .COUT(n12189));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam add_702_1.INIT0 = 16'hF000;
    defparam add_702_1.INIT1 = 16'hffff;
    defparam add_702_1.INJECT1_0 = "NO";
    defparam add_702_1.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_63 (.A0(phase_inc_carrGen[63]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11611), .S0(n880));
    defparam sub_37_add_2_63.INIT0 = 16'h5555;
    defparam sub_37_add_2_63.INIT1 = 16'h0000;
    defparam sub_37_add_2_63.INJECT1_0 = "NO";
    defparam sub_37_add_2_63.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_61 (.A0(phase_inc_carrGen[61]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[62]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11610), .COUT(n11611), .S0(n882), .S1(n881));
    defparam sub_37_add_2_61.INIT0 = 16'h5555;
    defparam sub_37_add_2_61.INIT1 = 16'h5555;
    defparam sub_37_add_2_61.INJECT1_0 = "NO";
    defparam sub_37_add_2_61.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_59 (.A0(phase_inc_carrGen[59]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[60]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11609), .COUT(n11610), .S0(n884), .S1(n883));
    defparam sub_37_add_2_59.INIT0 = 16'h5555;
    defparam sub_37_add_2_59.INIT1 = 16'h5555;
    defparam sub_37_add_2_59.INJECT1_0 = "NO";
    defparam sub_37_add_2_59.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_57 (.A0(phase_inc_carrGen[57]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[58]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11608), .COUT(n11609), .S0(n886), .S1(n885));
    defparam sub_37_add_2_57.INIT0 = 16'h5555;
    defparam sub_37_add_2_57.INIT1 = 16'h5555;
    defparam sub_37_add_2_57.INJECT1_0 = "NO";
    defparam sub_37_add_2_57.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_55 (.A0(phase_inc_carrGen[55]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[56]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11607), .COUT(n11608), .S0(n888), .S1(n887));
    defparam sub_37_add_2_55.INIT0 = 16'h5555;
    defparam sub_37_add_2_55.INIT1 = 16'h5555;
    defparam sub_37_add_2_55.INJECT1_0 = "NO";
    defparam sub_37_add_2_55.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_53 (.A0(phase_inc_carrGen[53]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[54]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11606), .COUT(n11607), .S0(n890), .S1(n889));
    defparam sub_37_add_2_53.INIT0 = 16'h5555;
    defparam sub_37_add_2_53.INIT1 = 16'h5555;
    defparam sub_37_add_2_53.INJECT1_0 = "NO";
    defparam sub_37_add_2_53.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_51 (.A0(phase_inc_carrGen[51]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[52]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11605), .COUT(n11606), .S0(n892), .S1(n891));
    defparam sub_37_add_2_51.INIT0 = 16'h5555;
    defparam sub_37_add_2_51.INIT1 = 16'h5555;
    defparam sub_37_add_2_51.INJECT1_0 = "NO";
    defparam sub_37_add_2_51.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_49 (.A0(phase_inc_carrGen[49]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[50]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11604), .COUT(n11605), .S0(n894), .S1(n893));
    defparam sub_37_add_2_49.INIT0 = 16'h5aaa;
    defparam sub_37_add_2_49.INIT1 = 16'h5aaa;
    defparam sub_37_add_2_49.INJECT1_0 = "NO";
    defparam sub_37_add_2_49.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_47 (.A0(phase_inc_carrGen[47]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[48]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11603), .COUT(n11604), .S0(n896), .S1(n895));
    defparam sub_37_add_2_47.INIT0 = 16'h5555;
    defparam sub_37_add_2_47.INIT1 = 16'h5aaa;
    defparam sub_37_add_2_47.INJECT1_0 = "NO";
    defparam sub_37_add_2_47.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_45 (.A0(phase_inc_carrGen[45]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[46]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11602), .COUT(n11603), .S0(n898), .S1(n897));
    defparam sub_37_add_2_45.INIT0 = 16'h5555;
    defparam sub_37_add_2_45.INIT1 = 16'h5aaa;
    defparam sub_37_add_2_45.INJECT1_0 = "NO";
    defparam sub_37_add_2_45.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_43 (.A0(phase_inc_carrGen[43]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[44]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11601), .COUT(n11602), .S0(n900), .S1(n899));
    defparam sub_37_add_2_43.INIT0 = 16'h5aaa;
    defparam sub_37_add_2_43.INIT1 = 16'h5aaa;
    defparam sub_37_add_2_43.INJECT1_0 = "NO";
    defparam sub_37_add_2_43.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_41 (.A0(phase_inc_carrGen[41]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[42]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11600), .COUT(n11601), .S0(n902), .S1(n901));
    defparam sub_37_add_2_41.INIT0 = 16'h5aaa;
    defparam sub_37_add_2_41.INIT1 = 16'h5aaa;
    defparam sub_37_add_2_41.INJECT1_0 = "NO";
    defparam sub_37_add_2_41.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_39 (.A0(phase_inc_carrGen[39]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[40]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11599), .COUT(n11600), .S0(n904), .S1(n903));
    defparam sub_37_add_2_39.INIT0 = 16'h5555;
    defparam sub_37_add_2_39.INIT1 = 16'h5aaa;
    defparam sub_37_add_2_39.INJECT1_0 = "NO";
    defparam sub_37_add_2_39.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_37 (.A0(phase_inc_carrGen[37]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[38]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11598), .COUT(n11599), .S0(n906), .S1(n905));
    defparam sub_37_add_2_37.INIT0 = 16'h5aaa;
    defparam sub_37_add_2_37.INIT1 = 16'h5aaa;
    defparam sub_37_add_2_37.INJECT1_0 = "NO";
    defparam sub_37_add_2_37.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_35 (.A0(phase_inc_carrGen[35]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[36]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11597), .COUT(n11598), .S0(n908), .S1(n907));
    defparam sub_37_add_2_35.INIT0 = 16'h5aaa;
    defparam sub_37_add_2_35.INIT1 = 16'h5555;
    defparam sub_37_add_2_35.INJECT1_0 = "NO";
    defparam sub_37_add_2_35.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_33 (.A0(phase_inc_carrGen[33]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[34]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11596), .COUT(n11597), .S0(n910), .S1(n909));
    defparam sub_37_add_2_33.INIT0 = 16'h5aaa;
    defparam sub_37_add_2_33.INIT1 = 16'h5aaa;
    defparam sub_37_add_2_33.INJECT1_0 = "NO";
    defparam sub_37_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_31 (.A0(phase_inc_carrGen[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[32]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11595), .COUT(n11596), .S0(n912), .S1(n911));
    defparam sub_37_add_2_31.INIT0 = 16'h5aaa;
    defparam sub_37_add_2_31.INIT1 = 16'h5aaa;
    defparam sub_37_add_2_31.INJECT1_0 = "NO";
    defparam sub_37_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_29 (.A0(phase_inc_carrGen[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11594), .COUT(n11595), .S0(n914), .S1(n913));
    defparam sub_37_add_2_29.INIT0 = 16'h5555;
    defparam sub_37_add_2_29.INIT1 = 16'h5aaa;
    defparam sub_37_add_2_29.INJECT1_0 = "NO";
    defparam sub_37_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_27 (.A0(phase_inc_carrGen[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11593), .COUT(n11594), .S0(n916), .S1(n915));
    defparam sub_37_add_2_27.INIT0 = 16'h5555;
    defparam sub_37_add_2_27.INIT1 = 16'h5aaa;
    defparam sub_37_add_2_27.INJECT1_0 = "NO";
    defparam sub_37_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_25 (.A0(phase_inc_carrGen[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11592), .COUT(n11593), .S0(n918), .S1(n917));
    defparam sub_37_add_2_25.INIT0 = 16'h5aaa;
    defparam sub_37_add_2_25.INIT1 = 16'h5555;
    defparam sub_37_add_2_25.INJECT1_0 = "NO";
    defparam sub_37_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_23 (.A0(phase_inc_carrGen[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11591), .COUT(n11592), .S0(n920), .S1(n919));
    defparam sub_37_add_2_23.INIT0 = 16'h5555;
    defparam sub_37_add_2_23.INIT1 = 16'h5555;
    defparam sub_37_add_2_23.INJECT1_0 = "NO";
    defparam sub_37_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_21 (.A0(phase_inc_carrGen[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11590), .COUT(n11591), .S0(n922), .S1(n921));
    defparam sub_37_add_2_21.INIT0 = 16'h5555;
    defparam sub_37_add_2_21.INIT1 = 16'h5555;
    defparam sub_37_add_2_21.INJECT1_0 = "NO";
    defparam sub_37_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_19 (.A0(phase_inc_carrGen[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11589), .COUT(n11590), .S0(n924), .S1(n923));
    defparam sub_37_add_2_19.INIT0 = 16'h5aaa;
    defparam sub_37_add_2_19.INIT1 = 16'h5aaa;
    defparam sub_37_add_2_19.INJECT1_0 = "NO";
    defparam sub_37_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_17 (.A0(phase_inc_carrGen[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11588), .COUT(n11589), .S0(n926), .S1(n925));
    defparam sub_37_add_2_17.INIT0 = 16'h5aaa;
    defparam sub_37_add_2_17.INIT1 = 16'h5aaa;
    defparam sub_37_add_2_17.INJECT1_0 = "NO";
    defparam sub_37_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_15 (.A0(phase_inc_carrGen[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11587), .COUT(n11588), .S0(n928), .S1(n927));
    defparam sub_37_add_2_15.INIT0 = 16'h5aaa;
    defparam sub_37_add_2_15.INIT1 = 16'h5aaa;
    defparam sub_37_add_2_15.INJECT1_0 = "NO";
    defparam sub_37_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_13 (.A0(phase_inc_carrGen[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11586), .COUT(n11587), .S0(n930), .S1(n929));
    defparam sub_37_add_2_13.INIT0 = 16'h5aaa;
    defparam sub_37_add_2_13.INIT1 = 16'h5aaa;
    defparam sub_37_add_2_13.INJECT1_0 = "NO";
    defparam sub_37_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_11 (.A0(phase_inc_carrGen[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11585), .COUT(n11586), .S0(n932), .S1(n931));
    defparam sub_37_add_2_11.INIT0 = 16'h5555;
    defparam sub_37_add_2_11.INIT1 = 16'h5aaa;
    defparam sub_37_add_2_11.INJECT1_0 = "NO";
    defparam sub_37_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_9 (.A0(phase_inc_carrGen[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11584), .COUT(n11585), .S0(n934), .S1(n933));
    defparam sub_37_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_37_add_2_9.INIT1 = 16'h5555;
    defparam sub_37_add_2_9.INJECT1_0 = "NO";
    defparam sub_37_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_7 (.A0(phase_inc_carrGen[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11583), .COUT(n11584), .S0(n936), .S1(n935));
    defparam sub_37_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_37_add_2_7.INIT1 = 16'h5555;
    defparam sub_37_add_2_7.INJECT1_0 = "NO";
    defparam sub_37_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_5 (.A0(phase_inc_carrGen[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11582), .COUT(n11583), .S0(n938), .S1(n937));
    defparam sub_37_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_37_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_37_add_2_5.INJECT1_0 = "NO";
    defparam sub_37_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_3 (.A0(phase_inc_carrGen[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11581), .COUT(n11582), .S0(n940), .S1(n939));
    defparam sub_37_add_2_3.INIT0 = 16'h5555;
    defparam sub_37_add_2_3.INIT1 = 16'h5555;
    defparam sub_37_add_2_3.INJECT1_0 = "NO";
    defparam sub_37_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_37_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(phase_inc_carrGen[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n11581), .S1(n941));
    defparam sub_37_add_2_1.INIT0 = 16'hF000;
    defparam sub_37_add_2_1.INIT1 = 16'h5555;
    defparam sub_37_add_2_1.INJECT1_0 = "NO";
    defparam sub_37_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_61 (.A0(phase_inc_carrGen[62]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[63]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11579), .S0(n944), .S1(n943));
    defparam sub_38_add_2_61.INIT0 = 16'h5555;
    defparam sub_38_add_2_61.INIT1 = 16'h5555;
    defparam sub_38_add_2_61.INJECT1_0 = "NO";
    defparam sub_38_add_2_61.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_59 (.A0(phase_inc_carrGen[60]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[61]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11578), .COUT(n11579), .S0(n946), .S1(n945));
    defparam sub_38_add_2_59.INIT0 = 16'h5555;
    defparam sub_38_add_2_59.INIT1 = 16'h5555;
    defparam sub_38_add_2_59.INJECT1_0 = "NO";
    defparam sub_38_add_2_59.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_57 (.A0(phase_inc_carrGen[58]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[59]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11577), .COUT(n11578), .S0(n948), .S1(n947));
    defparam sub_38_add_2_57.INIT0 = 16'h5555;
    defparam sub_38_add_2_57.INIT1 = 16'h5555;
    defparam sub_38_add_2_57.INJECT1_0 = "NO";
    defparam sub_38_add_2_57.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_55 (.A0(phase_inc_carrGen[56]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[57]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11576), .COUT(n11577), .S0(n950), .S1(n949));
    defparam sub_38_add_2_55.INIT0 = 16'h5555;
    defparam sub_38_add_2_55.INIT1 = 16'h5555;
    defparam sub_38_add_2_55.INJECT1_0 = "NO";
    defparam sub_38_add_2_55.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_53 (.A0(phase_inc_carrGen[54]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[55]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11575), .COUT(n11576), .S0(n952), .S1(n951));
    defparam sub_38_add_2_53.INIT0 = 16'h5555;
    defparam sub_38_add_2_53.INIT1 = 16'h5555;
    defparam sub_38_add_2_53.INJECT1_0 = "NO";
    defparam sub_38_add_2_53.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_51 (.A0(phase_inc_carrGen[52]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[53]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11574), .COUT(n11575), .S0(n954), .S1(n953));
    defparam sub_38_add_2_51.INIT0 = 16'h5555;
    defparam sub_38_add_2_51.INIT1 = 16'h5555;
    defparam sub_38_add_2_51.INJECT1_0 = "NO";
    defparam sub_38_add_2_51.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_49 (.A0(phase_inc_carrGen[50]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[51]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11573), .COUT(n11574), .S0(n956), .S1(n955));
    defparam sub_38_add_2_49.INIT0 = 16'h5555;
    defparam sub_38_add_2_49.INIT1 = 16'h5555;
    defparam sub_38_add_2_49.INJECT1_0 = "NO";
    defparam sub_38_add_2_49.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_47 (.A0(phase_inc_carrGen[48]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[49]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11572), .COUT(n11573), .S0(n958), .S1(n957));
    defparam sub_38_add_2_47.INIT0 = 16'h5555;
    defparam sub_38_add_2_47.INIT1 = 16'h5555;
    defparam sub_38_add_2_47.INJECT1_0 = "NO";
    defparam sub_38_add_2_47.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_45 (.A0(phase_inc_carrGen[46]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[47]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11571), .COUT(n11572), .S0(n960), .S1(n959));
    defparam sub_38_add_2_45.INIT0 = 16'h5555;
    defparam sub_38_add_2_45.INIT1 = 16'h5555;
    defparam sub_38_add_2_45.INJECT1_0 = "NO";
    defparam sub_38_add_2_45.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_43 (.A0(phase_inc_carrGen[44]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[45]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11570), .COUT(n11571), .S0(n962), .S1(n961));
    defparam sub_38_add_2_43.INIT0 = 16'h5aaa;
    defparam sub_38_add_2_43.INIT1 = 16'h5555;
    defparam sub_38_add_2_43.INJECT1_0 = "NO";
    defparam sub_38_add_2_43.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_41 (.A0(phase_inc_carrGen[42]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[43]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11569), .COUT(n11570), .S0(n964), .S1(n963));
    defparam sub_38_add_2_41.INIT0 = 16'h5aaa;
    defparam sub_38_add_2_41.INIT1 = 16'h5555;
    defparam sub_38_add_2_41.INJECT1_0 = "NO";
    defparam sub_38_add_2_41.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_39 (.A0(phase_inc_carrGen[40]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[41]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11568), .COUT(n11569), .S0(n966), .S1(n965));
    defparam sub_38_add_2_39.INIT0 = 16'h5555;
    defparam sub_38_add_2_39.INIT1 = 16'h5555;
    defparam sub_38_add_2_39.INJECT1_0 = "NO";
    defparam sub_38_add_2_39.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_37 (.A0(phase_inc_carrGen[38]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[39]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11567), .COUT(n11568), .S0(n968), .S1(n967));
    defparam sub_38_add_2_37.INIT0 = 16'h5aaa;
    defparam sub_38_add_2_37.INIT1 = 16'h5aaa;
    defparam sub_38_add_2_37.INJECT1_0 = "NO";
    defparam sub_38_add_2_37.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_35 (.A0(phase_inc_carrGen[36]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[37]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11566), .COUT(n11567), .S0(n970), .S1(n969));
    defparam sub_38_add_2_35.INIT0 = 16'h5aaa;
    defparam sub_38_add_2_35.INIT1 = 16'h5aaa;
    defparam sub_38_add_2_35.INJECT1_0 = "NO";
    defparam sub_38_add_2_35.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_33 (.A0(phase_inc_carrGen[34]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[35]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11565), .COUT(n11566), .S0(n972), .S1(n971));
    defparam sub_38_add_2_33.INIT0 = 16'h5555;
    defparam sub_38_add_2_33.INIT1 = 16'h5aaa;
    defparam sub_38_add_2_33.INJECT1_0 = "NO";
    defparam sub_38_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_31 (.A0(phase_inc_carrGen[32]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[33]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11564), .COUT(n11565), .S0(n974), .S1(n973));
    defparam sub_38_add_2_31.INIT0 = 16'h5555;
    defparam sub_38_add_2_31.INIT1 = 16'h5555;
    defparam sub_38_add_2_31.INJECT1_0 = "NO";
    defparam sub_38_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_29 (.A0(phase_inc_carrGen[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11563), .COUT(n11564), .S0(n976), .S1(n975));
    defparam sub_38_add_2_29.INIT0 = 16'h5555;
    defparam sub_38_add_2_29.INIT1 = 16'h5aaa;
    defparam sub_38_add_2_29.INJECT1_0 = "NO";
    defparam sub_38_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_27 (.A0(phase_inc_carrGen[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11562), .COUT(n11563), .S0(n978), .S1(n977));
    defparam sub_38_add_2_27.INIT0 = 16'h5aaa;
    defparam sub_38_add_2_27.INIT1 = 16'h5aaa;
    defparam sub_38_add_2_27.INJECT1_0 = "NO";
    defparam sub_38_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_25 (.A0(phase_inc_carrGen[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11561), .COUT(n11562), .S0(n980), .S1(n979));
    defparam sub_38_add_2_25.INIT0 = 16'h5aaa;
    defparam sub_38_add_2_25.INIT1 = 16'h5555;
    defparam sub_38_add_2_25.INJECT1_0 = "NO";
    defparam sub_38_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_23 (.A0(phase_inc_carrGen[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11560), .COUT(n11561), .S0(n982), .S1(n981));
    defparam sub_38_add_2_23.INIT0 = 16'h5aaa;
    defparam sub_38_add_2_23.INIT1 = 16'h5555;
    defparam sub_38_add_2_23.INJECT1_0 = "NO";
    defparam sub_38_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_21 (.A0(phase_inc_carrGen[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11559), .COUT(n11560), .S0(n984), .S1(n983));
    defparam sub_38_add_2_21.INIT0 = 16'h5555;
    defparam sub_38_add_2_21.INIT1 = 16'h5aaa;
    defparam sub_38_add_2_21.INJECT1_0 = "NO";
    defparam sub_38_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_19 (.A0(phase_inc_carrGen[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11558), .COUT(n11559), .S0(n986), .S1(n985));
    defparam sub_38_add_2_19.INIT0 = 16'h5555;
    defparam sub_38_add_2_19.INIT1 = 16'h5555;
    defparam sub_38_add_2_19.INJECT1_0 = "NO";
    defparam sub_38_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_17 (.A0(phase_inc_carrGen[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11557), .COUT(n11558), .S0(n988), .S1(n987));
    defparam sub_38_add_2_17.INIT0 = 16'h5555;
    defparam sub_38_add_2_17.INIT1 = 16'h5aaa;
    defparam sub_38_add_2_17.INJECT1_0 = "NO";
    defparam sub_38_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_15 (.A0(phase_inc_carrGen[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11556), .COUT(n11557), .S0(n990), .S1(n989));
    defparam sub_38_add_2_15.INIT0 = 16'h5555;
    defparam sub_38_add_2_15.INIT1 = 16'h5555;
    defparam sub_38_add_2_15.INJECT1_0 = "NO";
    defparam sub_38_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_13 (.A0(phase_inc_carrGen[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11555), .COUT(n11556), .S0(n992), .S1(n991));
    defparam sub_38_add_2_13.INIT0 = 16'h5aaa;
    defparam sub_38_add_2_13.INIT1 = 16'h5aaa;
    defparam sub_38_add_2_13.INJECT1_0 = "NO";
    defparam sub_38_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_11 (.A0(phase_inc_carrGen[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11554), .COUT(n11555), .S0(n994), .S1(n993));
    defparam sub_38_add_2_11.INIT0 = 16'h5555;
    defparam sub_38_add_2_11.INIT1 = 16'h5aaa;
    defparam sub_38_add_2_11.INJECT1_0 = "NO";
    defparam sub_38_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_9 (.A0(phase_inc_carrGen[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11553), .COUT(n11554), .S0(n996), .S1(n995));
    defparam sub_38_add_2_9.INIT0 = 16'h5555;
    defparam sub_38_add_2_9.INIT1 = 16'h5555;
    defparam sub_38_add_2_9.INJECT1_0 = "NO";
    defparam sub_38_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_7 (.A0(phase_inc_carrGen[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11552), .COUT(n11553), .S0(n998), .S1(n997));
    defparam sub_38_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_38_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_38_add_2_7.INJECT1_0 = "NO";
    defparam sub_38_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_5 (.A0(phase_inc_carrGen[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11551), .COUT(n11552), .S0(n1000), .S1(n999));
    defparam sub_38_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_38_add_2_5.INIT1 = 16'h5555;
    defparam sub_38_add_2_5.INJECT1_0 = "NO";
    defparam sub_38_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_3 (.A0(phase_inc_carrGen[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11550), .COUT(n11551), .S0(n1002), .S1(n1001));
    defparam sub_38_add_2_3.INIT0 = 16'h5555;
    defparam sub_38_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_38_add_2_3.INJECT1_0 = "NO";
    defparam sub_38_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_38_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(phase_inc_carrGen[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n11550), .S1(n1003));
    defparam sub_38_add_2_1.INIT0 = 16'hF000;
    defparam sub_38_add_2_1.INIT1 = 16'h5555;
    defparam sub_38_add_2_1.INJECT1_0 = "NO";
    defparam sub_38_add_2_1.INJECT1_1 = "NO";
    LUT4 mux_378_i13_3_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), 
         .C(o_Rx_Byte_c_3), .D(n2596), .Z(n2727)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i13_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_378_i20_4_lut_else_4_lut (.A(o_Rx_Byte_c_2), .B(o_Rx_Byte_c_3), 
         .C(n7319), .D(o_Rx_Byte_c_0), .Z(n13810)) /* synthesis lut_function=(!(A (B (C)+!B (D))+!A (B (C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i20_4_lut_else_4_lut.init = 16'h1d3f;
    LUT4 mux_367_i41_4_lut (.A(n2699), .B(n966), .C(n2215), .D(n13757), 
         .Z(n2240)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i41_4_lut.init = 16'hcfca;
    LUT4 mux_378_i41_4_lut (.A(o_Rx_Byte_c_2), .B(n7319), .C(o_Rx_Byte_c_3), 
         .D(n903), .Z(n2699)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(B+!(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i41_4_lut.init = 16'h9a1a;
    LUT4 mux_367_i42_4_lut (.A(n2698), .B(n965), .C(n2215), .D(n13757), 
         .Z(n2239)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i42_4_lut.init = 16'hcfca;
    LUT4 mux_367_i63_4_lut (.A(n881), .B(n944), .C(n2215), .D(n7986), 
         .Z(n2218)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i63_4_lut.init = 16'hcac0;
    LUT4 mux_375_i42_3_lut (.A(n7319), .B(n902), .C(o_Rx_Byte_c_2), .Z(n2567)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_375_i42_3_lut.init = 16'hdada;
    LUT4 mux_378_i55_4_lut_then_4_lut (.A(o_Rx_Byte_c_2), .B(o_Rx_Byte_c_3), 
         .C(n7319), .D(o_Rx_Byte_c_0), .Z(n13775)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i55_4_lut_then_4_lut.init = 16'he2c0;
    LUT4 mux_367_i39_4_lut (.A(n2701), .B(n968), .C(n2215), .D(n13757), 
         .Z(n2242)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i39_4_lut.init = 16'hc0ca;
    LUT4 mux_375_i39_3_lut (.A(n7319), .B(n905), .C(o_Rx_Byte_c_2), .Z(n2570)) /* synthesis lut_function=(A (B (C))+!A !(C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_375_i39_3_lut.init = 16'h8585;
    LUT4 mux_367_i40_4_lut (.A(n2700), .B(n967), .C(n2215), .D(n13757), 
         .Z(n2241)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i40_4_lut.init = 16'hcfca;
    LUT4 mux_367_i64_4_lut (.A(n880), .B(n943), .C(n2215), .D(n7986), 
         .Z(n2217)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i64_4_lut.init = 16'hcac0;
    LUT4 i2799_4_lut (.A(n7319), .B(o_Rx_Byte_c_3), .C(n904), .D(o_Rx_Byte_c_2), 
         .Z(n2700)) /* synthesis lut_function=(A (B (C (D)))+!A !((D)+!B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i2799_4_lut.init = 16'h8044;
    LUT4 mux_367_i61_4_lut (.A(n2548), .B(n946), .C(n2215), .D(n13753), 
         .Z(n2220)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i61_4_lut.init = 16'hcac0;
    LUT4 mux_378_i24_4_lut_then_4_lut (.A(o_Rx_Byte_c_2), .B(o_Rx_Byte_c_3), 
         .C(n7319), .D(o_Rx_Byte_c_0), .Z(n13817)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i24_4_lut_then_4_lut.init = 16'hd1c0;
    LUT4 mux_378_i24_4_lut_else_4_lut (.A(o_Rx_Byte_c_2), .B(o_Rx_Byte_c_3), 
         .C(n7319), .D(o_Rx_Byte_c_0), .Z(n13816)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i24_4_lut_else_4_lut.init = 16'h5140;
    LUT4 mux_375_i61_3_lut (.A(n7319), .B(n883), .C(o_Rx_Byte_c_2), .Z(n2548)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_375_i61_3_lut.init = 16'hdada;
    LUT4 mux_367_i62_4_lut (.A(n882), .B(n945), .C(n2215), .D(n7986), 
         .Z(n2219)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i62_4_lut.init = 16'hcac0;
    LUT4 mux_367_i37_4_lut (.A(n7695), .B(n970), .C(n2215), .D(n13757), 
         .Z(n2244)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i37_4_lut.init = 16'hc0ca;
    LUT4 mux_367_i59_4_lut (.A(n2681), .B(n948), .C(n2215), .D(n13757), 
         .Z(n2222)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i59_4_lut.init = 16'hc0ca;
    \CIC(width=72,decimation_ratio=4096)  CIC1Sin (.osc_clk(osc_clk), .\CICGain[1] (CICGain[1]), 
            .\CICGain[0] (CICGain[0]), .CIC1_out_clkSin(CIC1_out_clkSin), 
            .\CIC1_outSin[0] (CIC1_outSin[0]), .MixerOutSin({MixerOutSin}), 
            .GND_net(GND_net), .\CIC1_outSin[1] (CIC1_outSin[1]), .\CIC1_outSin[2] (CIC1_outSin[2]), 
            .\CIC1_outSin[3] (CIC1_outSin[3]), .\CIC1_outSin[4] (CIC1_outSin[4]), 
            .\CIC1_outSin[5] (CIC1_outSin[5]), .MYLED_c_0(MYLED_c_0), .MYLED_c_1(MYLED_c_1), 
            .MYLED_c_2(MYLED_c_2), .MYLED_c_3(MYLED_c_3), .MYLED_c_4(MYLED_c_4), 
            .MYLED_c_5(MYLED_c_5), .\d10[67] (d10_adj_2639[67]), .\d10[68] (d10_adj_2639[68]), 
            .\d10[69] (d10_adj_2639[69]), .\d10[70] (d10_adj_2639[70]), 
            .n63(n63), .\d_out_11__N_1818[2] (d_out_11__N_1818_adj_2663[2]), 
            .n64(n64), .\d_out_11__N_1818[3] (d_out_11__N_1818_adj_2663[3]), 
            .n70(n70), .n67(n67), .\d10[65] (d10_adj_2639[65]), .n68(n68), 
            .\d10[66] (d10_adj_2639[66]), .n65(n65), .\d10[63] (d10_adj_2639[63]), 
            .n66(n66), .\d10[64] (d10_adj_2639[64]), .\d10[61] (d10_adj_2639[61]), 
            .\d10[62] (d10_adj_2639[62]), .\d_out_11__N_1818[10] (d_out_11__N_1818_adj_2663[10]), 
            .n61(n61), .\d10[59] (d10_adj_2639[59]), .n62(n62), .\d10[60] (d10_adj_2639[60]), 
            .\d_out_11__N_1818[5] (d_out_11__N_1818_adj_2663[5]), .\d_out_11__N_1818[4] (d_out_11__N_1818_adj_2663[4]), 
            .\d_out_11__N_1818[6] (d_out_11__N_1818_adj_2663[6]), .\d_out_11__N_1818[7] (d_out_11__N_1818_adj_2663[7]), 
            .\d_out_11__N_1818[8] (d_out_11__N_1818_adj_2663[8]), .\d_out_11__N_1818[9] (d_out_11__N_1818_adj_2663[9]), 
            .\d10[71] (d10_adj_2639[71]), .\d_out_11__N_1818[11] (d_out_11__N_1818_adj_2663[11])) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(128[45] 134[2])
    LUT4 mux_375_i59_3_lut (.A(n7319), .B(n885), .C(o_Rx_Byte_c_2), .Z(n2550)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_375_i59_3_lut.init = 16'hdada;
    LUT4 mux_367_i60_4_lut (.A(n884), .B(n947), .C(n2215), .D(n7986), 
         .Z(n2221)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i60_4_lut.init = 16'hcac0;
    LUT4 mux_367_i57_4_lut (.A(n2683), .B(n950), .C(n2215), .D(n13757), 
         .Z(n2224)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i57_4_lut.init = 16'hc0ca;
    LUT4 mux_375_i57_3_lut (.A(n7319), .B(n887), .C(o_Rx_Byte_c_2), .Z(n2552)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_375_i57_3_lut.init = 16'hdada;
    LUT4 i2699_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), .C(n2310), 
         .D(o_Rx_Byte_c_3), .Z(n7695)) /* synthesis lut_function=(A ((C (D))+!B)+!A ((C+!(D))+!B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i2699_4_lut.init = 16'hf377;
    LUT4 i5912_4_lut (.A(n8210), .B(o_Rx_Byte_c_3), .C(o_Rx_Byte_c_6), 
         .D(n6), .Z(osc_clk_enable_1393)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i5912_4_lut.init = 16'h0001;
    LUT4 i1_2_lut (.A(o_Rx_Byte_c_2), .B(o_Rx_Byte_c_4), .Z(n6)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 i2844_2_lut (.A(n907), .B(n7319), .Z(n2310)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i2844_2_lut.init = 16'hbbbb;
    LUT4 mux_367_i38_4_lut (.A(n2702), .B(n969), .C(n2215), .D(n13757), 
         .Z(n2243)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i38_4_lut.init = 16'hcfca;
    LUT4 i2845_2_lut (.A(n906), .B(n7319), .Z(n2309)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i2845_2_lut.init = 16'hbbbb;
    LUT4 mux_367_i35_4_lut (.A(n13151), .B(n972), .C(n2215), .D(n9), 
         .Z(n2246)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i35_4_lut.init = 16'hc5cf;
    LUT4 mux_367_i58_4_lut (.A(n2682), .B(n949), .C(n2215), .D(n13757), 
         .Z(n2223)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i58_4_lut.init = 16'hcfca;
    LUT4 i1_3_lut (.A(n909), .B(o_Rx_Byte_c_3), .C(n7319), .Z(n9)) /* synthesis lut_function=(!(A (B)+!A !((C)+!B))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i1_3_lut.init = 16'h7373;
    LUT4 mux_375_i58_3_lut (.A(n7319), .B(n886), .C(o_Rx_Byte_c_2), .Z(n2551)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_375_i58_3_lut.init = 16'hdada;
    PFUMX i6066 (.BLUT(n13837), .ALUT(n13838), .C0(n895), .Z(n13839));
    PFUMX i6064 (.BLUT(n13822), .ALUT(n13823), .C0(n899), .Z(n13836));
    LUT4 mux_378_i27_4_lut_then_4_lut (.A(o_Rx_Byte_c_2), .B(o_Rx_Byte_c_3), 
         .C(n7319), .D(o_Rx_Byte_c_0), .Z(n13823)) /* synthesis lut_function=(A+!(B (C)+!B (D))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i27_4_lut_then_4_lut.init = 16'haebf;
    LUT4 mux_378_i27_4_lut_else_4_lut (.A(o_Rx_Byte_c_2), .B(o_Rx_Byte_c_3), 
         .C(n7319), .D(o_Rx_Byte_c_0), .Z(n13822)) /* synthesis lut_function=(!(A (B (C))+!A (B (C)+!B (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i27_4_lut_else_4_lut.init = 16'h2e3f;
    PFUMX i6062 (.BLUT(n13831), .ALUT(n13832), .C0(o_Rx_Byte_c_0), .Z(n13833));
    LUT4 i1709_2_lut_rep_170 (.A(n7319), .B(o_Rx_Byte_c_2), .Z(n13763)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i1709_2_lut_rep_170.init = 16'h8888;
    LUT4 mux_367_i36_4_lut (.A(n2704), .B(n971), .C(n2215), .D(n13757), 
         .Z(n2245)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i36_4_lut.init = 16'hcfca;
    LUT4 mux_375_i36_3_lut (.A(n7319), .B(n908), .C(o_Rx_Byte_c_2), .Z(n2573)) /* synthesis lut_function=(A (B (C))+!A !(C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_375_i36_3_lut.init = 16'h8585;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n7319), .B(o_Rx_Byte_c_2), .C(n13757), 
         .D(o_Rx_Byte_c_3), .Z(n7986)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0800;
    LUT4 i1_3_lut_adj_62 (.A(o_Rx_Byte_c_5), .B(o_Rx_DV_c_0), .C(o_Rx_Byte_c_7), 
         .Z(n8210)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_3_lut_adj_62.init = 16'hf7f7;
    LUT4 mux_367_i55_4_lut (.A(n13776), .B(n952), .C(n2215), .D(n13757), 
         .Z(n2226)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i55_4_lut.init = 16'hcfca;
    LUT4 mux_367_i33_4_lut (.A(n2707), .B(n974), .C(n2215), .D(n13757), 
         .Z(n2248)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i33_4_lut.init = 16'hc0ca;
    LUT4 i2842_2_lut (.A(n911), .B(n7319), .Z(n2314)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i2842_2_lut.init = 16'hbbbb;
    LUT4 mux_367_i34_4_lut (.A(n14103), .B(n973), .C(n2215), .D(n13757), 
         .Z(n2247)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i34_4_lut.init = 16'hcfca;
    PFUMX i6056 (.BLUT(n13822), .ALUT(n13823), .C0(n917), .Z(n13824));
    LUT4 mux_367_i31_4_lut (.A(n2709), .B(n976), .C(n2215), .D(n13757), 
         .Z(n2250)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i31_4_lut.init = 16'hc0ca;
    LUT4 i2840_2_lut (.A(n913), .B(n7319), .Z(n2316)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i2840_2_lut.init = 16'h8888;
    LUT4 mux_378_i7_4_lut_else_4_lut (.A(n937), .B(o_Rx_Byte_c_3), .C(o_Rx_Byte_c_2), 
         .D(n7319), .Z(n14095)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i7_4_lut_else_4_lut.init = 16'h8000;
    PFUMX i6052 (.BLUT(n13816), .ALUT(n13817), .C0(n920), .Z(n13818));
    PFUMX i6175 (.BLUT(n14095), .ALUT(n14096), .C0(o_Rx_Byte_c_0), .Z(n14097));
    LUT4 mux_367_i32_4_lut (.A(n2708), .B(n975), .C(n2215), .D(n13757), 
         .Z(n2249)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i32_4_lut.init = 16'hc0ca;
    PFUMX i6050 (.BLUT(n13822), .ALUT(n13823), .C0(n925), .Z(n13815));
    LUT4 mux_378_i43_4_lut_then_4_lut (.A(n901), .B(o_Rx_Byte_c_3), .C(o_Rx_Byte_c_2), 
         .D(n7319), .Z(n13832)) /* synthesis lut_function=(A (B+(C))+!A !(B (C (D))+!B !(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i43_4_lut_then_4_lut.init = 16'hbcfc;
    LUT4 mux_378_i43_4_lut_else_4_lut (.A(n901), .B(o_Rx_Byte_c_3), .C(o_Rx_Byte_c_2), 
         .D(n7319), .Z(n13831)) /* synthesis lut_function=(A (B+!(C))+!A !(B (C (D))+!B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i43_4_lut_else_4_lut.init = 16'h8fcf;
    PFUMX i6048 (.BLUT(n13810), .ALUT(n13811), .C0(n924), .Z(n13812));
    LUT4 mux_367_i56_4_lut (.A(n8992), .B(n951), .C(n2215), .D(n12946), 
         .Z(n2225)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i56_4_lut.init = 16'hcacf;
    LUT4 mux_375_i32_3_lut (.A(n7319), .B(n912), .C(o_Rx_Byte_c_2), .Z(n2577)) /* synthesis lut_function=(A (B (C))+!A !(C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_375_i32_3_lut.init = 16'h8585;
    LUT4 mux_367_i29_4_lut (.A(n2711), .B(n978), .C(n2215), .D(n13757), 
         .Z(n2252)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i29_4_lut.init = 16'hcfca;
    LUT4 mux_375_i29_3_lut (.A(n7319), .B(n915), .C(o_Rx_Byte_c_2), .Z(n2580)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_375_i29_3_lut.init = 16'hdada;
    LUT4 mux_378_i49_4_lut_then_4_lut (.A(o_Rx_Byte_c_2), .B(o_Rx_Byte_c_3), 
         .C(n7319), .D(o_Rx_Byte_c_0), .Z(n13838)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i49_4_lut_then_4_lut.init = 16'hc0e2;
    LUT4 mux_378_i49_4_lut_else_4_lut (.A(o_Rx_Byte_c_2), .B(o_Rx_Byte_c_3), 
         .C(n7319), .D(o_Rx_Byte_c_0), .Z(n13837)) /* synthesis lut_function=(!(A (B+(D))+!A !(B (C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i49_4_lut_else_4_lut.init = 16'h4062;
    LUT4 mux_367_i30_4_lut (.A(n2710), .B(n977), .C(n2215), .D(n13757), 
         .Z(n2251)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i30_4_lut.init = 16'hc0ca;
    LUT4 i2989_2_lut (.A(o_Rx_Byte_c_2), .B(n888), .Z(n8992)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i2989_2_lut.init = 16'h8888;
    PFUMX i6044 (.BLUT(n13804), .ALUT(n13805), .C0(n7319), .Z(n13806));
    LUT4 mux_375_i30_3_lut (.A(n7319), .B(n914), .C(o_Rx_Byte_c_2), .Z(n2579)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_375_i30_3_lut.init = 16'hdada;
    PFUMX i6042 (.BLUT(n13801), .ALUT(n13802), .C0(o_Rx_Byte_c_0), .Z(n13803));
    LUT4 mux_367_i27_4_lut (.A(n13824), .B(n980), .C(n2215), .D(n13757), 
         .Z(n2254)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i27_4_lut.init = 16'hcfca;
    LUT4 mux_367_i28_4_lut (.A(n2712), .B(n979), .C(n2215), .D(n13757), 
         .Z(n2253)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i28_4_lut.init = 16'hc0ca;
    PLL PLL1 (.XIn_c(XIn_c), .osc_clk(osc_clk), .GND_net(GND_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(154[5] 156[2])
    PFUMX i6038 (.BLUT(n13795), .ALUT(n13796), .C0(n934), .Z(n13797));
    LUT4 i5863_4_lut (.A(n9004), .B(n7986), .C(osc_clk_enable_1457), .D(n2215), 
         .Z(osc_clk_enable_1458)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i5863_4_lut.init = 16'h0010;
    LUT4 mux_375_i28_3_lut (.A(n7319), .B(n916), .C(o_Rx_Byte_c_2), .Z(n2581)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_375_i28_3_lut.init = 16'hdada;
    LUT4 mux_378_i22_4_lut_then_4_lut (.A(n922), .B(o_Rx_Byte_c_3), .C(o_Rx_Byte_c_2), 
         .D(n7319), .Z(n14099)) /* synthesis lut_function=(A (B+(C))+!A !(B (C (D))+!B !(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i22_4_lut_then_4_lut.init = 16'hbcfc;
    LUT4 i5_4_lut (.A(n9_adj_2616), .B(n7), .C(n13757), .D(n13767), 
         .Z(n8366)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut.init = 16'h8000;
    LUT4 mux_367_i25_4_lut (.A(n2715), .B(n982), .C(n2215), .D(n13757), 
         .Z(n2256)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i25_4_lut.init = 16'hc0ca;
    LUT4 i3_2_lut (.A(o_Rx_Byte_c_6), .B(n41), .Z(n9_adj_2616)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    PFUMX i6036 (.BLUT(n13792), .ALUT(n13793), .C0(n7319), .Z(n41));
    LUT4 i1_2_lut_adj_63 (.A(n9004), .B(n2215), .Z(n7)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i1_2_lut_adj_63.init = 16'h1111;
    PFUMX i6034 (.BLUT(n13810), .ALUT(n13811), .C0(n939), .Z(n13791));
    LUT4 i2798_4_lut (.A(n919), .B(o_Rx_Byte_c_3), .C(o_Rx_Byte_c_2), 
         .D(n7319), .Z(n2715)) /* synthesis lut_function=(A ((C)+!B)+!A !(B ((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i2798_4_lut.init = 16'hb3f3;
    LUT4 mux_367_i26_4_lut (.A(n2714), .B(n981), .C(n2215), .D(n13757), 
         .Z(n2255)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i26_4_lut.init = 16'hc0ca;
    LUT4 mux_378_i26_4_lut (.A(o_Rx_Byte_c_0), .B(n918), .C(o_Rx_Byte_c_3), 
         .D(n13763), .Z(n2714)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B+!(C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i26_4_lut.init = 16'hc5f5;
    LUT4 mux_367_i23_4_lut (.A(n2717), .B(n984), .C(n2215), .D(n13757), 
         .Z(n2258)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i23_4_lut.init = 16'hcfca;
    LUT4 mux_375_i23_3_lut (.A(n7319), .B(n921), .C(o_Rx_Byte_c_2), .Z(n2586)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_375_i23_3_lut.init = 16'hdada;
    PFUMX i6032 (.BLUT(n13837), .ALUT(n13838), .C0(n938), .Z(n13788));
    LUT4 mux_367_i24_4_lut (.A(n13818), .B(n983), .C(n2215), .D(n13757), 
         .Z(n2257)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i24_4_lut.init = 16'hc0ca;
    LUT4 mux_367_i21_4_lut (.A(n8980), .B(n986), .C(n2215), .D(n12946), 
         .Z(n2260)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i21_4_lut.init = 16'hcacf;
    LUT4 i2977_2_lut (.A(o_Rx_Byte_c_2), .B(n923), .Z(n8980)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i2977_2_lut.init = 16'h8888;
    FD1P3AX phase_inc_carrGen_i0_i2 (.D(n2936), .SP(osc_clk_enable_1396), 
            .CK(osc_clk), .Q(phase_inc_carrGen[2]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i2.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i3 (.D(n2935), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[3]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i3.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i4 (.D(n2934), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[4]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i4.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i5 (.D(n2933), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[5]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i5.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i6 (.D(n2932), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[6]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i6.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i7 (.D(n2931), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[7]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i7.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i8 (.D(n2930), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[8]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i8.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i9 (.D(n2929), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[9]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i9.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i10 (.D(n2928), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[10]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i10.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i11 (.D(n2927), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[11]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i11.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i12 (.D(n2926), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[12]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i12.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i13 (.D(n2925), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[13]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i13.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i14 (.D(n2924), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[14]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i14.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i15 (.D(n2923), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[15]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i15.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i16 (.D(n2922), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[16]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i16.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i17 (.D(n2921), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[17]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i17.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i18 (.D(n2920), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[18]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i18.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i19 (.D(n2919), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[19]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i19.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i20 (.D(n2918), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[20]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i20.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i21 (.D(n2917), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[21]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i21.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i22 (.D(n2916), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[22]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i22.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i23 (.D(n2915), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[23]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i23.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i24 (.D(n2914), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[24]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i24.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i25 (.D(n2913), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[25]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i25.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i26 (.D(n2912), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[26]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i26.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i27 (.D(n2911), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[27]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i27.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i28 (.D(n2910), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[28]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i28.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i29 (.D(n2909), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[29]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i29.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i30 (.D(n2908), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[30]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i30.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i31 (.D(n2907), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[31]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i31.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i32 (.D(n2906), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[32]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i32.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i33 (.D(n2905), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[33]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i33.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i34 (.D(n2904), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[34]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i34.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i35 (.D(n2903), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[35]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i35.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i36 (.D(n2902), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[36]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i36.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i37 (.D(n2901), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[37]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i37.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i38 (.D(n2900), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[38]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i38.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i39 (.D(n2899), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[39]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i39.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i40 (.D(n2898), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[40]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i40.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i41 (.D(n2897), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[41]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i41.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i42 (.D(n2896), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[42]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i42.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i43 (.D(n2895), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[43]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i43.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i44 (.D(n2894), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[44]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i44.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i45 (.D(n2893), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[45]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i45.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i46 (.D(n2892), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[46]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i46.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i47 (.D(n2891), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[47]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i47.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i48 (.D(n2890), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[48]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i48.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i49 (.D(n2889), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[49]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i49.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i50 (.D(n2888), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[50]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i50.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i51 (.D(n2887), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[51]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i51.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i52 (.D(n2886), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[52]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i52.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i53 (.D(n2885), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[53]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i53.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i54 (.D(n2884), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[54]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i54.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i55 (.D(n2883), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[55]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i55.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i56 (.D(n2882), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[56]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i56.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i57 (.D(n2881), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[57]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i57.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i58 (.D(n2880), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[58]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i58.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i59 (.D(n2879), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[59]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i59.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i60 (.D(n2878), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[60]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i60.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i61 (.D(n2877), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[61]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i61.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i62 (.D(n2876), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[62]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i62.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i63 (.D(n2875), .SP(osc_clk_enable_1457), 
            .CK(osc_clk), .Q(phase_inc_carrGen[63]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i63.GSR = "ENABLED";
    LUT4 mux_367_i22_4_lut (.A(n14100), .B(n985), .C(n2215), .D(n13757), 
         .Z(n2259)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i22_4_lut.init = 16'hcfca;
    PFUMX i6030 (.BLUT(n13783), .ALUT(n13775), .C0(n940), .Z(n13785));
    LUT4 mux_367_i19_4_lut (.A(n13815), .B(n988), .C(n2215), .D(n13757), 
         .Z(n2262)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i19_4_lut.init = 16'hc0ca;
    PFUMX i6179 (.BLUT(n14101), .ALUT(n14102), .C0(o_Rx_Byte_c_0), .Z(n14103));
    LUT4 i2355_2_lut (.A(o_Rx_Byte_c_2), .B(o_Rx_Byte_c_3), .Z(n2738)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i2355_2_lut.init = 16'h6666;
    GSR GSR_INST (.GSR(VCC_net));
    LUT4 mux_367_i20_4_lut (.A(n13812), .B(n987), .C(n2215), .D(n13757), 
         .Z(n2261)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i20_4_lut.init = 16'hcfca;
    TSALL TSALL_INST (.TSALL(GND_net));
    LUT4 mux_367_i17_4_lut (.A(n2723), .B(n990), .C(n2215), .D(n13757), 
         .Z(n2264)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i17_4_lut.init = 16'hc0ca;
    LUT4 mux_378_i17_4_lut (.A(o_Rx_Byte_c_0), .B(n2330), .C(o_Rx_Byte_c_3), 
         .D(o_Rx_Byte_c_2), .Z(n2723)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i17_4_lut.init = 16'hcafa;
    LUT4 i2828_2_lut (.A(n927), .B(n7319), .Z(n2330)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i2828_2_lut.init = 16'h8888;
    LUT4 mux_367_i18_4_lut (.A(n2722), .B(n989), .C(n2215), .D(n13757), 
         .Z(n2263)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i18_4_lut.init = 16'hcfca;
    LUT4 mux_375_i18_3_lut (.A(n7319), .B(n926), .C(o_Rx_Byte_c_2), .Z(n2591)) /* synthesis lut_function=(A (B (C))+!A !(C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_375_i18_3_lut.init = 16'h8585;
    LUT4 i5489_2_lut_rep_172 (.A(n7319), .B(o_Rx_Byte_c_4), .Z(n13765)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i5489_2_lut_rep_172.init = 16'heeee;
    LUT4 mux_367_i15_4_lut (.A(n2725), .B(n992), .C(n2215), .D(n13757), 
         .Z(n2266)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i15_4_lut.init = 16'hcfca;
    LUT4 mux_375_i15_3_lut (.A(n7319), .B(n929), .C(o_Rx_Byte_c_2), .Z(n2594)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_375_i15_3_lut.init = 16'hdada;
    LUT4 i1_3_lut_rep_164_4_lut (.A(n7319), .B(o_Rx_Byte_c_4), .C(o_Rx_Byte_c_0), 
         .D(n12872), .Z(n13757)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_3_lut_rep_164_4_lut.init = 16'h1000;
    LUT4 mux_367_i16_4_lut (.A(n2724), .B(n991), .C(n2215), .D(n13757), 
         .Z(n2265)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i16_4_lut.init = 16'hcfca;
    LUT4 mux_378_i16_4_lut (.A(o_Rx_Byte_c_0), .B(n2331), .C(o_Rx_Byte_c_3), 
         .D(o_Rx_Byte_c_2), .Z(n2724)) /* synthesis lut_function=(A (B (C (D)))+!A (B ((D)+!C)+!B !(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i16_4_lut.init = 16'hc505;
    LUT4 i2827_2_lut (.A(n928), .B(n7319), .Z(n2331)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i2827_2_lut.init = 16'hbbbb;
    LUT4 mux_367_i13_4_lut (.A(n2727), .B(n994), .C(n2215), .D(n13757), 
         .Z(n2268)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i13_4_lut.init = 16'hc0ca;
    LUT4 mux_375_i13_3_lut (.A(n7319), .B(n931), .C(o_Rx_Byte_c_2), .Z(n2596)) /* synthesis lut_function=(A (B (C))+!A !(C)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_375_i13_3_lut.init = 16'h8585;
    nco_sig ncoGen (.osc_clk(osc_clk), .\phase_accum[63] (phase_accum[63]), 
            .\phase_accum[62] (phase_accum[62]), .\phase_accum[61] (phase_accum[61]), 
            .\phase_accum[60] (phase_accum[60]), .\phase_accum[59] (phase_accum[59]), 
            .\phase_accum[58] (phase_accum[58]), .\phase_accum[57] (phase_accum[57]), 
            .\phase_accum[56] (phase_accum[56]), .sinGen_c(sinGen_c), .phase_inc_carrGen1({phase_inc_carrGen1}), 
            .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(108[10] 114[2])
    LUT4 i5897_4_lut (.A(n13806), .B(n12896), .C(o_Rx_Byte_c_4), .D(n57), 
         .Z(n9004)) /* synthesis lut_function=(!(A (B)+!A !((C+!(D))+!B))) */ ;
    defparam i5897_4_lut.init = 16'h7377;
    LUT4 i1_3_lut_rep_174 (.A(o_Rx_Byte_c_5), .B(o_Rx_DV_c_0), .C(o_Rx_Byte_c_7), 
         .Z(n13767)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_3_lut_rep_174.init = 16'h0808;
    LUT4 i1_2_lut_4_lut (.A(o_Rx_Byte_c_5), .B(o_Rx_DV_c_0), .C(o_Rx_Byte_c_7), 
         .D(o_Rx_Byte_c_6), .Z(n12896)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0800;
    LUT4 mux_367_i14_4_lut (.A(n2595), .B(n993), .C(n2215), .D(n13753), 
         .Z(n2267)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i14_4_lut.init = 16'hcacf;
    PFUMX i6177 (.BLUT(n14098), .ALUT(n14099), .C0(o_Rx_Byte_c_0), .Z(n14100));
    LUT4 i2802_3_lut (.A(n930), .B(o_Rx_Byte_c_2), .C(n7319), .Z(n2595)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam i2802_3_lut.init = 16'h8c8c;
    LUT4 mux_367_i11_4_lut (.A(n13803), .B(n996), .C(n2215), .D(n13757), 
         .Z(n2270)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i11_4_lut.init = 16'hc0ca;
    LUT4 i74_4_lut (.A(o_Rx_Byte_c_0), .B(n7319), .C(o_Rx_Byte_c_2), .D(o_Rx_Byte_c_3), 
         .Z(n57)) /* synthesis lut_function=(!(A (B (C)+!B (D))+!A (B+((D)+!C)))) */ ;
    defparam i74_4_lut.init = 16'h083a;
    \CIC(width=72,decimation_ratio=4096)_U1  CIC1Cos (.GND_net(GND_net), .osc_clk(osc_clk), 
            .CIC1_outCos({CIC1_outCos}), .\d10[59] (d10_adj_2639[59]), .\d10[60] (d10_adj_2639[60]), 
            .\d10[61] (d10_adj_2639[61]), .\d10[62] (d10_adj_2639[62]), 
            .\d10[63] (d10_adj_2639[63]), .\d10[64] (d10_adj_2639[64]), 
            .\d10[65] (d10_adj_2639[65]), .\d10[66] (d10_adj_2639[66]), 
            .\d10[67] (d10_adj_2639[67]), .\d10[68] (d10_adj_2639[68]), 
            .\d10[69] (d10_adj_2639[69]), .\d10[70] (d10_adj_2639[70]), 
            .\d10[71] (d10_adj_2639[71]), .\d_out_11__N_1818[2] (d_out_11__N_1818_adj_2663[2]), 
            .\d_out_11__N_1818[3] (d_out_11__N_1818_adj_2663[3]), .\d_out_11__N_1818[4] (d_out_11__N_1818_adj_2663[4]), 
            .\d_out_11__N_1818[5] (d_out_11__N_1818_adj_2663[5]), .\d_out_11__N_1818[6] (d_out_11__N_1818_adj_2663[6]), 
            .\d_out_11__N_1818[7] (d_out_11__N_1818_adj_2663[7]), .\d_out_11__N_1818[8] (d_out_11__N_1818_adj_2663[8]), 
            .\d_out_11__N_1818[9] (d_out_11__N_1818_adj_2663[9]), .\d_out_11__N_1818[10] (d_out_11__N_1818_adj_2663[10]), 
            .\d_out_11__N_1818[11] (d_out_11__N_1818_adj_2663[11]), .\CICGain[0] (CICGain[0]), 
            .n61(n61), .MixerOutCos({MixerOutCos}), .n62(n62), .n63(n63), 
            .n64(n64), .\CICGain[1] (CICGain[1]), .n65(n65), .n66(n66), 
            .n67(n67), .n68(n68), .n70(n70)) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(137[45] 143[2])
    PFUMX i6024 (.BLUT(n13783), .ALUT(n13775), .C0(n889), .Z(n13776));
    VLO i1 (.Z(GND_net));
    FD1P3JX phase_inc_carrGen_i0_i0 (.D(n2739), .SP(osc_clk_enable_1458), 
            .PD(n8366), .CK(osc_clk), .Q(phase_inc_carrGen[0]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(193[8] 234[4])
    defparam phase_inc_carrGen_i0_i0.GSR = "ENABLED";
    \uart_rx(CLKS_PER_BIT=87)  uart_rx1 (.\UartClk[2] (UartClk_adj_2711[2]), 
            .osc_clk(osc_clk), .i_Rx_Serial_c(i_Rx_Serial_c), .o_Rx_DV_c_0(o_Rx_DV_c_0), 
            .o_Rx_Byte_c_0(o_Rx_Byte_c_0), .n7319(n7319), .o_Rx_Byte_c_2(o_Rx_Byte_c_2), 
            .o_Rx_Byte_c_3(o_Rx_Byte_c_3), .o_Rx_Byte_c_4(o_Rx_Byte_c_4), 
            .o_Rx_Byte_c_5(o_Rx_Byte_c_5), .o_Rx_Byte_c_6(o_Rx_Byte_c_6), 
            .o_Rx_Byte_c_7(o_Rx_Byte_c_7), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(176[32] 181[2])
    LUT4 mux_378_i1_4_lut_4_lut (.A(o_Rx_Byte_c_0), .B(o_Rx_Byte_c_2), .C(o_Rx_Byte_c_3), 
         .D(n7319), .Z(n2739)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (B ((D)+!C)+!B (C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_378_i1_4_lut_4_lut.init = 16'h09c9;
    LUT4 mux_367_i12_4_lut (.A(n2728), .B(n995), .C(n2215), .D(n13757), 
         .Z(n2269)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(197[2] 233[6])
    defparam mux_367_i12_4_lut.init = 16'hc0ca;
    AMDemodulator AMDemodulator1 (.CIC1_out_clkSin(CIC1_out_clkSin), .\CIC1_outSin[0] (CIC1_outSin[0]), 
            .CIC1_outCos({CIC1_outCos}), .\DataInReg_11__N_1855[0] (DataInReg_11__N_1855[0]), 
            .GND_net(GND_net), .\CIC1_outSin[1] (CIC1_outSin[1]), .\CIC1_outSin[2] (CIC1_outSin[2]), 
            .\CIC1_outSin[3] (CIC1_outSin[3]), .\CIC1_outSin[4] (CIC1_outSin[4]), 
            .\CIC1_outSin[5] (CIC1_outSin[5]), .MYLED_c_0(MYLED_c_0), .MYLED_c_1(MYLED_c_1), 
            .MYLED_c_2(MYLED_c_2), .MYLED_c_3(MYLED_c_3), .MYLED_c_4(MYLED_c_4), 
            .MYLED_c_5(MYLED_c_5), .\DataInReg_11__N_1855[1] (DataInReg_11__N_1855[1]), 
            .\DataInReg_11__N_1855[2] (DataInReg_11__N_1855[2]), .\DataInReg_11__N_1855[3] (DataInReg_11__N_1855[3]), 
            .\DataInReg_11__N_1855[4] (DataInReg_11__N_1855[4]), .\DataInReg_11__N_1855[5] (DataInReg_11__N_1855[5]), 
            .\DataInReg_11__N_1855[6] (DataInReg_11__N_1855[6]), .\DataInReg_11__N_1855[7] (DataInReg_11__N_1855[7]), 
            .\DataInReg_11__N_1855[8] (DataInReg_11__N_1855[8]), .\DemodOut[9] (DemodOut[9]), 
            .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(168[15] 173[10])
    
endmodule
//
// Verilog Description of module Mixer
//

module Mixer (MixerOutCos, osc_clk, MixerOutSin, DiffOut_c, RFIn_c, 
            \LOCosine[2] , \LOCosine[3] , \LOCosine[6] , \LOCosine[7] , 
            \LOCosine[8] , \LOCosine[9] , \LOCosine[10] , \LOCosine[12] , 
            GND_net, \LOCosine[11] , \LOCosine[4] , \LOCosine[5] , \LOCosine[1] , 
            \LOSine[12] , \LOSine[10] , \LOSine[11] , \LOSine[8] , \LOSine[9] , 
            \LOSine[6] , \LOSine[7] , \LOSine[4] , \LOSine[5] , \LOSine[2] , 
            \LOSine[3] , \LOSine[1] ) /* synthesis syn_module_defined=1 */ ;
    output [11:0]MixerOutCos;
    input osc_clk;
    output [11:0]MixerOutSin;
    output DiffOut_c;
    input RFIn_c;
    input \LOCosine[2] ;
    input \LOCosine[3] ;
    input \LOCosine[6] ;
    input \LOCosine[7] ;
    input \LOCosine[8] ;
    input \LOCosine[9] ;
    input \LOCosine[10] ;
    input \LOCosine[12] ;
    input GND_net;
    input \LOCosine[11] ;
    input \LOCosine[4] ;
    input \LOCosine[5] ;
    input \LOCosine[1] ;
    input \LOSine[12] ;
    input \LOSine[10] ;
    input \LOSine[11] ;
    input \LOSine[8] ;
    input \LOSine[9] ;
    input \LOSine[6] ;
    input \LOSine[7] ;
    input \LOSine[4] ;
    input \LOSine[5] ;
    input \LOSine[2] ;
    input \LOSine[3] ;
    input \LOSine[1] ;
    
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(55[8:15])
    wire [11:0]MixerOutCos_11__N_223;
    wire [11:0]MixerOutSin_11__N_211;
    
    wire RFInR;
    wire [11:0]MixerOutCos_11__N_249;
    
    wire n11216, n11215, n11214, n11213, n11212, n11211, n11196;
    wire [11:0]MixerOutSin_11__N_235;
    
    wire n11195, n11194, n11193, n11192, n11191;
    
    FD1S3AX MixerOutCos_i4 (.D(MixerOutCos_11__N_223[4]), .CK(osc_clk), 
            .Q(MixerOutCos[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i4.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i3 (.D(MixerOutCos_11__N_223[3]), .CK(osc_clk), 
            .Q(MixerOutCos[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i3.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i0 (.D(MixerOutSin_11__N_211[0]), .CK(osc_clk), 
            .Q(MixerOutSin[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i0.GSR = "ENABLED";
    FD1S3AY RFInR_14 (.D(DiffOut_c), .CK(osc_clk), .Q(RFInR)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(23[10] 27[8])
    defparam RFInR_14.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i0 (.D(MixerOutCos_11__N_223[0]), .CK(osc_clk), 
            .Q(MixerOutCos[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i0.GSR = "ENABLED";
    FD1S3AY RFInR1_13 (.D(RFIn_c), .CK(osc_clk), .Q(DiffOut_c)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(23[10] 27[8])
    defparam RFInR1_13.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i2 (.D(MixerOutCos_11__N_223[2]), .CK(osc_clk), 
            .Q(MixerOutCos[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i2.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i1 (.D(MixerOutCos_11__N_223[1]), .CK(osc_clk), 
            .Q(MixerOutCos[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i1.GSR = "ENABLED";
    LUT4 MixerOutCos_11__I_0_i2_3_lut (.A(\LOCosine[2] ), .B(MixerOutCos_11__N_249[1]), 
         .C(RFInR), .Z(MixerOutCos_11__N_223[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i2_3_lut.init = 16'hcaca;
    FD1S3AX MixerOutSin_i7 (.D(MixerOutSin_11__N_211[7]), .CK(osc_clk), 
            .Q(MixerOutSin[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i7.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i6 (.D(MixerOutSin_11__N_211[6]), .CK(osc_clk), 
            .Q(MixerOutSin[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i6.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i5 (.D(MixerOutSin_11__N_211[5]), .CK(osc_clk), 
            .Q(MixerOutSin[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i5.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i4 (.D(MixerOutSin_11__N_211[4]), .CK(osc_clk), 
            .Q(MixerOutSin[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i4.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i3 (.D(MixerOutSin_11__N_211[3]), .CK(osc_clk), 
            .Q(MixerOutSin[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i3.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i2 (.D(MixerOutSin_11__N_211[2]), .CK(osc_clk), 
            .Q(MixerOutSin[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i2.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i1 (.D(MixerOutSin_11__N_211[1]), .CK(osc_clk), 
            .Q(MixerOutSin[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i1.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i8 (.D(MixerOutSin_11__N_211[8]), .CK(osc_clk), 
            .Q(MixerOutSin[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i8.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i9 (.D(MixerOutSin_11__N_211[9]), .CK(osc_clk), 
            .Q(MixerOutSin[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i9.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i10 (.D(MixerOutSin_11__N_211[10]), .CK(osc_clk), 
            .Q(MixerOutSin[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i10.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i11 (.D(MixerOutSin_11__N_211[11]), .CK(osc_clk), 
            .Q(MixerOutSin[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutSin_i11.GSR = "ENABLED";
    LUT4 MixerOutCos_11__I_0_i3_3_lut (.A(\LOCosine[3] ), .B(MixerOutCos_11__N_249[2]), 
         .C(RFInR), .Z(MixerOutCos_11__N_223[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i6_3_lut (.A(\LOCosine[6] ), .B(MixerOutCos_11__N_249[5]), 
         .C(RFInR), .Z(MixerOutCos_11__N_223[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i7_3_lut (.A(\LOCosine[7] ), .B(MixerOutCos_11__N_249[6]), 
         .C(RFInR), .Z(MixerOutCos_11__N_223[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i7_3_lut.init = 16'hcaca;
    FD1S3AX MixerOutCos_i5 (.D(MixerOutCos_11__N_223[5]), .CK(osc_clk), 
            .Q(MixerOutCos[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i5.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i6 (.D(MixerOutCos_11__N_223[6]), .CK(osc_clk), 
            .Q(MixerOutCos[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i6.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i7 (.D(MixerOutCos_11__N_223[7]), .CK(osc_clk), 
            .Q(MixerOutCos[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i7.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i8 (.D(MixerOutCos_11__N_223[8]), .CK(osc_clk), 
            .Q(MixerOutCos[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i8.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i9 (.D(MixerOutCos_11__N_223[9]), .CK(osc_clk), 
            .Q(MixerOutCos[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i9.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i10 (.D(MixerOutCos_11__N_223[10]), .CK(osc_clk), 
            .Q(MixerOutCos[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i10.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i11 (.D(MixerOutCos_11__N_223[11]), .CK(osc_clk), 
            .Q(MixerOutCos[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=2, LSE_LLINE=117, LSE_RLINE=125 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(32[10] 44[8])
    defparam MixerOutCos_i11.GSR = "ENABLED";
    LUT4 MixerOutCos_11__I_0_i8_3_lut (.A(\LOCosine[8] ), .B(MixerOutCos_11__N_249[7]), 
         .C(RFInR), .Z(MixerOutCos_11__N_223[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i9_3_lut (.A(\LOCosine[9] ), .B(MixerOutCos_11__N_249[8]), 
         .C(RFInR), .Z(MixerOutCos_11__N_223[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i10_3_lut (.A(\LOCosine[10] ), .B(MixerOutCos_11__N_249[9]), 
         .C(RFInR), .Z(MixerOutCos_11__N_223[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i10_3_lut.init = 16'hcaca;
    CCU2D unary_minus_7_add_3_13 (.A0(\LOCosine[12] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11216), .S0(MixerOutCos_11__N_249[11]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(42[26:33])
    defparam unary_minus_7_add_3_13.INIT0 = 16'hf555;
    defparam unary_minus_7_add_3_13.INIT1 = 16'h0000;
    defparam unary_minus_7_add_3_13.INJECT1_0 = "NO";
    defparam unary_minus_7_add_3_13.INJECT1_1 = "NO";
    CCU2D unary_minus_7_add_3_11 (.A0(\LOCosine[10] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOCosine[11] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11215), .COUT(n11216), .S0(MixerOutCos_11__N_249[9]), 
          .S1(MixerOutCos_11__N_249[10]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(42[26:33])
    defparam unary_minus_7_add_3_11.INIT0 = 16'hf555;
    defparam unary_minus_7_add_3_11.INIT1 = 16'hf555;
    defparam unary_minus_7_add_3_11.INJECT1_0 = "NO";
    defparam unary_minus_7_add_3_11.INJECT1_1 = "NO";
    CCU2D unary_minus_7_add_3_9 (.A0(\LOCosine[8] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOCosine[9] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11214), .COUT(n11215), .S0(MixerOutCos_11__N_249[7]), 
          .S1(MixerOutCos_11__N_249[8]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(42[26:33])
    defparam unary_minus_7_add_3_9.INIT0 = 16'hf555;
    defparam unary_minus_7_add_3_9.INIT1 = 16'hf555;
    defparam unary_minus_7_add_3_9.INJECT1_0 = "NO";
    defparam unary_minus_7_add_3_9.INJECT1_1 = "NO";
    CCU2D unary_minus_7_add_3_7 (.A0(\LOCosine[6] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOCosine[7] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11213), .COUT(n11214), .S0(MixerOutCos_11__N_249[5]), 
          .S1(MixerOutCos_11__N_249[6]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(42[26:33])
    defparam unary_minus_7_add_3_7.INIT0 = 16'hf555;
    defparam unary_minus_7_add_3_7.INIT1 = 16'hf555;
    defparam unary_minus_7_add_3_7.INJECT1_0 = "NO";
    defparam unary_minus_7_add_3_7.INJECT1_1 = "NO";
    CCU2D unary_minus_7_add_3_5 (.A0(\LOCosine[4] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOCosine[5] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11212), .COUT(n11213), .S0(MixerOutCos_11__N_249[3]), 
          .S1(MixerOutCos_11__N_249[4]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(42[26:33])
    defparam unary_minus_7_add_3_5.INIT0 = 16'hf555;
    defparam unary_minus_7_add_3_5.INIT1 = 16'hf555;
    defparam unary_minus_7_add_3_5.INJECT1_0 = "NO";
    defparam unary_minus_7_add_3_5.INJECT1_1 = "NO";
    CCU2D unary_minus_7_add_3_3 (.A0(\LOCosine[2] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOCosine[3] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11211), .COUT(n11212), .S0(MixerOutCos_11__N_249[1]), 
          .S1(MixerOutCos_11__N_249[2]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(42[26:33])
    defparam unary_minus_7_add_3_3.INIT0 = 16'hf555;
    defparam unary_minus_7_add_3_3.INIT1 = 16'hf555;
    defparam unary_minus_7_add_3_3.INJECT1_0 = "NO";
    defparam unary_minus_7_add_3_3.INJECT1_1 = "NO";
    CCU2D unary_minus_7_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOCosine[1] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n11211), .S1(MixerOutCos_11__N_249[0]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(42[26:33])
    defparam unary_minus_7_add_3_1.INIT0 = 16'hF000;
    defparam unary_minus_7_add_3_1.INIT1 = 16'h0aaa;
    defparam unary_minus_7_add_3_1.INJECT1_0 = "NO";
    defparam unary_minus_7_add_3_1.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_13 (.A0(\LOSine[12] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11196), .S0(MixerOutSin_11__N_235[11]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(41[26:33])
    defparam unary_minus_6_add_3_13.INIT0 = 16'hf555;
    defparam unary_minus_6_add_3_13.INIT1 = 16'h0000;
    defparam unary_minus_6_add_3_13.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_13.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_11 (.A0(\LOSine[10] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOSine[11] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11195), .COUT(n11196), .S0(MixerOutSin_11__N_235[9]), 
          .S1(MixerOutSin_11__N_235[10]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(41[26:33])
    defparam unary_minus_6_add_3_11.INIT0 = 16'hf555;
    defparam unary_minus_6_add_3_11.INIT1 = 16'hf555;
    defparam unary_minus_6_add_3_11.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_11.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_9 (.A0(\LOSine[8] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOSine[9] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11194), .COUT(n11195), .S0(MixerOutSin_11__N_235[7]), 
          .S1(MixerOutSin_11__N_235[8]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(41[26:33])
    defparam unary_minus_6_add_3_9.INIT0 = 16'hf555;
    defparam unary_minus_6_add_3_9.INIT1 = 16'hf555;
    defparam unary_minus_6_add_3_9.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_9.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_7 (.A0(\LOSine[6] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOSine[7] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11193), .COUT(n11194), .S0(MixerOutSin_11__N_235[5]), 
          .S1(MixerOutSin_11__N_235[6]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(41[26:33])
    defparam unary_minus_6_add_3_7.INIT0 = 16'hf555;
    defparam unary_minus_6_add_3_7.INIT1 = 16'hf555;
    defparam unary_minus_6_add_3_7.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_7.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_5 (.A0(\LOSine[4] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOSine[5] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11192), .COUT(n11193), .S0(MixerOutSin_11__N_235[3]), 
          .S1(MixerOutSin_11__N_235[4]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(41[26:33])
    defparam unary_minus_6_add_3_5.INIT0 = 16'hf555;
    defparam unary_minus_6_add_3_5.INIT1 = 16'hf555;
    defparam unary_minus_6_add_3_5.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_5.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_3 (.A0(\LOSine[2] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOSine[3] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11191), .COUT(n11192), .S0(MixerOutSin_11__N_235[1]), 
          .S1(MixerOutSin_11__N_235[2]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(41[26:33])
    defparam unary_minus_6_add_3_3.INIT0 = 16'hf555;
    defparam unary_minus_6_add_3_3.INIT1 = 16'hf555;
    defparam unary_minus_6_add_3_3.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_3.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\LOSine[1] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n11191), .S1(MixerOutSin_11__N_235[0]));   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(41[26:33])
    defparam unary_minus_6_add_3_1.INIT0 = 16'hF000;
    defparam unary_minus_6_add_3_1.INIT1 = 16'h0aaa;
    defparam unary_minus_6_add_3_1.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_1.INJECT1_1 = "NO";
    LUT4 MixerOutCos_11__I_0_i11_3_lut (.A(\LOCosine[11] ), .B(MixerOutCos_11__N_249[10]), 
         .C(RFInR), .Z(MixerOutCos_11__N_223[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i12_3_lut (.A(\LOCosine[12] ), .B(MixerOutCos_11__N_249[11]), 
         .C(RFInR), .Z(MixerOutCos_11__N_223[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i4_3_lut (.A(\LOCosine[4] ), .B(MixerOutCos_11__N_249[3]), 
         .C(RFInR), .Z(MixerOutCos_11__N_223[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i1_3_lut (.A(\LOSine[1] ), .B(MixerOutSin_11__N_235[0]), 
         .C(RFInR), .Z(MixerOutSin_11__N_211[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i1_3_lut (.A(\LOCosine[1] ), .B(MixerOutCos_11__N_249[0]), 
         .C(RFInR), .Z(MixerOutCos_11__N_223[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i8_3_lut (.A(\LOSine[8] ), .B(MixerOutSin_11__N_235[7]), 
         .C(RFInR), .Z(MixerOutSin_11__N_211[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i7_3_lut (.A(\LOSine[7] ), .B(MixerOutSin_11__N_235[6]), 
         .C(RFInR), .Z(MixerOutSin_11__N_211[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i6_3_lut (.A(\LOSine[6] ), .B(MixerOutSin_11__N_235[5]), 
         .C(RFInR), .Z(MixerOutSin_11__N_211[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i5_3_lut (.A(\LOSine[5] ), .B(MixerOutSin_11__N_235[4]), 
         .C(RFInR), .Z(MixerOutSin_11__N_211[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i4_3_lut (.A(\LOSine[4] ), .B(MixerOutSin_11__N_235[3]), 
         .C(RFInR), .Z(MixerOutSin_11__N_211[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i3_3_lut (.A(\LOSine[3] ), .B(MixerOutSin_11__N_235[2]), 
         .C(RFInR), .Z(MixerOutSin_11__N_211[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i5_3_lut (.A(\LOCosine[5] ), .B(MixerOutCos_11__N_249[4]), 
         .C(RFInR), .Z(MixerOutCos_11__N_223[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutCos_11__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i2_3_lut (.A(\LOSine[2] ), .B(MixerOutSin_11__N_235[1]), 
         .C(RFInR), .Z(MixerOutSin_11__N_211[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i9_3_lut (.A(\LOSine[9] ), .B(MixerOutSin_11__N_235[8]), 
         .C(RFInR), .Z(MixerOutSin_11__N_211[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i10_3_lut (.A(\LOSine[10] ), .B(MixerOutSin_11__N_235[9]), 
         .C(RFInR), .Z(MixerOutSin_11__N_211[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i11_3_lut (.A(\LOSine[11] ), .B(MixerOutSin_11__N_235[10]), 
         .C(RFInR), .Z(MixerOutSin_11__N_211[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i12_3_lut (.A(\LOSine[12] ), .B(MixerOutSin_11__N_235[11]), 
         .C(RFInR), .Z(MixerOutSin_11__N_211[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/mixer.v(40[9] 43[12])
    defparam MixerOutSin_11__I_0_i12_3_lut.init = 16'hcaca;
    
endmodule
//
// Verilog Description of module PWM
//

module PWM (osc_clk, \DataInReg_11__N_1855[0] , PWMOut_c, \DataInReg_11__N_1855[1] , 
            \DataInReg_11__N_1855[2] , \DataInReg_11__N_1855[3] , \DataInReg_11__N_1855[4] , 
            \DataInReg_11__N_1855[5] , \DataInReg_11__N_1855[6] , \DataInReg_11__N_1855[7] , 
            \DataInReg_11__N_1855[8] , GND_net, \DemodOut[9] ) /* synthesis syn_module_defined=1 */ ;
    input osc_clk;
    input \DataInReg_11__N_1855[0] ;
    output PWMOut_c;
    input \DataInReg_11__N_1855[1] ;
    input \DataInReg_11__N_1855[2] ;
    input \DataInReg_11__N_1855[3] ;
    input \DataInReg_11__N_1855[4] ;
    input \DataInReg_11__N_1855[5] ;
    input \DataInReg_11__N_1855[6] ;
    input \DataInReg_11__N_1855[7] ;
    input \DataInReg_11__N_1855[8] ;
    input GND_net;
    input \DemodOut[9] ;
    
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(55[8:15])
    wire [11:0]DataInReg;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(10[12:21])
    
    wire osc_clk_enable_1392, PWMOut_N_1868;
    wire [9:0]counter;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(7[11:18])
    wire [9:0]n45;
    
    wire n15;
    wire [11:0]n3822;
    
    wire n11, n17, n12, n11114, n11113, n11112, n11111, n11110, 
        n11616, n11615, n11614, n11613, n11612;
    
    FD1P3AX DataInReg__i1 (.D(\DataInReg_11__N_1855[0] ), .SP(osc_clk_enable_1392), 
            .CK(osc_clk), .Q(DataInReg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=146, LSE_RLINE=152 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i1.GSR = "ENABLED";
    FD1S3AX PWMOut_15 (.D(PWMOut_N_1868), .CK(osc_clk), .Q(PWMOut_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=146, LSE_RLINE=152 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam PWMOut_15.GSR = "ENABLED";
    FD1S3AX counter_929__i0 (.D(n45[0]), .CK(osc_clk), .Q(counter[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_929__i0.GSR = "ENABLED";
    LUT4 i5_2_lut (.A(counter[2]), .B(counter[9]), .Z(n15)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(26[7:19])
    defparam i5_2_lut.init = 16'heeee;
    FD1P3AX DataInReg__i2 (.D(\DataInReg_11__N_1855[1] ), .SP(osc_clk_enable_1392), 
            .CK(osc_clk), .Q(DataInReg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=146, LSE_RLINE=152 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i2.GSR = "ENABLED";
    FD1P3AX DataInReg__i3 (.D(\DataInReg_11__N_1855[2] ), .SP(osc_clk_enable_1392), 
            .CK(osc_clk), .Q(DataInReg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=146, LSE_RLINE=152 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i3.GSR = "ENABLED";
    FD1P3AX DataInReg__i4 (.D(\DataInReg_11__N_1855[3] ), .SP(osc_clk_enable_1392), 
            .CK(osc_clk), .Q(DataInReg[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=146, LSE_RLINE=152 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i4.GSR = "ENABLED";
    FD1P3AX DataInReg__i5 (.D(\DataInReg_11__N_1855[4] ), .SP(osc_clk_enable_1392), 
            .CK(osc_clk), .Q(DataInReg[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=146, LSE_RLINE=152 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i5.GSR = "ENABLED";
    FD1P3AX DataInReg__i6 (.D(\DataInReg_11__N_1855[5] ), .SP(osc_clk_enable_1392), 
            .CK(osc_clk), .Q(DataInReg[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=146, LSE_RLINE=152 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i6.GSR = "ENABLED";
    FD1P3AX DataInReg__i7 (.D(\DataInReg_11__N_1855[6] ), .SP(osc_clk_enable_1392), 
            .CK(osc_clk), .Q(DataInReg[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=146, LSE_RLINE=152 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i7.GSR = "ENABLED";
    FD1P3AX DataInReg__i8 (.D(\DataInReg_11__N_1855[7] ), .SP(osc_clk_enable_1392), 
            .CK(osc_clk), .Q(DataInReg[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=146, LSE_RLINE=152 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i8.GSR = "ENABLED";
    FD1P3AX DataInReg__i9 (.D(\DataInReg_11__N_1855[8] ), .SP(osc_clk_enable_1392), 
            .CK(osc_clk), .Q(DataInReg[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=146, LSE_RLINE=152 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i9.GSR = "ENABLED";
    FD1P3AX DataInReg__i10 (.D(n3822[9]), .SP(osc_clk_enable_1392), .CK(osc_clk), 
            .Q(DataInReg[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=146, LSE_RLINE=152 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(23[8] 35[5])
    defparam DataInReg__i10.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(counter[0]), .B(counter[5]), .Z(n11)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(26[7:19])
    defparam i1_2_lut.init = 16'heeee;
    FD1S3AX counter_929__i1 (.D(n45[1]), .CK(osc_clk), .Q(counter[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_929__i1.GSR = "ENABLED";
    FD1S3AX counter_929__i2 (.D(n45[2]), .CK(osc_clk), .Q(counter[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_929__i2.GSR = "ENABLED";
    FD1S3AX counter_929__i3 (.D(n45[3]), .CK(osc_clk), .Q(counter[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_929__i3.GSR = "ENABLED";
    FD1S3AX counter_929__i4 (.D(n45[4]), .CK(osc_clk), .Q(counter[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_929__i4.GSR = "ENABLED";
    FD1S3AX counter_929__i5 (.D(n45[5]), .CK(osc_clk), .Q(counter[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_929__i5.GSR = "ENABLED";
    FD1S3AX counter_929__i6 (.D(n45[6]), .CK(osc_clk), .Q(counter[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_929__i6.GSR = "ENABLED";
    FD1S3AX counter_929__i7 (.D(n45[7]), .CK(osc_clk), .Q(counter[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_929__i7.GSR = "ENABLED";
    FD1S3AX counter_929__i8 (.D(n45[8]), .CK(osc_clk), .Q(counter[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_929__i8.GSR = "ENABLED";
    FD1S3AX counter_929__i9 (.D(n45[9]), .CK(osc_clk), .Q(counter[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_929__i9.GSR = "ENABLED";
    LUT4 i5915_4_lut (.A(n17), .B(n15), .C(n11), .D(n12), .Z(osc_clk_enable_1392)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(26[7:19])
    defparam i5915_4_lut.init = 16'h0001;
    LUT4 i7_4_lut (.A(counter[4]), .B(counter[1]), .C(counter[6]), .D(counter[8]), 
         .Z(n17)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(26[7:19])
    defparam i7_4_lut.init = 16'hfffe;
    CCU2D sub_718_add_2_11 (.A0(DataInReg[9]), .B0(counter[9]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11114), .S1(PWMOut_N_1868));
    defparam sub_718_add_2_11.INIT0 = 16'h5999;
    defparam sub_718_add_2_11.INIT1 = 16'h0000;
    defparam sub_718_add_2_11.INJECT1_0 = "NO";
    defparam sub_718_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_718_add_2_9 (.A0(DataInReg[7]), .B0(counter[7]), .C0(GND_net), 
          .D0(GND_net), .A1(DataInReg[8]), .B1(counter[8]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11113), .COUT(n11114));
    defparam sub_718_add_2_9.INIT0 = 16'h5999;
    defparam sub_718_add_2_9.INIT1 = 16'h5999;
    defparam sub_718_add_2_9.INJECT1_0 = "NO";
    defparam sub_718_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_718_add_2_7 (.A0(DataInReg[5]), .B0(counter[5]), .C0(GND_net), 
          .D0(GND_net), .A1(DataInReg[6]), .B1(counter[6]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11112), .COUT(n11113));
    defparam sub_718_add_2_7.INIT0 = 16'h5999;
    defparam sub_718_add_2_7.INIT1 = 16'h5999;
    defparam sub_718_add_2_7.INJECT1_0 = "NO";
    defparam sub_718_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_718_add_2_5 (.A0(DataInReg[3]), .B0(counter[3]), .C0(GND_net), 
          .D0(GND_net), .A1(DataInReg[4]), .B1(counter[4]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11111), .COUT(n11112));
    defparam sub_718_add_2_5.INIT0 = 16'h5999;
    defparam sub_718_add_2_5.INIT1 = 16'h5999;
    defparam sub_718_add_2_5.INJECT1_0 = "NO";
    defparam sub_718_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_718_add_2_3 (.A0(DataInReg[1]), .B0(counter[1]), .C0(GND_net), 
          .D0(GND_net), .A1(DataInReg[2]), .B1(counter[2]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11110), .COUT(n11111));
    defparam sub_718_add_2_3.INIT0 = 16'h5999;
    defparam sub_718_add_2_3.INIT1 = 16'h5999;
    defparam sub_718_add_2_3.INJECT1_0 = "NO";
    defparam sub_718_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_718_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(DataInReg[0]), .B1(counter[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n11110));
    defparam sub_718_add_2_1.INIT0 = 16'h0000;
    defparam sub_718_add_2_1.INIT1 = 16'h5999;
    defparam sub_718_add_2_1.INJECT1_0 = "NO";
    defparam sub_718_add_2_1.INJECT1_1 = "NO";
    CCU2D counter_929_add_4_11 (.A0(counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11616), .S0(n45[9]));   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_929_add_4_11.INIT0 = 16'hfaaa;
    defparam counter_929_add_4_11.INIT1 = 16'h0000;
    defparam counter_929_add_4_11.INJECT1_0 = "NO";
    defparam counter_929_add_4_11.INJECT1_1 = "NO";
    CCU2D counter_929_add_4_9 (.A0(counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11615), .COUT(n11616), .S0(n45[7]), .S1(n45[8]));   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_929_add_4_9.INIT0 = 16'hfaaa;
    defparam counter_929_add_4_9.INIT1 = 16'hfaaa;
    defparam counter_929_add_4_9.INJECT1_0 = "NO";
    defparam counter_929_add_4_9.INJECT1_1 = "NO";
    CCU2D counter_929_add_4_7 (.A0(counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11614), .COUT(n11615), .S0(n45[5]), .S1(n45[6]));   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_929_add_4_7.INIT0 = 16'hfaaa;
    defparam counter_929_add_4_7.INIT1 = 16'hfaaa;
    defparam counter_929_add_4_7.INJECT1_0 = "NO";
    defparam counter_929_add_4_7.INJECT1_1 = "NO";
    CCU2D counter_929_add_4_5 (.A0(counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11613), .COUT(n11614), .S0(n45[3]), .S1(n45[4]));   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_929_add_4_5.INIT0 = 16'hfaaa;
    defparam counter_929_add_4_5.INIT1 = 16'hfaaa;
    defparam counter_929_add_4_5.INJECT1_0 = "NO";
    defparam counter_929_add_4_5.INJECT1_1 = "NO";
    CCU2D counter_929_add_4_3 (.A0(counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11612), .COUT(n11613), .S0(n45[1]), .S1(n45[2]));   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_929_add_4_3.INIT0 = 16'hfaaa;
    defparam counter_929_add_4_3.INIT1 = 16'hfaaa;
    defparam counter_929_add_4_3.INJECT1_0 = "NO";
    defparam counter_929_add_4_3.INJECT1_1 = "NO";
    CCU2D counter_929_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n11612), .S1(n45[0]));   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(25[14:29])
    defparam counter_929_add_4_1.INIT0 = 16'hF000;
    defparam counter_929_add_4_1.INIT1 = 16'h0555;
    defparam counter_929_add_4_1.INJECT1_0 = "NO";
    defparam counter_929_add_4_1.INJECT1_1 = "NO";
    LUT4 i2_2_lut (.A(counter[7]), .B(counter[3]), .Z(n12)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(26[7:19])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i1091_1_lut (.A(\DemodOut[9] ), .Z(n3822[9])) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/pwm.v(26[3] 27[35])
    defparam i1091_1_lut.init = 16'h5555;
    
endmodule
//
// Verilog Description of module \uart_tx(CLKS_PER_BIT=87) 
//

module \uart_tx(CLKS_PER_BIT=87)  (\UartClk[2] , o_Rx_Byte_c_0, n12872, 
            n7319, o_Rx_Byte_c_4, n2215, o_Tx_Serial_c, o_Rx_DV_c_0, 
            o_Rx_Byte_c_7, o_Rx_Byte_c_2, osc_clk, o_Rx_Byte_c_6, o_Rx_Byte_c_5, 
            o_Rx_Byte_c_3, GND_net, n13765, n13753, n13151) /* synthesis syn_module_defined=1 */ ;
    output \UartClk[2] ;
    input o_Rx_Byte_c_0;
    output n12872;
    input n7319;
    input o_Rx_Byte_c_4;
    output n2215;
    output o_Tx_Serial_c;
    input o_Rx_DV_c_0;
    input o_Rx_Byte_c_7;
    input o_Rx_Byte_c_2;
    input osc_clk;
    input o_Rx_Byte_c_6;
    input o_Rx_Byte_c_5;
    input o_Rx_Byte_c_3;
    input GND_net;
    input n13765;
    output n13753;
    output n13151;
    
    wire \UartClk[2]  /* synthesis SET_AS_NETWORK=\uart_tx1/UartClk[2], is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(37[14:21])
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(55[8:15])
    wire [7:0]r_Tx_Data;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(34[16:25])
    wire [2:0]r_Bit_Index;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(33[16:27])
    
    wire n13261, n13262, n13263, UartClk_2_enable_5, n3, n13046;
    wire [2:0]r_SM_Main;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(31[16:25])
    
    wire n13013;
    wire [2:0]r_SM_Main_2__N_2530;
    
    wire n7667, n3_adj_2612;
    wire [15:0]n121;
    
    wire UartClk_2_enable_41, n8364;
    wire [15:0]n69;
    
    wire n39, UartClk_2_enable_40, n13147;
    wire [2:0]n30;
    wire [2:0]n17;
    
    wire n13260, n9244, n13258, n13259;
    wire [15:0]r_Clock_Count;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(32[17:30])
    
    wire n12242, n12241, n12240, n12239, n3_adj_2614, n12238, n12237, 
        n12236, n12235, n13755, n3_adj_2615, n13766, n11625, n7, 
        n50, n6, n8994, n13031;
    
    LUT4 i5812_3_lut (.A(r_Tx_Data[2]), .B(r_Tx_Data[3]), .C(r_Bit_Index[0]), 
         .Z(n13261)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5812_3_lut.init = 16'hcaca;
    PFUMX i5814 (.BLUT(n13261), .ALUT(n13262), .C0(r_Bit_Index[2]), .Z(n13263));
    FD1P3AX r_Bit_Index_i2 (.D(n3), .SP(UartClk_2_enable_5), .CK(\UartClk[2] ), 
            .Q(r_Bit_Index[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=184, LSE_RLINE=191 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(45[10] 148[8])
    defparam r_Bit_Index_i2.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(o_Rx_Byte_c_0), .B(n12872), .C(n7319), .D(o_Rx_Byte_c_4), 
         .Z(n2215)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(48[7] 147[14])
    defparam i1_4_lut.init = 16'h4000;
    FD1P3AX r_Bit_Index_i1 (.D(n13046), .SP(UartClk_2_enable_5), .CK(\UartClk[2] ), 
            .Q(r_Bit_Index[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=184, LSE_RLINE=191 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(45[10] 148[8])
    defparam r_Bit_Index_i1.GSR = "ENABLED";
    FD1S3IX r_SM_Main_i2 (.D(r_SM_Main_2__N_2530[1]), .CK(\UartClk[2] ), 
            .CD(n13013), .Q(r_SM_Main[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=184, LSE_RLINE=191 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(45[10] 148[8])
    defparam r_SM_Main_i2.GSR = "ENABLED";
    FD1S3IX r_SM_Main_i0 (.D(n7667), .CK(\UartClk[2] ), .CD(r_SM_Main[2]), 
            .Q(r_SM_Main[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=184, LSE_RLINE=191 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(45[10] 148[8])
    defparam r_SM_Main_i0.GSR = "ENABLED";
    FD1P3AX r_Bit_Index_i0 (.D(n3_adj_2612), .SP(UartClk_2_enable_5), .CK(\UartClk[2] ), 
            .Q(r_Bit_Index[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=184, LSE_RLINE=191 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(45[10] 148[8])
    defparam r_Bit_Index_i0.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_935__i0 (.D(n69[0]), .SP(UartClk_2_enable_41), 
            .CD(n8364), .CK(\UartClk[2] ), .Q(n121[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935__i0.GSR = "ENABLED";
    FD1P3AX o_Tx_Serial_47 (.D(n39), .SP(UartClk_2_enable_41), .CK(\UartClk[2] ), 
            .Q(o_Tx_Serial_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=184, LSE_RLINE=191 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(45[10] 148[8])
    defparam o_Tx_Serial_47.GSR = "ENABLED";
    FD1P3AX r_Tx_Data_i0 (.D(o_Rx_Byte_c_0), .SP(UartClk_2_enable_40), .CK(\UartClk[2] ), 
            .Q(r_Tx_Data[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=184, LSE_RLINE=191 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(45[10] 148[8])
    defparam r_Tx_Data_i0.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_55 (.A(n13147), .B(o_Rx_DV_c_0), .C(o_Rx_Byte_c_7), 
         .D(o_Rx_Byte_c_2), .Z(n12872)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_55.init = 16'h0008;
    FD1S3AX UartClk_933_965__i0 (.D(n17[0]), .CK(osc_clk), .Q(n30[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(42[15:29])
    defparam UartClk_933_965__i0.GSR = "ENABLED";
    L6MUX21 i3242 (.D0(n13260), .D1(n13263), .SD(r_Bit_Index[1]), .Z(n9244));
    PFUMX i5811 (.BLUT(n13258), .ALUT(n13259), .C0(r_Bit_Index[0]), .Z(n13260));
    LUT4 i1_1_lut_rep_180 (.A(r_SM_Main[2]), .Z(UartClk_2_enable_41)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1_1_lut_rep_180.init = 16'h5555;
    LUT4 i2361_4_lut_4_lut (.A(r_SM_Main[2]), .B(r_SM_Main[0]), .C(r_SM_Main[1]), 
         .D(r_SM_Main_2__N_2530[1]), .Z(n8364)) /* synthesis lut_function=(!(A+!(B (D)+!B ((D)+!C)))) */ ;
    defparam i2361_4_lut_4_lut.init = 16'h5501;
    LUT4 i5899_3_lut (.A(r_SM_Main[2]), .B(r_SM_Main[1]), .C(r_SM_Main[0]), 
         .Z(n13013)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i5899_3_lut.init = 16'hbfbf;
    LUT4 i1_3_lut (.A(o_Rx_Byte_c_6), .B(o_Rx_Byte_c_5), .C(o_Rx_Byte_c_3), 
         .Z(n13147)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_3_lut.init = 16'h0808;
    FD1P3IX r_Clock_Count_935__i15 (.D(n69[15]), .SP(UartClk_2_enable_41), 
            .CD(n8364), .CK(\UartClk[2] ), .Q(r_Clock_Count[15])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935__i15.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_935__i14 (.D(n69[14]), .SP(UartClk_2_enable_41), 
            .CD(n8364), .CK(\UartClk[2] ), .Q(r_Clock_Count[14])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935__i14.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_935__i13 (.D(n69[13]), .SP(UartClk_2_enable_41), 
            .CD(n8364), .CK(\UartClk[2] ), .Q(r_Clock_Count[13])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935__i13.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_935__i12 (.D(n69[12]), .SP(UartClk_2_enable_41), 
            .CD(n8364), .CK(\UartClk[2] ), .Q(r_Clock_Count[12])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935__i12.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_935__i11 (.D(n69[11]), .SP(UartClk_2_enable_41), 
            .CD(n8364), .CK(\UartClk[2] ), .Q(r_Clock_Count[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935__i11.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_935__i10 (.D(n69[10]), .SP(UartClk_2_enable_41), 
            .CD(n8364), .CK(\UartClk[2] ), .Q(r_Clock_Count[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935__i10.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_935__i9 (.D(n69[9]), .SP(UartClk_2_enable_41), 
            .CD(n8364), .CK(\UartClk[2] ), .Q(r_Clock_Count[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935__i9.GSR = "ENABLED";
    CCU2D r_Clock_Count_935_add_4_17 (.A0(r_Clock_Count[15]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12242), .S0(n69[15]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935_add_4_17.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_935_add_4_17.INIT1 = 16'h0000;
    defparam r_Clock_Count_935_add_4_17.INJECT1_0 = "NO";
    defparam r_Clock_Count_935_add_4_17.INJECT1_1 = "NO";
    FD1P3IX r_Clock_Count_935__i8 (.D(n69[8]), .SP(UartClk_2_enable_41), 
            .CD(n8364), .CK(\UartClk[2] ), .Q(r_Clock_Count[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935__i8.GSR = "ENABLED";
    CCU2D r_Clock_Count_935_add_4_15 (.A0(r_Clock_Count[13]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[14]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12241), .COUT(n12242), .S0(n69[13]), 
          .S1(n69[14]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935_add_4_15.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_935_add_4_15.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_935_add_4_15.INJECT1_0 = "NO";
    defparam r_Clock_Count_935_add_4_15.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_935_add_4_13 (.A0(r_Clock_Count[11]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[12]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12240), .COUT(n12241), .S0(n69[11]), 
          .S1(n69[12]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935_add_4_13.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_935_add_4_13.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_935_add_4_13.INJECT1_0 = "NO";
    defparam r_Clock_Count_935_add_4_13.INJECT1_1 = "NO";
    FD1P3IX r_Clock_Count_935__i7 (.D(n69[7]), .SP(UartClk_2_enable_41), 
            .CD(n8364), .CK(\UartClk[2] ), .Q(r_Clock_Count[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935__i7.GSR = "ENABLED";
    CCU2D r_Clock_Count_935_add_4_11 (.A0(r_Clock_Count[9]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[10]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12239), .COUT(n12240), .S0(n69[9]), 
          .S1(n69[10]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935_add_4_11.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_935_add_4_11.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_935_add_4_11.INJECT1_0 = "NO";
    defparam r_Clock_Count_935_add_4_11.INJECT1_1 = "NO";
    FD1P3IX r_Clock_Count_935__i6 (.D(n69[6]), .SP(UartClk_2_enable_41), 
            .CD(n8364), .CK(\UartClk[2] ), .Q(r_Clock_Count[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935__i6.GSR = "ENABLED";
    FD1S3IX r_SM_Main_i1 (.D(n3_adj_2614), .CK(\UartClk[2] ), .CD(r_SM_Main[2]), 
            .Q(r_SM_Main[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=184, LSE_RLINE=191 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(45[10] 148[8])
    defparam r_SM_Main_i1.GSR = "ENABLED";
    CCU2D r_Clock_Count_935_add_4_9 (.A0(r_Clock_Count[7]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[8]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12238), .COUT(n12239), .S0(n69[7]), 
          .S1(n69[8]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935_add_4_9.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_935_add_4_9.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_935_add_4_9.INJECT1_0 = "NO";
    defparam r_Clock_Count_935_add_4_9.INJECT1_1 = "NO";
    FD1P3IX r_Clock_Count_935__i5 (.D(n69[5]), .SP(UartClk_2_enable_41), 
            .CD(n8364), .CK(\UartClk[2] ), .Q(r_Clock_Count[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935__i5.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_935__i4 (.D(n69[4]), .SP(UartClk_2_enable_41), 
            .CD(n8364), .CK(\UartClk[2] ), .Q(r_Clock_Count[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935__i4.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_935__i3 (.D(n69[3]), .SP(UartClk_2_enable_41), 
            .CD(n8364), .CK(\UartClk[2] ), .Q(r_Clock_Count[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935__i3.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_935__i2 (.D(n69[2]), .SP(UartClk_2_enable_41), 
            .CD(n8364), .CK(\UartClk[2] ), .Q(r_Clock_Count[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935__i2.GSR = "ENABLED";
    CCU2D r_Clock_Count_935_add_4_7 (.A0(r_Clock_Count[5]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[6]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12237), .COUT(n12238), .S0(n69[5]), 
          .S1(n69[6]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935_add_4_7.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_935_add_4_7.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_935_add_4_7.INJECT1_0 = "NO";
    defparam r_Clock_Count_935_add_4_7.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_935_add_4_5 (.A0(r_Clock_Count[3]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[4]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12236), .COUT(n12237), .S0(n69[3]), 
          .S1(n69[4]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935_add_4_5.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_935_add_4_5.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_935_add_4_5.INJECT1_0 = "NO";
    defparam r_Clock_Count_935_add_4_5.INJECT1_1 = "NO";
    FD1P3AX r_Tx_Data_i1 (.D(n7319), .SP(UartClk_2_enable_40), .CK(\UartClk[2] ), 
            .Q(r_Tx_Data[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=184, LSE_RLINE=191 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(45[10] 148[8])
    defparam r_Tx_Data_i1.GSR = "ENABLED";
    FD1P3AX r_Tx_Data_i2 (.D(o_Rx_Byte_c_2), .SP(UartClk_2_enable_40), .CK(\UartClk[2] ), 
            .Q(r_Tx_Data[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=184, LSE_RLINE=191 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(45[10] 148[8])
    defparam r_Tx_Data_i2.GSR = "ENABLED";
    FD1P3AX r_Tx_Data_i3 (.D(o_Rx_Byte_c_3), .SP(UartClk_2_enable_40), .CK(\UartClk[2] ), 
            .Q(r_Tx_Data[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=184, LSE_RLINE=191 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(45[10] 148[8])
    defparam r_Tx_Data_i3.GSR = "ENABLED";
    FD1P3AX r_Tx_Data_i4 (.D(o_Rx_Byte_c_4), .SP(UartClk_2_enable_40), .CK(\UartClk[2] ), 
            .Q(r_Tx_Data[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=184, LSE_RLINE=191 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(45[10] 148[8])
    defparam r_Tx_Data_i4.GSR = "ENABLED";
    FD1P3AX r_Tx_Data_i5 (.D(o_Rx_Byte_c_5), .SP(UartClk_2_enable_40), .CK(\UartClk[2] ), 
            .Q(r_Tx_Data[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=184, LSE_RLINE=191 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(45[10] 148[8])
    defparam r_Tx_Data_i5.GSR = "ENABLED";
    FD1P3AX r_Tx_Data_i6 (.D(o_Rx_Byte_c_6), .SP(UartClk_2_enable_40), .CK(\UartClk[2] ), 
            .Q(r_Tx_Data[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=184, LSE_RLINE=191 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(45[10] 148[8])
    defparam r_Tx_Data_i6.GSR = "ENABLED";
    FD1P3AX r_Tx_Data_i7 (.D(o_Rx_Byte_c_7), .SP(UartClk_2_enable_40), .CK(\UartClk[2] ), 
            .Q(r_Tx_Data[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=184, LSE_RLINE=191 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(45[10] 148[8])
    defparam r_Tx_Data_i7.GSR = "ENABLED";
    CCU2D r_Clock_Count_935_add_4_3 (.A0(r_Clock_Count[1]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[2]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12235), .COUT(n12236), .S0(n69[1]), 
          .S1(n69[2]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935_add_4_3.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_935_add_4_3.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_935_add_4_3.INJECT1_0 = "NO";
    defparam r_Clock_Count_935_add_4_3.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_935_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n121[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n12235), .S1(n69[0]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935_add_4_1.INIT0 = 16'hF000;
    defparam r_Clock_Count_935_add_4_1.INIT1 = 16'h0555;
    defparam r_Clock_Count_935_add_4_1.INJECT1_0 = "NO";
    defparam r_Clock_Count_935_add_4_1.INJECT1_1 = "NO";
    LUT4 i1_3_lut_rep_162 (.A(r_SM_Main[0]), .B(r_SM_Main_2__N_2530[1]), 
         .C(r_SM_Main[1]), .Z(n13755)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(45[10] 148[8])
    defparam i1_3_lut_rep_162.init = 16'h4040;
    LUT4 i1_2_lut_4_lut (.A(r_SM_Main[0]), .B(r_SM_Main_2__N_2530[1]), .C(r_SM_Main[1]), 
         .D(r_Bit_Index[0]), .Z(n3_adj_2612)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(45[10] 148[8])
    defparam i1_2_lut_4_lut.init = 16'h0040;
    LUT4 i1679_2_lut_rep_160_4_lut (.A(n13765), .B(n12872), .C(o_Rx_Byte_c_0), 
         .D(o_Rx_Byte_c_3), .Z(n13753)) /* synthesis lut_function=(A (D)+!A !(B (C+!(D))+!B !(D))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(48[7] 147[14])
    defparam i1679_2_lut_rep_160_4_lut.init = 16'hbf00;
    LUT4 i1_2_lut_4_lut_adj_56 (.A(n13765), .B(n12872), .C(o_Rx_Byte_c_0), 
         .D(o_Rx_Byte_c_2), .Z(n13151)) /* synthesis lut_function=(A (D)+!A !(B (C+!(D))+!B !(D))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(48[7] 147[14])
    defparam i1_2_lut_4_lut_adj_56.init = 16'hbf00;
    LUT4 i5809_3_lut (.A(r_Tx_Data[0]), .B(r_Tx_Data[4]), .C(r_Bit_Index[2]), 
         .Z(n13258)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5809_3_lut.init = 16'hcaca;
    LUT4 i7_3_lut (.A(n3_adj_2615), .B(r_SM_Main_2__N_2530[1]), .C(r_SM_Main[0]), 
         .Z(n7667)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(31[16:25])
    defparam i7_3_lut.init = 16'h3a3a;
    FD1S3AX UartClk_933_965__i1 (.D(n17[1]), .CK(osc_clk), .Q(n30[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(42[15:29])
    defparam UartClk_933_965__i1.GSR = "ENABLED";
    FD1S3AX UartClk_933_965__i2 (.D(n17[2]), .CK(osc_clk), .Q(\UartClk[2] )) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(42[15:29])
    defparam UartClk_933_965__i2.GSR = "ENABLED";
    LUT4 i6_4_lut (.A(o_Rx_DV_c_0), .B(n13766), .C(r_SM_Main[1]), .D(r_SM_Main_2__N_2530[1]), 
         .Z(n3_adj_2615)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(31[16:25])
    defparam i6_4_lut.init = 16'hca0a;
    CCU2D UartClk_933_965_add_4_3 (.A0(n30[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\UartClk[2] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11625), .S0(n17[1]), .S1(n17[2]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(42[15:29])
    defparam UartClk_933_965_add_4_3.INIT0 = 16'hfaaa;
    defparam UartClk_933_965_add_4_3.INIT1 = 16'hfaaa;
    defparam UartClk_933_965_add_4_3.INJECT1_0 = "NO";
    defparam UartClk_933_965_add_4_3.INJECT1_1 = "NO";
    CCU2D UartClk_933_965_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n30[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n11625), .S1(n17[0]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(42[15:29])
    defparam UartClk_933_965_add_4_1.INIT0 = 16'hF000;
    defparam UartClk_933_965_add_4_1.INIT1 = 16'h0555;
    defparam UartClk_933_965_add_4_1.INJECT1_0 = "NO";
    defparam UartClk_933_965_add_4_1.INJECT1_1 = "NO";
    LUT4 i20_3_lut (.A(r_SM_Main[0]), .B(r_SM_Main[1]), .C(r_SM_Main_2__N_2530[1]), 
         .Z(n3_adj_2614)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(31[16:25])
    defparam i20_3_lut.init = 16'h6c6c;
    LUT4 i5813_3_lut (.A(r_Tx_Data[6]), .B(r_Tx_Data[7]), .C(r_Bit_Index[0]), 
         .Z(n13262)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5813_3_lut.init = 16'hcaca;
    LUT4 i5810_3_lut (.A(r_Tx_Data[1]), .B(r_Tx_Data[5]), .C(r_Bit_Index[2]), 
         .Z(n13259)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5810_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_57 (.A(n13755), .B(r_Bit_Index[2]), .C(r_Bit_Index[1]), 
         .D(r_Bit_Index[0]), .Z(n3)) /* synthesis lut_function=(!((B (C (D))+!B !(C (D)))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(45[10] 148[8])
    defparam i1_4_lut_adj_57.init = 16'h2888;
    LUT4 i3244_3_lut (.A(r_SM_Main[0]), .B(n9244), .C(r_SM_Main[1]), .Z(n39)) /* synthesis lut_function=(A (C)+!A (B+!(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(31[16:25])
    defparam i3244_3_lut.init = 16'he5e5;
    FD1P3IX r_Clock_Count_935__i1 (.D(n69[1]), .SP(UartClk_2_enable_41), 
            .CD(n8364), .CK(\UartClk[2] ), .Q(r_Clock_Count[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam r_Clock_Count_935__i1.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_173 (.A(r_Bit_Index[0]), .B(r_Bit_Index[2]), .C(r_Bit_Index[1]), 
         .Z(n13766)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut_rep_173.init = 16'h8080;
    LUT4 i1_4_lut_3_lut (.A(r_Bit_Index[0]), .B(r_Bit_Index[1]), .C(n13755), 
         .Z(n13046)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;
    defparam i1_4_lut_3_lut.init = 16'h6060;
    LUT4 i1_4_lut_adj_58 (.A(n7), .B(n50), .C(r_Clock_Count[11]), .D(n6), 
         .Z(r_SM_Main_2__N_2530[1])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam i1_4_lut_adj_58.init = 16'hfffe;
    LUT4 i2_2_lut (.A(r_Clock_Count[9]), .B(r_Clock_Count[15]), .Z(n7)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i72_4_lut (.A(r_Clock_Count[5]), .B(r_Clock_Count[6]), .C(n8994), 
         .D(r_Clock_Count[4]), .Z(n50)) /* synthesis lut_function=(A (B)+!A (B (C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(32[17:30])
    defparam i72_4_lut.init = 16'hc888;
    LUT4 i1_3_lut_4_lut (.A(r_SM_Main[0]), .B(r_SM_Main[2]), .C(r_SM_Main_2__N_2530[1]), 
         .D(r_SM_Main[1]), .Z(UartClk_2_enable_5)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h1011;
    LUT4 i2_3_lut_4_lut (.A(r_SM_Main[0]), .B(r_SM_Main[2]), .C(o_Rx_DV_c_0), 
         .D(r_SM_Main[1]), .Z(UartClk_2_enable_40)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_4_lut_adj_59 (.A(r_Clock_Count[7]), .B(r_Clock_Count[8]), .C(r_Clock_Count[13]), 
         .D(n13031), .Z(n6)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam i1_4_lut_adj_59.init = 16'hfffe;
    LUT4 i2991_3_lut (.A(r_Clock_Count[1]), .B(r_Clock_Count[3]), .C(r_Clock_Count[2]), 
         .Z(n8994)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i2991_3_lut.init = 16'hecec;
    LUT4 i2_3_lut (.A(r_Clock_Count[12]), .B(r_Clock_Count[14]), .C(r_Clock_Count[10]), 
         .Z(n13031)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(123[34:54])
    defparam i2_3_lut.init = 16'hfefe;
    
endmodule
//
// Verilog Description of module SinCos
//

module SinCos (osc_clk, VCC_net, GND_net, \phase_accum[57] , \phase_accum[58] , 
            \phase_accum[59] , \phase_accum[60] , \phase_accum[61] , \phase_accum[62] , 
            \phase_accum[63] , \LOSine[1] , \LOSine[2] , \LOSine[3] , 
            \LOSine[4] , \LOSine[5] , \LOSine[6] , \LOSine[7] , \LOSine[8] , 
            \LOSine[9] , \LOSine[10] , \LOSine[11] , \LOSine[12] , \LOCosine[1] , 
            \LOCosine[2] , \LOCosine[3] , \LOCosine[4] , \LOCosine[5] , 
            \LOCosine[6] , \LOCosine[7] , \LOCosine[8] , \LOCosine[9] , 
            \LOCosine[10] , \LOCosine[11] , \LOCosine[12] , \phase_accum[56] ) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input osc_clk;
    input VCC_net;
    input GND_net;
    input \phase_accum[57] ;
    input \phase_accum[58] ;
    input \phase_accum[59] ;
    input \phase_accum[60] ;
    input \phase_accum[61] ;
    input \phase_accum[62] ;
    input \phase_accum[63] ;
    output \LOSine[1] ;
    output \LOSine[2] ;
    output \LOSine[3] ;
    output \LOSine[4] ;
    output \LOSine[5] ;
    output \LOSine[6] ;
    output \LOSine[7] ;
    output \LOSine[8] ;
    output \LOSine[9] ;
    output \LOSine[10] ;
    output \LOSine[11] ;
    output \LOSine[12] ;
    output \LOCosine[1] ;
    output \LOCosine[2] ;
    output \LOCosine[3] ;
    output \LOCosine[4] ;
    output \LOCosine[5] ;
    output \LOCosine[6] ;
    output \LOCosine[7] ;
    output \LOCosine[8] ;
    output \LOCosine[9] ;
    output \LOCosine[10] ;
    output \LOCosine[11] ;
    output \LOCosine[12] ;
    input \phase_accum[56] ;
    
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(55[8:15])
    
    wire rom_addr0_r_1, rom_addr0_r_1_inv, rom_addr0_r_2, rom_addr0_r_3, 
        rom_addr0_r_4, rom_addr0_r_5, mx_ctrl_r, mx_ctrl_r_1, rom_addr0_r, 
        rom_addr0_r_n, rom_addr0_r_6, rom_dout_11, rom_dout_11_ffin, 
        rom_dout_10, rom_dout_10_ffin, rom_dout_9, rom_dout_9_ffin, 
        rom_dout_8, rom_dout_8_ffin, rom_dout_7, rom_dout_7_ffin, rom_dout_6, 
        rom_dout_6_ffin, rom_dout_5, rom_dout_5_ffin, rom_dout_4, rom_dout_4_ffin, 
        rom_dout_3, rom_dout_3_ffin, rom_dout_2, rom_dout_2_ffin, rom_dout_1, 
        rom_dout_1_ffin, rom_dout, rom_dout_ffin, rom_dout_25, rom_dout_25_ffin, 
        rom_dout_24, rom_dout_24_ffin, rom_dout_23, rom_dout_23_ffin, 
        rom_dout_22, rom_dout_22_ffin, rom_dout_21, rom_dout_21_ffin, 
        rom_dout_20, rom_dout_20_ffin, rom_dout_19, rom_dout_19_ffin, 
        rom_dout_18, rom_dout_18_ffin, rom_dout_17, rom_dout_17_ffin, 
        rom_dout_16, rom_dout_16_ffin, rom_dout_15, rom_dout_15_ffin, 
        rom_dout_14, rom_dout_14_ffin, rom_dout_13, rom_dout_13_ffin, 
        cosromoutsel_i, cosromoutsel, sinromoutsel, sinout_pre_1, sinout_pre_2, 
        sinout_pre_3, sinout_pre_4, sinout_pre_5, sinout_pre_6, sinout_pre_7, 
        sinout_pre_8, sinout_pre_9, sinout_pre_10, sinout_pre_11, sinout_pre_12, 
        cosout_pre_1, cosout_pre_2, cosout_pre_3, cosout_pre_4, cosout_pre_5, 
        cosout_pre_6, cosout_pre_7, cosout_pre_8, cosout_pre_9, cosout_pre_10, 
        cosout_pre_11, cosout_pre_12, rom_addr0_r_inv, co0, rom_addr0_r_n_1, 
        rom_addr0_r_n_2, rom_addr0_r_2_inv, co1, rom_addr0_r_n_3, rom_addr0_r_n_4, 
        rom_addr0_r_3_inv, rom_addr0_r_4_inv, co2, rom_addr0_r_n_5, 
        rom_addr0_r_5_inv, rom_dout_12_ffin, rom_addr0_r_7, rom_addr0_r_8, 
        rom_addr0_r_9, rom_addr0_r_10, rom_addr0_r_11, rom_dout_s_n_1, 
        rom_dout_s_n_2, co0_1, rom_dout_1_inv, rom_dout_2_inv, co1_1, 
        rom_dout_s_n_3, rom_dout_s_n_4, rom_dout_3_inv, rom_dout_4_inv, 
        co2_1, rom_dout_s_n_5, rom_dout_s_n_6, rom_dout_5_inv, rom_dout_6_inv, 
        co3, rom_dout_s_n_7, rom_dout_s_n_8, rom_dout_7_inv, rom_dout_8_inv, 
        co4, rom_dout_s_n_9, rom_dout_s_n_10, rom_dout_9_inv, rom_dout_10_inv, 
        co5, rom_dout_s_n_11, rom_dout_s_n_12, rom_dout_11_inv, rom_dout_12_inv, 
        rom_dout_13_inv, co0_2, rom_dout_c_n_1, rom_dout_c_n_2, rom_dout_14_inv, 
        rom_dout_15_inv, co1_2, rom_dout_c_n_3, rom_dout_c_n_4, rom_dout_16_inv, 
        rom_dout_17_inv, co2_2, rom_dout_c_n_5, rom_dout_c_n_6, rom_dout_18_inv, 
        rom_dout_19_inv, co3_1, rom_dout_c_n_7, rom_dout_c_n_8, rom_dout_20_inv, 
        rom_dout_21_inv, co4_1, rom_dout_c_n_9, rom_dout_c_n_10, rom_dout_22_inv, 
        rom_dout_23_inv, co5_1, rom_dout_c_n_11, rom_dout_c_n_12, rom_dout_24_inv, 
        rom_dout_25_inv, rom_dout_12, rom_dout_inv, func_or_inet, lx_ne0, 
        lx_ne0_inv, out_sel_i, rom_dout_s_1, rom_dout_s_2, rom_dout_s_3, 
        rom_dout_s_4, rom_dout_s_5, rom_dout_s_6, rom_dout_s_7, rom_dout_s_8, 
        rom_dout_s_9, rom_dout_s_10, rom_dout_s_11, rom_dout_s_12, rom_dout_c_1, 
        rom_dout_c_2, rom_dout_c_3, rom_dout_c_4, rom_dout_c_5, rom_dout_c_6, 
        rom_dout_c_7, rom_dout_c_8, rom_dout_c_9, rom_dout_c_10, rom_dout_c_11, 
        rom_dout_c_12, out_sel;
    
    INV INV_29 (.A(rom_addr0_r_1), .Z(rom_addr0_r_1_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    FD1P3DX FF_61 (.D(\phase_accum[57] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(rom_addr0_r_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(312[13:88])
    defparam FF_61.GSR = "ENABLED";
    FD1P3DX FF_60 (.D(\phase_accum[58] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(rom_addr0_r_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(315[13:88])
    defparam FF_60.GSR = "ENABLED";
    FD1P3DX FF_59 (.D(\phase_accum[59] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(rom_addr0_r_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(318[13:88])
    defparam FF_59.GSR = "ENABLED";
    FD1P3DX FF_58 (.D(\phase_accum[60] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(rom_addr0_r_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(321[13:88])
    defparam FF_58.GSR = "ENABLED";
    FD1P3DX FF_57 (.D(\phase_accum[61] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(rom_addr0_r_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(324[13:88])
    defparam FF_57.GSR = "ENABLED";
    FD1P3DX FF_56 (.D(\phase_accum[62] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(mx_ctrl_r)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(327[13:84])
    defparam FF_56.GSR = "ENABLED";
    FD1P3DX FF_55 (.D(\phase_accum[63] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(mx_ctrl_r_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(330[13:86])
    defparam FF_55.GSR = "ENABLED";
    MUX21 muxb_57 (.D0(rom_addr0_r), .D1(rom_addr0_r_n), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    FD1P3DX FF_53 (.D(rom_dout_11_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(355[13] 356[25])
    defparam FF_53.GSR = "ENABLED";
    FD1P3DX FF_52 (.D(rom_dout_10_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(359[13] 360[25])
    defparam FF_52.GSR = "ENABLED";
    FD1P3DX FF_51 (.D(rom_dout_9_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(363[13] 364[24])
    defparam FF_51.GSR = "ENABLED";
    FD1P3DX FF_50 (.D(rom_dout_8_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(367[13] 368[24])
    defparam FF_50.GSR = "ENABLED";
    FD1P3DX FF_49 (.D(rom_dout_7_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(371[13] 372[24])
    defparam FF_49.GSR = "ENABLED";
    FD1P3DX FF_48 (.D(rom_dout_6_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(375[13] 376[24])
    defparam FF_48.GSR = "ENABLED";
    FD1P3DX FF_47 (.D(rom_dout_5_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(379[13] 380[24])
    defparam FF_47.GSR = "ENABLED";
    FD1P3DX FF_46 (.D(rom_dout_4_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(383[13] 384[24])
    defparam FF_46.GSR = "ENABLED";
    FD1P3DX FF_45 (.D(rom_dout_3_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(387[13] 388[24])
    defparam FF_45.GSR = "ENABLED";
    FD1P3DX FF_44 (.D(rom_dout_2_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(391[13] 392[24])
    defparam FF_44.GSR = "ENABLED";
    FD1P3DX FF_43 (.D(rom_dout_1_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(395[13] 396[24])
    defparam FF_43.GSR = "ENABLED";
    FD1P3DX FF_42 (.D(rom_dout_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(399[13] 400[22])
    defparam FF_42.GSR = "ENABLED";
    FD1P3DX FF_41 (.D(rom_dout_25_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_25)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(403[13] 404[25])
    defparam FF_41.GSR = "ENABLED";
    FD1P3DX FF_40 (.D(rom_dout_24_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_24)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(407[13] 408[25])
    defparam FF_40.GSR = "ENABLED";
    FD1P3DX FF_39 (.D(rom_dout_23_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_23)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(411[13] 412[25])
    defparam FF_39.GSR = "ENABLED";
    FD1P3DX FF_38 (.D(rom_dout_22_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_22)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(415[13] 416[25])
    defparam FF_38.GSR = "ENABLED";
    FD1P3DX FF_37 (.D(rom_dout_21_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(419[13] 420[25])
    defparam FF_37.GSR = "ENABLED";
    FD1P3DX FF_36 (.D(rom_dout_20_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(423[13] 424[25])
    defparam FF_36.GSR = "ENABLED";
    FD1P3DX FF_35 (.D(rom_dout_19_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(427[13] 428[25])
    defparam FF_35.GSR = "ENABLED";
    FD1P3DX FF_34 (.D(rom_dout_18_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(431[13] 432[25])
    defparam FF_34.GSR = "ENABLED";
    FD1P3DX FF_33 (.D(rom_dout_17_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(435[13] 436[25])
    defparam FF_33.GSR = "ENABLED";
    FD1P3DX FF_32 (.D(rom_dout_16_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(439[13] 440[25])
    defparam FF_32.GSR = "ENABLED";
    FD1P3DX FF_31 (.D(rom_dout_15_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(443[13] 444[25])
    defparam FF_31.GSR = "ENABLED";
    FD1P3DX FF_30 (.D(rom_dout_14_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(447[13] 448[25])
    defparam FF_30.GSR = "ENABLED";
    FD1P3DX FF_29 (.D(rom_dout_13_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(451[13] 452[25])
    defparam FF_29.GSR = "ENABLED";
    FD1P3DX FF_28 (.D(cosromoutsel_i), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(cosromoutsel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(455[13] 456[26])
    defparam FF_28.GSR = "ENABLED";
    FD1P3DX FF_27 (.D(mx_ctrl_r_1), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(sinromoutsel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(459[13] 460[26])
    defparam FF_27.GSR = "ENABLED";
    FD1P3DX FF_24 (.D(sinout_pre_1), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[1] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(599[13] 600[21])
    defparam FF_24.GSR = "ENABLED";
    FD1P3DX FF_23 (.D(sinout_pre_2), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[2] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(603[13] 604[21])
    defparam FF_23.GSR = "ENABLED";
    FD1P3DX FF_22 (.D(sinout_pre_3), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[3] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(607[13] 608[21])
    defparam FF_22.GSR = "ENABLED";
    FD1P3DX FF_21 (.D(sinout_pre_4), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[4] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(611[13] 612[21])
    defparam FF_21.GSR = "ENABLED";
    FD1P3DX FF_20 (.D(sinout_pre_5), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[5] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(615[13] 616[21])
    defparam FF_20.GSR = "ENABLED";
    FD1P3DX FF_19 (.D(sinout_pre_6), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[6] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(619[13] 620[21])
    defparam FF_19.GSR = "ENABLED";
    FD1P3DX FF_18 (.D(sinout_pre_7), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[7] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(623[13] 624[21])
    defparam FF_18.GSR = "ENABLED";
    FD1P3DX FF_17 (.D(sinout_pre_8), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[8] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(627[13] 628[21])
    defparam FF_17.GSR = "ENABLED";
    FD1P3DX FF_16 (.D(sinout_pre_9), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[9] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(631[13] 632[21])
    defparam FF_16.GSR = "ENABLED";
    FD1P3DX FF_15 (.D(sinout_pre_10), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[10] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(635[13] 636[22])
    defparam FF_15.GSR = "ENABLED";
    FD1P3DX FF_14 (.D(sinout_pre_11), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[11] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(639[13] 640[22])
    defparam FF_14.GSR = "ENABLED";
    FD1P3DX FF_13 (.D(sinout_pre_12), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOSine[12] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(643[13] 644[22])
    defparam FF_13.GSR = "ENABLED";
    FD1P3DX FF_11 (.D(cosout_pre_1), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[1] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(650[13] 651[23])
    defparam FF_11.GSR = "ENABLED";
    FD1P3DX FF_10 (.D(cosout_pre_2), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[2] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(654[13] 655[23])
    defparam FF_10.GSR = "ENABLED";
    FD1P3DX FF_9 (.D(cosout_pre_3), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[3] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(658[13] 659[23])
    defparam FF_9.GSR = "ENABLED";
    FD1P3DX FF_8 (.D(cosout_pre_4), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[4] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(662[13] 663[23])
    defparam FF_8.GSR = "ENABLED";
    FD1P3DX FF_7 (.D(cosout_pre_5), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[5] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(666[13] 667[23])
    defparam FF_7.GSR = "ENABLED";
    FD1P3DX FF_6 (.D(cosout_pre_6), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[6] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(670[13] 671[23])
    defparam FF_6.GSR = "ENABLED";
    FD1P3DX FF_5 (.D(cosout_pre_7), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[7] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(674[13] 675[23])
    defparam FF_5.GSR = "ENABLED";
    FD1P3DX FF_4 (.D(cosout_pre_8), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[8] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(678[13] 679[23])
    defparam FF_4.GSR = "ENABLED";
    FD1P3DX FF_3 (.D(cosout_pre_9), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[9] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(682[13] 683[23])
    defparam FF_3.GSR = "ENABLED";
    FD1P3DX FF_2 (.D(cosout_pre_10), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[10] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(686[13] 687[24])
    defparam FF_2.GSR = "ENABLED";
    FD1P3DX FF_1 (.D(cosout_pre_11), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[11] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(690[13] 691[24])
    defparam FF_1.GSR = "ENABLED";
    FD1P3DX FF_0 (.D(cosout_pre_12), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(\LOCosine[12] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(694[13] 695[24])
    defparam FF_0.GSR = "ENABLED";
    FADD2B neg_rom_addr0_r_n_0 (.A0(GND_net), .A1(rom_addr0_r_inv), .B0(GND_net), 
           .B1(VCC_net), .CI(GND_net), .COUT(co0), .S1(rom_addr0_r_n)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    FADD2B neg_rom_addr0_r_n_1 (.A0(rom_addr0_r_1_inv), .A1(rom_addr0_r_2_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co0), .COUT(co1), .S0(rom_addr0_r_n_1), 
           .S1(rom_addr0_r_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    FADD2B neg_rom_addr0_r_n_2 (.A0(rom_addr0_r_3_inv), .A1(rom_addr0_r_4_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co1), .COUT(co2), .S0(rom_addr0_r_n_3), 
           .S1(rom_addr0_r_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    FADD2B neg_rom_addr0_r_n_3 (.A0(rom_addr0_r_5_inv), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co2), .S0(rom_addr0_r_n_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    ROM64X1A triglut_1_0_25 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_12_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_25.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    FADD2B neg_rom_dout_s_n_1 (.A0(rom_dout_1_inv), .A1(rom_dout_2_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co0_1), .COUT(co1_1), .S0(rom_dout_s_n_1), 
           .S1(rom_dout_s_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    FADD2B neg_rom_dout_s_n_2 (.A0(rom_dout_3_inv), .A1(rom_dout_4_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co1_1), .COUT(co2_1), .S0(rom_dout_s_n_3), 
           .S1(rom_dout_s_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    FADD2B neg_rom_dout_s_n_3 (.A0(rom_dout_5_inv), .A1(rom_dout_6_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co2_1), .COUT(co3), .S0(rom_dout_s_n_5), 
           .S1(rom_dout_s_n_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    FADD2B neg_rom_dout_s_n_4 (.A0(rom_dout_7_inv), .A1(rom_dout_8_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co3), .COUT(co4), .S0(rom_dout_s_n_7), 
           .S1(rom_dout_s_n_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    FADD2B neg_rom_dout_s_n_5 (.A0(rom_dout_9_inv), .A1(rom_dout_10_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co4), .COUT(co5), .S0(rom_dout_s_n_9), 
           .S1(rom_dout_s_n_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    FADD2B neg_rom_dout_s_n_6 (.A0(rom_dout_11_inv), .A1(rom_dout_12_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co5), .S0(rom_dout_s_n_11), 
           .S1(rom_dout_s_n_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_30 (.A(rom_addr0_r_2), .Z(rom_addr0_r_2_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    FADD2B neg_rom_dout_c_n_0 (.A0(GND_net), .A1(rom_dout_13_inv), .B0(GND_net), 
           .B1(VCC_net), .CI(GND_net), .COUT(co0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    FADD2B neg_rom_dout_c_n_1 (.A0(rom_dout_14_inv), .A1(rom_dout_15_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co0_2), .COUT(co1_2), .S0(rom_dout_c_n_1), 
           .S1(rom_dout_c_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    FADD2B neg_rom_dout_c_n_2 (.A0(rom_dout_16_inv), .A1(rom_dout_17_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co1_2), .COUT(co2_2), .S0(rom_dout_c_n_3), 
           .S1(rom_dout_c_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    FADD2B neg_rom_dout_c_n_3 (.A0(rom_dout_18_inv), .A1(rom_dout_19_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co2_2), .COUT(co3_1), .S0(rom_dout_c_n_5), 
           .S1(rom_dout_c_n_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    FADD2B neg_rom_dout_c_n_4 (.A0(rom_dout_20_inv), .A1(rom_dout_21_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co3_1), .COUT(co4_1), .S0(rom_dout_c_n_7), 
           .S1(rom_dout_c_n_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    FADD2B neg_rom_dout_c_n_5 (.A0(rom_dout_22_inv), .A1(rom_dout_23_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co4_1), .COUT(co5_1), .S0(rom_dout_c_n_9), 
           .S1(rom_dout_c_n_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    FADD2B neg_rom_dout_c_n_6 (.A0(rom_dout_24_inv), .A1(rom_dout_25_inv), 
           .B0(GND_net), .B1(GND_net), .CI(co5_1), .S0(rom_dout_c_n_11), 
           .S1(rom_dout_c_n_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_31 (.A(rom_addr0_r_3), .Z(rom_addr0_r_3_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_32 (.A(rom_addr0_r_4), .Z(rom_addr0_r_4_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_33 (.A(rom_addr0_r_5), .Z(rom_addr0_r_5_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_28 (.A(rom_addr0_r), .Z(rom_addr0_r_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    XOR2 XOR2_t1 (.A(mx_ctrl_r), .B(mx_ctrl_r_1), .Z(cosromoutsel_i)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(241[10:70])
    INV INV_27 (.A(rom_dout_12), .Z(rom_dout_12_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_26 (.A(rom_dout_11), .Z(rom_dout_11_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_25 (.A(rom_dout_10), .Z(rom_dout_10_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_24 (.A(rom_dout_9), .Z(rom_dout_9_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_23 (.A(rom_dout_8), .Z(rom_dout_8_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_22 (.A(rom_dout_7), .Z(rom_dout_7_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_21 (.A(rom_dout_6), .Z(rom_dout_6_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_20 (.A(rom_dout_5), .Z(rom_dout_5_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_19 (.A(rom_dout_4), .Z(rom_dout_4_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_18 (.A(rom_dout_3), .Z(rom_dout_3_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_17 (.A(rom_dout_2), .Z(rom_dout_2_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_16 (.A(rom_dout_1), .Z(rom_dout_1_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_15 (.A(rom_dout), .Z(rom_dout_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_14 (.A(rom_dout_25), .Z(rom_dout_25_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_13 (.A(rom_dout_24), .Z(rom_dout_24_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_12 (.A(rom_dout_23), .Z(rom_dout_23_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_11 (.A(rom_dout_22), .Z(rom_dout_22_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_10 (.A(rom_dout_21), .Z(rom_dout_21_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_9 (.A(rom_dout_20), .Z(rom_dout_20_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_8 (.A(rom_dout_19), .Z(rom_dout_19_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_7 (.A(rom_dout_18), .Z(rom_dout_18_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_6 (.A(rom_dout_17), .Z(rom_dout_17_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_5 (.A(rom_dout_16), .Z(rom_dout_16_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_4 (.A(rom_dout_15), .Z(rom_dout_15_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_3 (.A(rom_dout_14), .Z(rom_dout_14_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    INV INV_2 (.A(rom_dout_13), .Z(rom_dout_13_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    ROM16X1A LUT4_1 (.AD0(rom_addr0_r_9), .AD1(rom_addr0_r_8), .AD2(rom_addr0_r_7), 
            .AD3(rom_addr0_r_6), .DO0(func_or_inet)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam LUT4_1.initval = 16'b1111111111111110;
    ROM16X1A LUT4_0 (.AD0(GND_net), .AD1(rom_addr0_r_11), .AD2(rom_addr0_r_10), 
            .AD3(func_or_inet), .DO0(lx_ne0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam LUT4_0.initval = 16'b1111111111111110;
    INV INV_1 (.A(lx_ne0), .Z(lx_ne0_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    AND2 AND2_t0 (.A(mx_ctrl_r), .B(lx_ne0_inv), .Z(out_sel_i)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(305[10:64])
    FD1P3DX FF_62 (.D(\phase_accum[56] ), .SP(VCC_net), .CK(osc_clk), 
            .CD(GND_net), .Q(rom_addr0_r)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(309[13:86])
    defparam FF_62.GSR = "ENABLED";
    MUX21 muxb_56 (.D0(rom_addr0_r_1), .D1(rom_addr0_r_n_1), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_55 (.D0(rom_addr0_r_2), .D1(rom_addr0_r_n_2), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_54 (.D0(rom_addr0_r_3), .D1(rom_addr0_r_n_3), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_53 (.D0(rom_addr0_r_4), .D1(rom_addr0_r_n_4), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_52 (.D0(rom_addr0_r_5), .D1(rom_addr0_r_n_5), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    FD1P3DX FF_54 (.D(rom_dout_12_ffin), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(rom_dout_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(351[13] 352[25])
    defparam FF_54.GSR = "ENABLED";
    MUX21 muxb_50 (.D0(rom_dout_1), .D1(rom_dout_s_n_1), .SD(sinromoutsel), 
          .Z(rom_dout_s_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_49 (.D0(rom_dout_2), .D1(rom_dout_s_n_2), .SD(sinromoutsel), 
          .Z(rom_dout_s_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_48 (.D0(rom_dout_3), .D1(rom_dout_s_n_3), .SD(sinromoutsel), 
          .Z(rom_dout_s_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_47 (.D0(rom_dout_4), .D1(rom_dout_s_n_4), .SD(sinromoutsel), 
          .Z(rom_dout_s_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_46 (.D0(rom_dout_5), .D1(rom_dout_s_n_5), .SD(sinromoutsel), 
          .Z(rom_dout_s_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_45 (.D0(rom_dout_6), .D1(rom_dout_s_n_6), .SD(sinromoutsel), 
          .Z(rom_dout_s_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_44 (.D0(rom_dout_7), .D1(rom_dout_s_n_7), .SD(sinromoutsel), 
          .Z(rom_dout_s_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_43 (.D0(rom_dout_8), .D1(rom_dout_s_n_8), .SD(sinromoutsel), 
          .Z(rom_dout_s_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_42 (.D0(rom_dout_9), .D1(rom_dout_s_n_9), .SD(sinromoutsel), 
          .Z(rom_dout_s_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_41 (.D0(rom_dout_10), .D1(rom_dout_s_n_10), .SD(sinromoutsel), 
          .Z(rom_dout_s_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_40 (.D0(rom_dout_11), .D1(rom_dout_s_n_11), .SD(sinromoutsel), 
          .Z(rom_dout_s_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_39 (.D0(rom_dout_12), .D1(rom_dout_s_n_12), .SD(sinromoutsel), 
          .Z(rom_dout_s_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_37 (.D0(rom_dout_14), .D1(rom_dout_c_n_1), .SD(cosromoutsel), 
          .Z(rom_dout_c_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_36 (.D0(rom_dout_15), .D1(rom_dout_c_n_2), .SD(cosromoutsel), 
          .Z(rom_dout_c_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_35 (.D0(rom_dout_16), .D1(rom_dout_c_n_3), .SD(cosromoutsel), 
          .Z(rom_dout_c_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_34 (.D0(rom_dout_17), .D1(rom_dout_c_n_4), .SD(cosromoutsel), 
          .Z(rom_dout_c_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_33 (.D0(rom_dout_18), .D1(rom_dout_c_n_5), .SD(cosromoutsel), 
          .Z(rom_dout_c_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_32 (.D0(rom_dout_19), .D1(rom_dout_c_n_6), .SD(cosromoutsel), 
          .Z(rom_dout_c_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_31 (.D0(rom_dout_20), .D1(rom_dout_c_n_7), .SD(cosromoutsel), 
          .Z(rom_dout_c_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_30 (.D0(rom_dout_21), .D1(rom_dout_c_n_8), .SD(cosromoutsel), 
          .Z(rom_dout_c_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_29 (.D0(rom_dout_22), .D1(rom_dout_c_n_9), .SD(cosromoutsel), 
          .Z(rom_dout_c_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_28 (.D0(rom_dout_23), .D1(rom_dout_c_n_10), .SD(cosromoutsel), 
          .Z(rom_dout_c_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_27 (.D0(rom_dout_24), .D1(rom_dout_c_n_11), .SD(cosromoutsel), 
          .Z(rom_dout_c_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_26 (.D0(rom_dout_25), .D1(rom_dout_c_n_12), .SD(cosromoutsel), 
          .Z(rom_dout_c_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    FD1P3DX FF_26 (.D(out_sel_i), .SP(VCC_net), .CK(osc_clk), .CD(GND_net), 
            .Q(out_sel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/sincos.v(541[13:83])
    defparam FF_26.GSR = "ENABLED";
    MUX21 muxb_24 (.D0(rom_dout_s_1), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_23 (.D0(rom_dout_s_2), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_22 (.D0(rom_dout_s_3), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_21 (.D0(rom_dout_s_4), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_20 (.D0(rom_dout_s_5), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_19 (.D0(rom_dout_s_6), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_18 (.D0(rom_dout_s_7), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_17 (.D0(rom_dout_s_8), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_16 (.D0(rom_dout_s_9), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_15 (.D0(rom_dout_s_10), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_14 (.D0(rom_dout_s_11), .D1(VCC_net), .SD(out_sel), .Z(sinout_pre_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_13 (.D0(rom_dout_s_12), .D1(mx_ctrl_r_1), .SD(out_sel), 
          .Z(sinout_pre_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_11 (.D0(rom_dout_c_1), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_10 (.D0(rom_dout_c_2), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_9 (.D0(rom_dout_c_3), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_8 (.D0(rom_dout_c_4), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_7 (.D0(rom_dout_c_5), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_6 (.D0(rom_dout_c_6), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_5 (.D0(rom_dout_c_7), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_4 (.D0(rom_dout_c_8), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_3 (.D0(rom_dout_c_9), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_2 (.D0(rom_dout_c_10), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_1 (.D0(rom_dout_c_11), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    MUX21 muxb_0 (.D0(rom_dout_c_12), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    ROM64X1A triglut_1_0_24 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_11_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_24.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    ROM64X1A triglut_1_0_23 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_10_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_23.initval = 64'b1111111111111111111111111111111111111111110000000000000000000000;
    ROM64X1A triglut_1_0_22 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_9_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_22.initval = 64'b1111111111111111111111111111100000000000001111111111100000000000;
    ROM64X1A triglut_1_0_21 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_8_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_21.initval = 64'b1111111111111111111100000000011111110000001111110000011111000000;
    ROM64X1A triglut_1_0_20 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_7_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_20.initval = 64'b1111111111111100000011111000011110001110001110001110011100111000;
    ROM64X1A triglut_1_0_19 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_6_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_19.initval = 64'b1111111111000011100011100110011001001101101101001001011010110100;
    ROM64X1A triglut_1_0_18 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_5_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_18.initval = 64'b1111111000110011011010010101010100101001001001101100110001100110;
    ROM64X1A triglut_1_0_17 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_4_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_17.initval = 64'b1111100100101010110011000000000001110011011010110101010110101010;
    ROM64X1A triglut_1_0_16 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_3_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_16.initval = 64'b1110010110011100010101001111111101101010110011100000000011110000;
    ROM64X1A triglut_1_0_15 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_2_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_15.initval = 64'b1101000010100011001111010111110011001100010101100000000011001100;
    ROM64X1A triglut_1_0_14 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_1_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_14.initval = 64'b1111011011100010010110111011101001110011000000100111110010101010;
    ROM64X1A triglut_1_0_13 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_13.initval = 64'b1000100101001010011001010111111001010010011110001001001001111000;
    ROM64X1A triglut_1_0_12 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_25_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_12.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    ROM64X1A triglut_1_0_11 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_24_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_11.initval = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    ROM64X1A triglut_1_0_10 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_23_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_10.initval = 64'b0000000000000000000001111111111111111111111111111111111111111110;
    ROM64X1A triglut_1_0_9 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_22_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_9.initval = 64'b0000000000111111111110000000000000111111111111111111111111111110;
    ROM64X1A triglut_1_0_8 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_21_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_8.initval = 64'b0000011111000001111110000001111111000000000111111111111111111110;
    ROM64X1A triglut_1_0_7 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_20_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_7.initval = 64'b0011100111001110001110001110001111000011111000000111111111111110;
    ROM64X1A triglut_1_0_6 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_19_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_6.initval = 64'b0101101011010010010110110110010011001100111000111000011111111110;
    ROM64X1A triglut_1_0_5 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_18_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_5.initval = 64'b1100110001100110110010010010100101010101001011011001100011111110;
    ROM64X1A triglut_1_0_4 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_17_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_4.initval = 64'b1010101101010101101011011001110000000000011001101010100100111110;
    ROM64X1A triglut_1_0_3 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_16_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_3.initval = 64'b0001111000000000111001101010110111111110010101000111001101001110;
    ROM64X1A triglut_1_0_2 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_15_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_2.initval = 64'b0110011000000000110101000110011001111101011110011000101000010110;
    ROM64X1A triglut_1_0_1 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_14_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_1.initval = 64'b1010101001111100100000011001110010111011101101001000111011011110;
    ROM64X1A triglut_1_0_0 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_13_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    defparam triglut_1_0_0.initval = 64'b0011110010010010001111001001010011111101010011001010010100100010;
    FADD2B neg_rom_dout_s_n_0 (.A0(GND_net), .A1(rom_dout_inv), .B0(GND_net), 
           .B1(VCC_net), .CI(GND_net), .COUT(co0_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=98, LSE_RLINE=105 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(98[8] 105[2])
    
endmodule
//
// Verilog Description of module \CIC(width=72,decimation_ratio=4096) 
//

module \CIC(width=72,decimation_ratio=4096)  (osc_clk, \CICGain[1] , \CICGain[0] , 
            CIC1_out_clkSin, \CIC1_outSin[0] , MixerOutSin, GND_net, 
            \CIC1_outSin[1] , \CIC1_outSin[2] , \CIC1_outSin[3] , \CIC1_outSin[4] , 
            \CIC1_outSin[5] , MYLED_c_0, MYLED_c_1, MYLED_c_2, MYLED_c_3, 
            MYLED_c_4, MYLED_c_5, \d10[67] , \d10[68] , \d10[69] , 
            \d10[70] , n63, \d_out_11__N_1818[2] , n64, \d_out_11__N_1818[3] , 
            n70, n67, \d10[65] , n68, \d10[66] , n65, \d10[63] , 
            n66, \d10[64] , \d10[61] , \d10[62] , \d_out_11__N_1818[10] , 
            n61, \d10[59] , n62, \d10[60] , \d_out_11__N_1818[5] , 
            \d_out_11__N_1818[4] , \d_out_11__N_1818[6] , \d_out_11__N_1818[7] , 
            \d_out_11__N_1818[8] , \d_out_11__N_1818[9] , \d10[71] , \d_out_11__N_1818[11] ) /* synthesis syn_module_defined=1 */ ;
    input osc_clk;
    input \CICGain[1] ;
    input \CICGain[0] ;
    output CIC1_out_clkSin;
    output \CIC1_outSin[0] ;
    input [11:0]MixerOutSin;
    input GND_net;
    output \CIC1_outSin[1] ;
    output \CIC1_outSin[2] ;
    output \CIC1_outSin[3] ;
    output \CIC1_outSin[4] ;
    output \CIC1_outSin[5] ;
    output MYLED_c_0;
    output MYLED_c_1;
    output MYLED_c_2;
    output MYLED_c_3;
    output MYLED_c_4;
    output MYLED_c_5;
    input \d10[67] ;
    input \d10[68] ;
    input \d10[69] ;
    input \d10[70] ;
    input n63;
    output \d_out_11__N_1818[2] ;
    input n64;
    output \d_out_11__N_1818[3] ;
    input n70;
    input n67;
    input \d10[65] ;
    input n68;
    input \d10[66] ;
    input n65;
    input \d10[63] ;
    input n66;
    input \d10[64] ;
    input \d10[61] ;
    input \d10[62] ;
    output \d_out_11__N_1818[10] ;
    input n61;
    input \d10[59] ;
    input n62;
    input \d10[60] ;
    output \d_out_11__N_1818[5] ;
    output \d_out_11__N_1818[4] ;
    output \d_out_11__N_1818[6] ;
    output \d_out_11__N_1818[7] ;
    output \d_out_11__N_1818[8] ;
    output \d_out_11__N_1818[9] ;
    input \d10[71] ;
    output \d_out_11__N_1818[11] ;
    
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(55[8:15])
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(67[6:21])
    wire [71:0]d_d_tmp;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(30[33:40])
    
    wire osc_clk_enable_1395;
    wire [71:0]d_tmp;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(30[26:31])
    
    wire n65_c, n133;
    wire [71:0]d_out_11__N_1818;
    
    wire n12089;
    wire [71:0]d2;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(36[26:28])
    
    wire n4190;
    wire [35:0]n4191;
    wire [71:0]d1;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(35[26:28])
    wire [71:0]d2_71__N_489;
    
    wire n12090, osc_clk_enable_62;
    wire [71:0]d5;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(39[26:28])
    wire [71:0]d3;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(37[26:28])
    wire [71:0]d3_71__N_561;
    wire [71:0]d4;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(38[26:28])
    wire [71:0]d4_71__N_633;
    wire [71:0]d5_71__N_705;
    wire [71:0]d6;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(43[26:28])
    wire [71:0]d6_71__N_1458;
    wire [71:0]d_d6;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(43[30:34])
    
    wire n11723, n5558;
    wire [35:0]n5559;
    wire [71:0]d7_71__N_1530;
    
    wire n11724, d_clk_tmp, n8331, v_comb;
    wire [71:0]d7;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(44[26:28])
    wire [71:0]d_d7;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(44[30:34])
    wire [71:0]d8;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(45[26:28])
    wire [71:0]d8_71__N_1602;
    wire [71:0]d_d8;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(45[30:34])
    wire [71:0]d9;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(46[26:28])
    wire [71:0]d9_71__N_1674;
    wire [71:0]d_d9;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(46[30:34])
    wire [71:0]d1_71__N_417;
    wire [15:0]count;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(50[14:19])
    wire [15:0]count_15__N_1441;
    
    wire n12088, n12087, n68_c;
    wire [71:0]d10;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(47[26:29])
    
    wire n138, n12086, n12085, n12084, n12083, n12082, n12081, 
        n12080, n12079, n12078, n12073;
    wire [35:0]n4343;
    
    wire n12072, n66_c, n134, n21, n19, n15, n16, n31, n63_c, 
        n131, n64_c, n132, n11726, n11727, n11722, n11721, n11720, 
        n11719, n11718, n11717, n11716, n11715, n11714, n11713, 
        n11712, n11711, n11710, n11706;
    wire [35:0]n5711;
    
    wire n11705, n11704, n11703, n11702, n11701, n11700, n13254, 
        n11699, n11698, n11697, n12071, n11696, n11695, d_clk_tmp_N_1830, 
        n11694, n11693, n12864, n11692, n11691, n67_c, n135, n12070, 
        n61_c, n13252, n13, n13238, n14123, n12261, n4038, n11725, 
        n12260, n12259;
    wire [35:0]n4495;
    
    wire osc_clk_enable_146, n136, n11746, n11745, n11744, n11743, 
        n11742, n11741, n11740, n11739, n11738, n11737, n11736, 
        n11735, n13778, n11734, n11733, n11732, n11731, n11730, 
        n11729, n12069, n12068, n12067, n12066, n12065, n12064, 
        n12063, n12062, n12061, n12060, n12059, n12058, n12057, 
        osc_clk_enable_196, osc_clk_enable_246, osc_clk_enable_296, osc_clk_enable_346, 
        osc_clk_enable_396, osc_clk_enable_446, osc_clk_enable_496, osc_clk_enable_546, 
        osc_clk_enable_596, osc_clk_enable_646, osc_clk_enable_696;
    wire [71:0]d10_71__N_1746;
    
    wire n12054, n4342, n12053, n12052, n12051, n12050, n12049, 
        n12048, n12047, n12046, n12045, n12044, n12043, n8367;
    wire [15:0]n375;
    
    wire n12258, n12257, n12256, n11408;
    wire [35:0]n6319;
    
    wire n11407, n11406, n11405, n11404, n11403, n11402, n11401, 
        n11400, n11399, n11398, n11397, n11396, n11395, n11394, 
        n11393, n11392, n11391, n11390;
    wire [35:0]n6357;
    
    wire n11389, n11388, n11387, n11386, n11385, n11384, n11383, 
        n11382, n11381, n11380, n11379, n11378, n11377, n11376, 
        n11375, n11374, n11373, n11372;
    wire [35:0]n6471;
    
    wire n11371, n11370, n11369, n11368, n11367, n11366, n11365, 
        n11364, n11363, n11362, n11361, n11360, n11359, n11358, 
        n11357, n12042, n12255, n11690, n12254, n12253, n12252, 
        n12251, n12250, n12249, n12248, n12041, n12040, n12039, 
        n12038, n12037, n12032, n12031, n12247, n12246, n13777, 
        n7, n12245, n12244, n12030, n11689, n12029, n11687, n5710, 
        n11686, n11685, n12028, n12027, n12026, n12025, n12024, 
        n12023, n12022;
    wire [35:0]n4647;
    
    wire n137, n12021, n12020, n11684, n11683, n11682, n12019, 
        n11681, n11356, n11355, n11353, n6470, n11352, n11351, 
        n11350, n11349, n11348, n11347, n11346, n11345, n11344, 
        n11343, n11342, n11341, n11340, n11339, n11338, n11337, 
        n11336, n11256;
    wire [35:0]n6927;
    
    wire n11255, n11254, n11253, n11252, n11251, n11250, n11249, 
        n11248, n11247, n11246, n11245, n11244, n11243, n11242, 
        n11241, n11240, n11239, n11237, n6926, n11236, n11235, 
        n11234, n11233, n11232, n11231, n11230, n11229, n11228, 
        n11227, n11226, n11225, n11224, n11223, n11222, n11221, 
        n11220, n11189;
    wire [35:0]n4077;
    
    wire n11188, n11187, n11186, n11185, n11184, n6318, n62_c, 
        n12018, n12017, n12016, n13799, n13798, n12013, n4494, 
        n12116, n12012, n12011, n12010, n12009, n12008, n12007, 
        n12006, n12005, n12004, n11680, n11679, n11678, n11677, 
        n11676, n11675, n11674, n11673, n11672, n11671, n11670, 
        n70_c, n13808, n13807, n11183, n11182, n11181, n11180, 
        n11179, n11178, n11177, n11176, n11175, n11174, n11173, 
        n11172, n11168, n11167, n11166, n11165, n11164, n11163, 
        n11162, n11161, n11160, n11159, n11158, n11157, n11156, 
        n11155, n11154, n11153, n11152, n11151, n11109, n11108, 
        n11107, n11106, n11105, n11104, n11103, n11102, n11101, 
        n11100, n11099, n11098, n11097, n11096, n11095, n11094, 
        n11093, n11092, n11091, n11090, n11089, n11088, n11087, 
        n11086, n11085, n11084, n11083, n11082, n11081, n11080, 
        n11079, n11078, n11077, n11076, n11075, n11074, n11019, 
        n11018, n11017, n11016, n11015, n11014, n11013, n11012, 
        n11011, n11010, n11009, n11008, n11007, n11006, n11005, 
        n11004, n11003, n11002, n10980, n10979, n10978, n10977, 
        n10976, n10975, n10974, n10973, n10972, n10971, n10970, 
        n10969, n10968, n10967, n10966, n10965, n10964, n10963, 
        n10886, n10885, n10884, n10883, n10882, n10881, n10880, 
        n10879, n10859, n4646, n10858, n10857, n10856, n10855, 
        n10854, n10853, n10852, n10851, n10850, n10849, n10848, 
        n10847, n10846, n10845, n10844, n10843, n10842, n10840, 
        n10839, n10838, n10837, n10836, n10835, n10834, n10833, 
        n10832, n10831, n10830, n10829, n10828, n10827, n10826, 
        n10825, n10824, n10823, n10821, n10820, n10819, n10818, 
        n10817, n10816, n10815, n10814, n10813, n10812, n10811, 
        n10810, n10809, n10808, n10807, n10806, n10805, n10804, 
        n10802, n10801, n10800, n10799, n10798, n10797, n10796, 
        n10795, n10794, n10793, n10792, n10791, n10790, n10789, 
        n10788, n10787, n10786, n10785, n140, n131_adj_2576, n13820, 
        n13819, n132_adj_2579, n12003, n140_adj_2582, n137_adj_2585, 
        n138_adj_2588, n135_adj_2591, n136_adj_2594, n133_adj_2596, 
        n134_adj_2598, n12002, n12001, n12000, n11999, n11998, n11997, 
        n11996, n11991, n11990, n11989, n11988, n11987, n11986, 
        n11985, n11984, n11983, n11982, n11981, n12134, n12133, 
        n12132, n12131, n12130, n12129, n12128, n12127, n12126, 
        n12125, n12124, n12123, n12122, n11980, n12121, n12120, 
        n12119, n11979, n12118, n11978, n12114, n12113, n11977, 
        n12112, n12111, n12110, n12109, n12108, n12107, n12106, 
        n12105, n12104, n12103, n12102, n12101, n12100, n12099, 
        n11976, n12098, n12095, n12094, n11975, n12093, n11972, 
        n11971, n11970, n11969, n11968, n11967, n11966, n11965, 
        n11964, n12092, n11963, n11962, n11961, n11960, n11959, 
        n11958, n11957, n11956, n11955, n12091;
    
    FD1P3AX d_d_tmp_i0_i4 (.D(d_tmp[4]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i3 (.D(d_tmp[3]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i2 (.D(d_tmp[2]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i1 (.D(d_tmp[1]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i1.GSR = "ENABLED";
    LUT4 shift_right_31_i205_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65_c), .D(n133), .Z(d_out_11__N_1818[4])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i205_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_989_25 (.A0(d2[58]), .B0(n4190), .C0(n4191[22]), .D0(d1[58]), 
          .A1(d2[59]), .B1(n4190), .C1(n4191[23]), .D1(d1[59]), .CIN(n12089), 
          .COUT(n12090), .S0(d2_71__N_489[58]), .S1(d2_71__N_489[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_989_25.INIT0 = 16'h74b8;
    defparam add_989_25.INIT1 = 16'h74b8;
    defparam add_989_25.INJECT1_0 = "NO";
    defparam add_989_25.INJECT1_1 = "NO";
    FD1P3AX d_d_tmp_i0_i0 (.D(d_tmp[0]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i0.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i71 (.D(d5[71]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i70 (.D(d5[70]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i69 (.D(d5[69]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i69.GSR = "ENABLED";
    FD1S3AX d2_i0 (.D(d2_71__N_489[0]), .CK(osc_clk), .Q(d2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i0.GSR = "ENABLED";
    FD1S3AX d3_i0 (.D(d3_71__N_561[0]), .CK(osc_clk), .Q(d3[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i0.GSR = "ENABLED";
    FD1S3AX d4_i0 (.D(d4_71__N_633[0]), .CK(osc_clk), .Q(d4[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i0.GSR = "ENABLED";
    FD1S3AX d5_i0 (.D(d5_71__N_705[0]), .CK(osc_clk), .Q(d5[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i0.GSR = "ENABLED";
    FD1P3AX d6_i0_i0 (.D(d6_71__N_1458[0]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i0 (.D(d6[0]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i0.GSR = "ENABLED";
    CCU2D add_1034_29 (.A0(d_d6[62]), .B0(n5558), .C0(n5559[26]), .D0(d6[62]), 
          .A1(d_d6[63]), .B1(n5558), .C1(n5559[27]), .D1(d6[63]), .CIN(n11723), 
          .COUT(n11724), .S0(d7_71__N_1530[62]), .S1(d7_71__N_1530[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1034_29.INIT0 = 16'hb874;
    defparam add_1034_29.INIT1 = 16'hb874;
    defparam add_1034_29.INJECT1_0 = "NO";
    defparam add_1034_29.INJECT1_1 = "NO";
    FD1S3JX d_clk_tmp_65 (.D(n8331), .CK(osc_clk), .PD(osc_clk_enable_62), 
            .Q(d_clk_tmp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_clk_tmp_65.GSR = "ENABLED";
    FD1S3AX v_comb_66 (.D(osc_clk_enable_62), .CK(osc_clk), .Q(v_comb)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66.GSR = "ENABLED";
    FD1S3AX d_clk_67 (.D(d_clk_tmp), .CK(osc_clk), .Q(CIC1_out_clkSin)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_clk_67.GSR = "ENABLED";
    FD1P3AX d7_i0_i0 (.D(d7_71__N_1530[0]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i0 (.D(d7[0]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d8_i0_i0 (.D(d8_71__N_1602[0]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i0 (.D(d8[0]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d9_i0_i0 (.D(d9_71__N_1674[0]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i0 (.D(d9[0]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_out_i0_i0 (.D(d_out_11__N_1818[0]), .SP(osc_clk_enable_1395), 
            .CK(osc_clk), .Q(\CIC1_outSin[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i0.GSR = "ENABLED";
    FD1S3AX d1_i0 (.D(d1_71__N_417[0]), .CK(osc_clk), .Q(d1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i0.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i68 (.D(d5[68]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i68.GSR = "ENABLED";
    FD1S3IX count__i0 (.D(count_15__N_1441[0]), .CK(osc_clk), .CD(osc_clk_enable_62), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i0.GSR = "ENABLED";
    LUT4 i4828_2_lut (.A(MixerOutSin[0]), .B(d1[0]), .Z(d1_71__N_417[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4828_2_lut.init = 16'h6666;
    FD1P3AX d_tmp_i0_i67 (.D(d5[67]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i67.GSR = "ENABLED";
    CCU2D add_989_23 (.A0(d2[56]), .B0(n4190), .C0(n4191[20]), .D0(d1[56]), 
          .A1(d2[57]), .B1(n4190), .C1(n4191[21]), .D1(d1[57]), .CIN(n12088), 
          .COUT(n12089), .S0(d2_71__N_489[56]), .S1(d2_71__N_489[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_989_23.INIT0 = 16'h74b8;
    defparam add_989_23.INIT1 = 16'h74b8;
    defparam add_989_23.INJECT1_0 = "NO";
    defparam add_989_23.INJECT1_1 = "NO";
    CCU2D add_989_21 (.A0(d2[54]), .B0(n4190), .C0(n4191[18]), .D0(d1[54]), 
          .A1(d2[55]), .B1(n4190), .C1(n4191[19]), .D1(d1[55]), .CIN(n12087), 
          .COUT(n12088), .S0(d2_71__N_489[54]), .S1(d2_71__N_489[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_989_21.INIT0 = 16'h74b8;
    defparam add_989_21.INIT1 = 16'h74b8;
    defparam add_989_21.INJECT1_0 = "NO";
    defparam add_989_21.INJECT1_1 = "NO";
    FD1P3AX d_tmp_i0_i66 (.D(d5[66]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i65 (.D(d5[65]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i65.GSR = "ENABLED";
    LUT4 shift_right_31_i138_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n68_c), .D(d10[66]), .Z(n138)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i138_3_lut_4_lut.init = 16'hf960;
    FD1P3AX d_tmp_i0_i64 (.D(d5[64]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i64.GSR = "ENABLED";
    CCU2D add_989_19 (.A0(d2[52]), .B0(n4190), .C0(n4191[16]), .D0(d1[52]), 
          .A1(d2[53]), .B1(n4190), .C1(n4191[17]), .D1(d1[53]), .CIN(n12086), 
          .COUT(n12087), .S0(d2_71__N_489[52]), .S1(d2_71__N_489[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_989_19.INIT0 = 16'h74b8;
    defparam add_989_19.INIT1 = 16'h74b8;
    defparam add_989_19.INJECT1_0 = "NO";
    defparam add_989_19.INJECT1_1 = "NO";
    CCU2D add_989_17 (.A0(d2[50]), .B0(n4190), .C0(n4191[14]), .D0(d1[50]), 
          .A1(d2[51]), .B1(n4190), .C1(n4191[15]), .D1(d1[51]), .CIN(n12085), 
          .COUT(n12086), .S0(d2_71__N_489[50]), .S1(d2_71__N_489[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_989_17.INIT0 = 16'h74b8;
    defparam add_989_17.INIT1 = 16'h74b8;
    defparam add_989_17.INJECT1_0 = "NO";
    defparam add_989_17.INJECT1_1 = "NO";
    CCU2D add_989_15 (.A0(d2[48]), .B0(n4190), .C0(n4191[12]), .D0(d1[48]), 
          .A1(d2[49]), .B1(n4190), .C1(n4191[13]), .D1(d1[49]), .CIN(n12084), 
          .COUT(n12085), .S0(d2_71__N_489[48]), .S1(d2_71__N_489[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_989_15.INIT0 = 16'h74b8;
    defparam add_989_15.INIT1 = 16'h74b8;
    defparam add_989_15.INJECT1_0 = "NO";
    defparam add_989_15.INJECT1_1 = "NO";
    CCU2D add_989_13 (.A0(d2[46]), .B0(n4190), .C0(n4191[10]), .D0(d1[46]), 
          .A1(d2[47]), .B1(n4190), .C1(n4191[11]), .D1(d1[47]), .CIN(n12083), 
          .COUT(n12084), .S0(d2_71__N_489[46]), .S1(d2_71__N_489[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_989_13.INIT0 = 16'h74b8;
    defparam add_989_13.INIT1 = 16'h74b8;
    defparam add_989_13.INJECT1_0 = "NO";
    defparam add_989_13.INJECT1_1 = "NO";
    CCU2D add_989_11 (.A0(d2[44]), .B0(n4190), .C0(n4191[8]), .D0(d1[44]), 
          .A1(d2[45]), .B1(n4190), .C1(n4191[9]), .D1(d1[45]), .CIN(n12082), 
          .COUT(n12083), .S0(d2_71__N_489[44]), .S1(d2_71__N_489[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_989_11.INIT0 = 16'h74b8;
    defparam add_989_11.INIT1 = 16'h74b8;
    defparam add_989_11.INJECT1_0 = "NO";
    defparam add_989_11.INJECT1_1 = "NO";
    CCU2D add_989_9 (.A0(d2[42]), .B0(n4190), .C0(n4191[6]), .D0(d1[42]), 
          .A1(d2[43]), .B1(n4190), .C1(n4191[7]), .D1(d1[43]), .CIN(n12081), 
          .COUT(n12082), .S0(d2_71__N_489[42]), .S1(d2_71__N_489[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_989_9.INIT0 = 16'h74b8;
    defparam add_989_9.INIT1 = 16'h74b8;
    defparam add_989_9.INJECT1_0 = "NO";
    defparam add_989_9.INJECT1_1 = "NO";
    CCU2D add_989_7 (.A0(d2[40]), .B0(n4190), .C0(n4191[4]), .D0(d1[40]), 
          .A1(d2[41]), .B1(n4190), .C1(n4191[5]), .D1(d1[41]), .CIN(n12080), 
          .COUT(n12081), .S0(d2_71__N_489[40]), .S1(d2_71__N_489[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_989_7.INIT0 = 16'h74b8;
    defparam add_989_7.INIT1 = 16'h74b8;
    defparam add_989_7.INJECT1_0 = "NO";
    defparam add_989_7.INJECT1_1 = "NO";
    CCU2D add_989_5 (.A0(d2[38]), .B0(n4190), .C0(n4191[2]), .D0(d1[38]), 
          .A1(d2[39]), .B1(n4190), .C1(n4191[3]), .D1(d1[39]), .CIN(n12079), 
          .COUT(n12080), .S0(d2_71__N_489[38]), .S1(d2_71__N_489[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_989_5.INIT0 = 16'h74b8;
    defparam add_989_5.INIT1 = 16'h74b8;
    defparam add_989_5.INJECT1_0 = "NO";
    defparam add_989_5.INJECT1_1 = "NO";
    CCU2D add_989_3 (.A0(d2[36]), .B0(n4190), .C0(n4191[0]), .D0(d1[36]), 
          .A1(d2[37]), .B1(n4190), .C1(n4191[1]), .D1(d1[37]), .CIN(n12078), 
          .COUT(n12079), .S0(d2_71__N_489[36]), .S1(d2_71__N_489[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_989_3.INIT0 = 16'h74b8;
    defparam add_989_3.INIT1 = 16'h74b8;
    defparam add_989_3.INJECT1_0 = "NO";
    defparam add_989_3.INJECT1_1 = "NO";
    CCU2D add_989_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n4190), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n12078));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_989_1.INIT0 = 16'hF000;
    defparam add_989_1.INIT1 = 16'h0555;
    defparam add_989_1.INJECT1_0 = "NO";
    defparam add_989_1.INJECT1_1 = "NO";
    CCU2D add_993_36 (.A0(d2[70]), .B0(d3[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[71]), .B1(d3[71]), .C1(GND_net), .D1(GND_net), .CIN(n12073), 
          .S0(n4343[34]), .S1(n4343[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_993_36.INIT0 = 16'h5666;
    defparam add_993_36.INIT1 = 16'h5666;
    defparam add_993_36.INJECT1_0 = "NO";
    defparam add_993_36.INJECT1_1 = "NO";
    CCU2D add_993_34 (.A0(d2[68]), .B0(d3[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[69]), .B1(d3[69]), .C1(GND_net), .D1(GND_net), .CIN(n12072), 
          .COUT(n12073), .S0(n4343[32]), .S1(n4343[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_993_34.INIT0 = 16'h5666;
    defparam add_993_34.INIT1 = 16'h5666;
    defparam add_993_34.INJECT1_0 = "NO";
    defparam add_993_34.INJECT1_1 = "NO";
    FD1P3AX d_tmp_i0_i63 (.D(d5[63]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i63.GSR = "ENABLED";
    LUT4 shift_right_31_i206_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66_c), .D(n134), .Z(d_out_11__N_1818[5])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i206_3_lut_4_lut.init = 16'hfe10;
    FD1P3AX d_tmp_i0_i62 (.D(d5[62]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i62.GSR = "ENABLED";
    LUT4 i11_4_lut (.A(n21), .B(n19), .C(n15), .D(n16), .Z(n31)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(80[22:52])
    defparam i11_4_lut.init = 16'hfffe;
    FD1P3AX d_d_tmp_i0_i6 (.D(d_tmp[6]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i61 (.D(d5[61]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i60 (.D(d5[60]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i59 (.D(d5[59]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i58 (.D(d5[58]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i57 (.D(d5[57]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i56 (.D(d5[56]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i55 (.D(d5[55]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i54 (.D(d5[54]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i53 (.D(d5[53]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i52 (.D(d5[52]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i51 (.D(d5[51]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i50 (.D(d5[50]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i50.GSR = "ENABLED";
    LUT4 shift_right_31_i203_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63_c), .D(n131), .Z(d_out_11__N_1818[2])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i203_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i204_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64_c), .D(n132), .Z(d_out_11__N_1818[3])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i204_3_lut_4_lut.init = 16'hfe10;
    FD1P3AX d_tmp_i0_i49 (.D(d5[49]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i49.GSR = "ENABLED";
    CCU2D add_1034_35 (.A0(d_d6[68]), .B0(n5558), .C0(n5559[32]), .D0(d6[68]), 
          .A1(d_d6[69]), .B1(n5558), .C1(n5559[33]), .D1(d6[69]), .CIN(n11726), 
          .COUT(n11727), .S0(d7_71__N_1530[68]), .S1(d7_71__N_1530[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1034_35.INIT0 = 16'hb874;
    defparam add_1034_35.INIT1 = 16'hb874;
    defparam add_1034_35.INJECT1_0 = "NO";
    defparam add_1034_35.INJECT1_1 = "NO";
    FD1P3AX d_tmp_i0_i48 (.D(d5[48]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i47 (.D(d5[47]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i47.GSR = "ENABLED";
    CCU2D add_1034_27 (.A0(d_d6[60]), .B0(n5558), .C0(n5559[24]), .D0(d6[60]), 
          .A1(d_d6[61]), .B1(n5558), .C1(n5559[25]), .D1(d6[61]), .CIN(n11722), 
          .COUT(n11723), .S0(d7_71__N_1530[60]), .S1(d7_71__N_1530[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1034_27.INIT0 = 16'hb874;
    defparam add_1034_27.INIT1 = 16'hb874;
    defparam add_1034_27.INJECT1_0 = "NO";
    defparam add_1034_27.INJECT1_1 = "NO";
    CCU2D add_1034_25 (.A0(d_d6[58]), .B0(n5558), .C0(n5559[22]), .D0(d6[58]), 
          .A1(d_d6[59]), .B1(n5558), .C1(n5559[23]), .D1(d6[59]), .CIN(n11721), 
          .COUT(n11722), .S0(d7_71__N_1530[58]), .S1(d7_71__N_1530[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1034_25.INIT0 = 16'hb874;
    defparam add_1034_25.INIT1 = 16'hb874;
    defparam add_1034_25.INJECT1_0 = "NO";
    defparam add_1034_25.INJECT1_1 = "NO";
    CCU2D add_1034_23 (.A0(d_d6[56]), .B0(n5558), .C0(n5559[20]), .D0(d6[56]), 
          .A1(d_d6[57]), .B1(n5558), .C1(n5559[21]), .D1(d6[57]), .CIN(n11720), 
          .COUT(n11721), .S0(d7_71__N_1530[56]), .S1(d7_71__N_1530[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1034_23.INIT0 = 16'hb874;
    defparam add_1034_23.INIT1 = 16'hb874;
    defparam add_1034_23.INJECT1_0 = "NO";
    defparam add_1034_23.INJECT1_1 = "NO";
    CCU2D add_1034_21 (.A0(d_d6[54]), .B0(n5558), .C0(n5559[18]), .D0(d6[54]), 
          .A1(d_d6[55]), .B1(n5558), .C1(n5559[19]), .D1(d6[55]), .CIN(n11719), 
          .COUT(n11720), .S0(d7_71__N_1530[54]), .S1(d7_71__N_1530[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1034_21.INIT0 = 16'hb874;
    defparam add_1034_21.INIT1 = 16'hb874;
    defparam add_1034_21.INJECT1_0 = "NO";
    defparam add_1034_21.INJECT1_1 = "NO";
    FD1P3AX d_tmp_i0_i46 (.D(d5[46]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i46.GSR = "ENABLED";
    CCU2D add_1034_19 (.A0(d_d6[52]), .B0(n5558), .C0(n5559[16]), .D0(d6[52]), 
          .A1(d_d6[53]), .B1(n5558), .C1(n5559[17]), .D1(d6[53]), .CIN(n11718), 
          .COUT(n11719), .S0(d7_71__N_1530[52]), .S1(d7_71__N_1530[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1034_19.INIT0 = 16'hb874;
    defparam add_1034_19.INIT1 = 16'hb874;
    defparam add_1034_19.INJECT1_0 = "NO";
    defparam add_1034_19.INJECT1_1 = "NO";
    FD1P3AX d_tmp_i0_i45 (.D(d5[45]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i45.GSR = "ENABLED";
    CCU2D add_1034_17 (.A0(d_d6[50]), .B0(n5558), .C0(n5559[14]), .D0(d6[50]), 
          .A1(d_d6[51]), .B1(n5558), .C1(n5559[15]), .D1(d6[51]), .CIN(n11717), 
          .COUT(n11718), .S0(d7_71__N_1530[50]), .S1(d7_71__N_1530[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1034_17.INIT0 = 16'hb874;
    defparam add_1034_17.INIT1 = 16'hb874;
    defparam add_1034_17.INJECT1_0 = "NO";
    defparam add_1034_17.INJECT1_1 = "NO";
    CCU2D add_1034_15 (.A0(d_d6[48]), .B0(n5558), .C0(n5559[12]), .D0(d6[48]), 
          .A1(d_d6[49]), .B1(n5558), .C1(n5559[13]), .D1(d6[49]), .CIN(n11716), 
          .COUT(n11717), .S0(d7_71__N_1530[48]), .S1(d7_71__N_1530[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1034_15.INIT0 = 16'hb874;
    defparam add_1034_15.INIT1 = 16'hb874;
    defparam add_1034_15.INJECT1_0 = "NO";
    defparam add_1034_15.INJECT1_1 = "NO";
    CCU2D add_1034_13 (.A0(d_d6[46]), .B0(n5558), .C0(n5559[10]), .D0(d6[46]), 
          .A1(d_d6[47]), .B1(n5558), .C1(n5559[11]), .D1(d6[47]), .CIN(n11715), 
          .COUT(n11716), .S0(d7_71__N_1530[46]), .S1(d7_71__N_1530[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1034_13.INIT0 = 16'hb874;
    defparam add_1034_13.INIT1 = 16'hb874;
    defparam add_1034_13.INJECT1_0 = "NO";
    defparam add_1034_13.INJECT1_1 = "NO";
    CCU2D add_1034_11 (.A0(d_d6[44]), .B0(n5558), .C0(n5559[8]), .D0(d6[44]), 
          .A1(d_d6[45]), .B1(n5558), .C1(n5559[9]), .D1(d6[45]), .CIN(n11714), 
          .COUT(n11715), .S0(d7_71__N_1530[44]), .S1(d7_71__N_1530[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1034_11.INIT0 = 16'hb874;
    defparam add_1034_11.INIT1 = 16'hb874;
    defparam add_1034_11.INJECT1_0 = "NO";
    defparam add_1034_11.INJECT1_1 = "NO";
    CCU2D add_1034_9 (.A0(d_d6[42]), .B0(n5558), .C0(n5559[6]), .D0(d6[42]), 
          .A1(d_d6[43]), .B1(n5558), .C1(n5559[7]), .D1(d6[43]), .CIN(n11713), 
          .COUT(n11714), .S0(d7_71__N_1530[42]), .S1(d7_71__N_1530[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1034_9.INIT0 = 16'hb874;
    defparam add_1034_9.INIT1 = 16'hb874;
    defparam add_1034_9.INJECT1_0 = "NO";
    defparam add_1034_9.INJECT1_1 = "NO";
    CCU2D add_1034_7 (.A0(d_d6[40]), .B0(n5558), .C0(n5559[4]), .D0(d6[40]), 
          .A1(d_d6[41]), .B1(n5558), .C1(n5559[5]), .D1(d6[41]), .CIN(n11712), 
          .COUT(n11713), .S0(d7_71__N_1530[40]), .S1(d7_71__N_1530[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1034_7.INIT0 = 16'hb874;
    defparam add_1034_7.INIT1 = 16'hb874;
    defparam add_1034_7.INJECT1_0 = "NO";
    defparam add_1034_7.INJECT1_1 = "NO";
    CCU2D add_1034_5 (.A0(d_d6[38]), .B0(n5558), .C0(n5559[2]), .D0(d6[38]), 
          .A1(d_d6[39]), .B1(n5558), .C1(n5559[3]), .D1(d6[39]), .CIN(n11711), 
          .COUT(n11712), .S0(d7_71__N_1530[38]), .S1(d7_71__N_1530[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1034_5.INIT0 = 16'hb874;
    defparam add_1034_5.INIT1 = 16'hb874;
    defparam add_1034_5.INJECT1_0 = "NO";
    defparam add_1034_5.INJECT1_1 = "NO";
    CCU2D add_1034_3 (.A0(d_d6[36]), .B0(n5558), .C0(n5559[0]), .D0(d6[36]), 
          .A1(d_d6[37]), .B1(n5558), .C1(n5559[1]), .D1(d6[37]), .CIN(n11710), 
          .COUT(n11711), .S0(d7_71__N_1530[36]), .S1(d7_71__N_1530[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1034_3.INIT0 = 16'hb874;
    defparam add_1034_3.INIT1 = 16'hb874;
    defparam add_1034_3.INJECT1_0 = "NO";
    defparam add_1034_3.INJECT1_1 = "NO";
    CCU2D add_1034_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5558), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11710));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1034_1.INIT0 = 16'hF000;
    defparam add_1034_1.INIT1 = 16'h0555;
    defparam add_1034_1.INJECT1_0 = "NO";
    defparam add_1034_1.INJECT1_1 = "NO";
    CCU2D add_1038_37 (.A0(d7[71]), .B0(d_d7[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11706), 
          .S0(n5711[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1038_37.INIT0 = 16'h5999;
    defparam add_1038_37.INIT1 = 16'h0000;
    defparam add_1038_37.INJECT1_0 = "NO";
    defparam add_1038_37.INJECT1_1 = "NO";
    CCU2D add_1038_35 (.A0(d7[69]), .B0(d_d7[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[70]), .B1(d_d7[70]), .C1(GND_net), .D1(GND_net), .CIN(n11705), 
          .COUT(n11706), .S0(n5711[33]), .S1(n5711[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1038_35.INIT0 = 16'h5999;
    defparam add_1038_35.INIT1 = 16'h5999;
    defparam add_1038_35.INJECT1_0 = "NO";
    defparam add_1038_35.INJECT1_1 = "NO";
    CCU2D add_1038_33 (.A0(d7[67]), .B0(d_d7[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[68]), .B1(d_d7[68]), .C1(GND_net), .D1(GND_net), .CIN(n11704), 
          .COUT(n11705), .S0(n5711[31]), .S1(n5711[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1038_33.INIT0 = 16'h5999;
    defparam add_1038_33.INIT1 = 16'h5999;
    defparam add_1038_33.INJECT1_0 = "NO";
    defparam add_1038_33.INJECT1_1 = "NO";
    CCU2D add_1038_31 (.A0(d7[65]), .B0(d_d7[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[66]), .B1(d_d7[66]), .C1(GND_net), .D1(GND_net), .CIN(n11703), 
          .COUT(n11704), .S0(n5711[29]), .S1(n5711[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1038_31.INIT0 = 16'h5999;
    defparam add_1038_31.INIT1 = 16'h5999;
    defparam add_1038_31.INJECT1_0 = "NO";
    defparam add_1038_31.INJECT1_1 = "NO";
    CCU2D add_1038_29 (.A0(d7[63]), .B0(d_d7[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[64]), .B1(d_d7[64]), .C1(GND_net), .D1(GND_net), .CIN(n11702), 
          .COUT(n11703), .S0(n5711[27]), .S1(n5711[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1038_29.INIT0 = 16'h5999;
    defparam add_1038_29.INIT1 = 16'h5999;
    defparam add_1038_29.INJECT1_0 = "NO";
    defparam add_1038_29.INJECT1_1 = "NO";
    CCU2D add_1038_27 (.A0(d7[61]), .B0(d_d7[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[62]), .B1(d_d7[62]), .C1(GND_net), .D1(GND_net), .CIN(n11701), 
          .COUT(n11702), .S0(n5711[25]), .S1(n5711[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1038_27.INIT0 = 16'h5999;
    defparam add_1038_27.INIT1 = 16'h5999;
    defparam add_1038_27.INJECT1_0 = "NO";
    defparam add_1038_27.INJECT1_1 = "NO";
    CCU2D add_1038_25 (.A0(d7[59]), .B0(d_d7[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[60]), .B1(d_d7[60]), .C1(GND_net), .D1(GND_net), .CIN(n11700), 
          .COUT(n11701), .S0(n5711[23]), .S1(n5711[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1038_25.INIT0 = 16'h5999;
    defparam add_1038_25.INIT1 = 16'h5999;
    defparam add_1038_25.INJECT1_0 = "NO";
    defparam add_1038_25.INJECT1_1 = "NO";
    LUT4 i5805_4_lut (.A(count[9]), .B(count[2]), .C(count[7]), .D(count[1]), 
         .Z(n13254)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5805_4_lut.init = 16'h8000;
    CCU2D add_1038_23 (.A0(d7[57]), .B0(d_d7[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[58]), .B1(d_d7[58]), .C1(GND_net), .D1(GND_net), .CIN(n11699), 
          .COUT(n11700), .S0(n5711[21]), .S1(n5711[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1038_23.INIT0 = 16'h5999;
    defparam add_1038_23.INIT1 = 16'h5999;
    defparam add_1038_23.INJECT1_0 = "NO";
    defparam add_1038_23.INJECT1_1 = "NO";
    CCU2D add_1038_21 (.A0(d7[55]), .B0(d_d7[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[56]), .B1(d_d7[56]), .C1(GND_net), .D1(GND_net), .CIN(n11698), 
          .COUT(n11699), .S0(n5711[19]), .S1(n5711[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1038_21.INIT0 = 16'h5999;
    defparam add_1038_21.INIT1 = 16'h5999;
    defparam add_1038_21.INJECT1_0 = "NO";
    defparam add_1038_21.INJECT1_1 = "NO";
    CCU2D add_1038_19 (.A0(d7[53]), .B0(d_d7[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[54]), .B1(d_d7[54]), .C1(GND_net), .D1(GND_net), .CIN(n11697), 
          .COUT(n11698), .S0(n5711[17]), .S1(n5711[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1038_19.INIT0 = 16'h5999;
    defparam add_1038_19.INIT1 = 16'h5999;
    defparam add_1038_19.INJECT1_0 = "NO";
    defparam add_1038_19.INJECT1_1 = "NO";
    CCU2D add_993_32 (.A0(d2[66]), .B0(d3[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[67]), .B1(d3[67]), .C1(GND_net), .D1(GND_net), .CIN(n12071), 
          .COUT(n12072), .S0(n4343[30]), .S1(n4343[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_993_32.INIT0 = 16'h5666;
    defparam add_993_32.INIT1 = 16'h5666;
    defparam add_993_32.INJECT1_0 = "NO";
    defparam add_993_32.INJECT1_1 = "NO";
    FD1P3AX d_tmp_i0_i44 (.D(d5[44]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i44.GSR = "ENABLED";
    CCU2D add_1038_17 (.A0(d7[51]), .B0(d_d7[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[52]), .B1(d_d7[52]), .C1(GND_net), .D1(GND_net), .CIN(n11696), 
          .COUT(n11697), .S0(n5711[15]), .S1(n5711[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1038_17.INIT0 = 16'h5999;
    defparam add_1038_17.INIT1 = 16'h5999;
    defparam add_1038_17.INJECT1_0 = "NO";
    defparam add_1038_17.INJECT1_1 = "NO";
    LUT4 i7_4_lut (.A(count[10]), .B(count[1]), .C(count[5]), .D(count[6]), 
         .Z(n19)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(80[22:52])
    defparam i7_4_lut.init = 16'hfffe;
    FD1P3AX d_tmp_i0_i43 (.D(d5[43]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i42 (.D(d5[42]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i41 (.D(d5[41]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i40 (.D(d5[40]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i39 (.D(d5[39]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i38 (.D(d5[38]), .SP(osc_clk_enable_62), .CK(osc_clk), 
            .Q(d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i38.GSR = "ENABLED";
    CCU2D add_1038_15 (.A0(d7[49]), .B0(d_d7[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[50]), .B1(d_d7[50]), .C1(GND_net), .D1(GND_net), .CIN(n11695), 
          .COUT(n11696), .S0(n5711[13]), .S1(n5711[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1038_15.INIT0 = 16'h5999;
    defparam add_1038_15.INIT1 = 16'h5999;
    defparam add_1038_15.INJECT1_0 = "NO";
    defparam add_1038_15.INJECT1_1 = "NO";
    FD1P3AX d_tmp_i0_i37 (.D(d5[37]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i37.GSR = "ENABLED";
    LUT4 i3_2_lut (.A(count[8]), .B(count[7]), .Z(n15)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(80[22:52])
    defparam i3_2_lut.init = 16'heeee;
    CCU2D add_1038_13 (.A0(d7[47]), .B0(d_d7[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[48]), .B1(d_d7[48]), .C1(GND_net), .D1(GND_net), .CIN(n11694), 
          .COUT(n11695), .S0(n5711[11]), .S1(n5711[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1038_13.INIT0 = 16'h5999;
    defparam add_1038_13.INIT1 = 16'h5999;
    defparam add_1038_13.INJECT1_0 = "NO";
    defparam add_1038_13.INJECT1_1 = "NO";
    FD1P3AX d_tmp_i0_i36 (.D(d5[36]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i36.GSR = "ENABLED";
    CCU2D add_1038_11 (.A0(d7[45]), .B0(d_d7[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[46]), .B1(d_d7[46]), .C1(GND_net), .D1(GND_net), .CIN(n11693), 
          .COUT(n11694), .S0(n5711[9]), .S1(n5711[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1038_11.INIT0 = 16'h5999;
    defparam add_1038_11.INIT1 = 16'h5999;
    defparam add_1038_11.INJECT1_0 = "NO";
    defparam add_1038_11.INJECT1_1 = "NO";
    FD1P3AX d_tmp_i0_i35 (.D(d5[35]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i34 (.D(d5[34]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i33 (.D(d5[33]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i32 (.D(d5[32]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i31 (.D(d5[31]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i30 (.D(d5[30]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i30.GSR = "ENABLED";
    LUT4 i4_2_lut (.A(n12864), .B(count[2]), .Z(n16)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(80[22:52])
    defparam i4_2_lut.init = 16'heeee;
    CCU2D add_1038_9 (.A0(d7[43]), .B0(d_d7[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[44]), .B1(d_d7[44]), .C1(GND_net), .D1(GND_net), .CIN(n11692), 
          .COUT(n11693), .S0(n5711[7]), .S1(n5711[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1038_9.INIT0 = 16'h5999;
    defparam add_1038_9.INIT1 = 16'h5999;
    defparam add_1038_9.INJECT1_0 = "NO";
    defparam add_1038_9.INJECT1_1 = "NO";
    CCU2D add_1038_7 (.A0(d7[41]), .B0(d_d7[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[42]), .B1(d_d7[42]), .C1(GND_net), .D1(GND_net), .CIN(n11691), 
          .COUT(n11692), .S0(n5711[5]), .S1(n5711[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1038_7.INIT0 = 16'h5999;
    defparam add_1038_7.INIT1 = 16'h5999;
    defparam add_1038_7.INJECT1_0 = "NO";
    defparam add_1038_7.INJECT1_1 = "NO";
    FD1P3AX d_tmp_i0_i29 (.D(d5[29]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i28 (.D(d5[28]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i27 (.D(d5[27]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i26 (.D(d5[26]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i26.GSR = "ENABLED";
    LUT4 shift_right_31_i207_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n67_c), .D(n135), .Z(d_out_11__N_1818[6])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i207_3_lut_4_lut.init = 16'hfe10;
    FD1P3AX d_tmp_i0_i25 (.D(d5[25]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i24 (.D(d5[24]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i23 (.D(d5[23]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i22 (.D(d5[22]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i21 (.D(d5[21]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i20 (.D(d5[20]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i19 (.D(d5[19]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i18 (.D(d5[18]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i17 (.D(d5[17]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i16 (.D(d5[16]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i16.GSR = "ENABLED";
    CCU2D add_993_30 (.A0(d2[64]), .B0(d3[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[65]), .B1(d3[65]), .C1(GND_net), .D1(GND_net), .CIN(n12070), 
          .COUT(n12071), .S0(n4343[28]), .S1(n4343[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_993_30.INIT0 = 16'h5666;
    defparam add_993_30.INIT1 = 16'h5666;
    defparam add_993_30.INJECT1_0 = "NO";
    defparam add_993_30.INJECT1_1 = "NO";
    LUT4 i4815_2_lut (.A(d1[36]), .B(d2[36]), .Z(n4191[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4815_2_lut.init = 16'h6666;
    LUT4 shift_right_31_i61_3_lut (.A(d10[60]), .B(d10[61]), .C(\CICGain[0] ), 
         .Z(n61_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i61_3_lut.init = 16'hcaca;
    FD1P3AX d_tmp_i0_i15 (.D(d5[15]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i14 (.D(d5[14]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i13 (.D(d5[13]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i12 (.D(d5[12]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i11 (.D(d5[11]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i10 (.D(d5[10]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i9 (.D(d5[9]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i8 (.D(d5[8]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i8.GSR = "ENABLED";
    LUT4 i5855_4_lut_rep_195 (.A(n13252), .B(n13), .C(n13254), .D(n13238), 
         .Z(n14123)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i5855_4_lut_rep_195.init = 16'h2000;
    CCU2D add_982_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n12261), 
          .S0(n4038));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_982_cout.INIT0 = 16'h0000;
    defparam add_982_cout.INIT1 = 16'h0000;
    defparam add_982_cout.INJECT1_0 = "NO";
    defparam add_982_cout.INJECT1_1 = "NO";
    CCU2D add_1034_33 (.A0(d_d6[66]), .B0(n5558), .C0(n5559[30]), .D0(d6[66]), 
          .A1(d_d6[67]), .B1(n5558), .C1(n5559[31]), .D1(d6[67]), .CIN(n11725), 
          .COUT(n11726), .S0(d7_71__N_1530[66]), .S1(d7_71__N_1530[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1034_33.INIT0 = 16'hb874;
    defparam add_1034_33.INIT1 = 16'hb874;
    defparam add_1034_33.INJECT1_0 = "NO";
    defparam add_1034_33.INJECT1_1 = "NO";
    CCU2D add_982_36 (.A0(MixerOutSin[11]), .B0(d1[34]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[35]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12260), .COUT(n12261), .S0(d1_71__N_417[34]), 
          .S1(d1_71__N_417[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_982_36.INIT0 = 16'h5666;
    defparam add_982_36.INIT1 = 16'h5666;
    defparam add_982_36.INJECT1_0 = "NO";
    defparam add_982_36.INJECT1_1 = "NO";
    CCU2D add_982_34 (.A0(MixerOutSin[11]), .B0(d1[32]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[33]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12259), .COUT(n12260), .S0(d1_71__N_417[32]), 
          .S1(d1_71__N_417[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_982_34.INIT0 = 16'h5666;
    defparam add_982_34.INIT1 = 16'h5666;
    defparam add_982_34.INJECT1_0 = "NO";
    defparam add_982_34.INJECT1_1 = "NO";
    FD1P3AX d_tmp_i0_i7 (.D(d5[7]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i6 (.D(d5[6]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i5 (.D(d5[5]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i4 (.D(d5[4]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i3 (.D(d5[3]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i3.GSR = "ENABLED";
    LUT4 i4809_2_lut (.A(d3[36]), .B(d4[36]), .Z(n4495[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4809_2_lut.init = 16'h6666;
    FD1P3AX d_d_tmp_i0_i71 (.D(d_tmp[71]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i70 (.D(d_tmp[70]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i69 (.D(d_tmp[69]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i68 (.D(d_tmp[68]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i67 (.D(d_tmp[67]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i66 (.D(d_tmp[66]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i65 (.D(d_tmp[65]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i64 (.D(d_tmp[64]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i63 (.D(d_tmp[63]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i62 (.D(d_tmp[62]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i61 (.D(d_tmp[61]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i60 (.D(d_tmp[60]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i59 (.D(d_tmp[59]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i58 (.D(d_tmp[58]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i57 (.D(d_tmp[57]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i56 (.D(d_tmp[56]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i55 (.D(d_tmp[55]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i54 (.D(d_tmp[54]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i53 (.D(d_tmp[53]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i52 (.D(d_tmp[52]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i51 (.D(d_tmp[51]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i50 (.D(d_tmp[50]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i49 (.D(d_tmp[49]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i48 (.D(d_tmp[48]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i47 (.D(d_tmp[47]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i46 (.D(d_tmp[46]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i45 (.D(d_tmp[45]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i44 (.D(d_tmp[44]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i43 (.D(d_tmp[43]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i42 (.D(d_tmp[42]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i41 (.D(d_tmp[41]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i40 (.D(d_tmp[40]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i39 (.D(d_tmp[39]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i38 (.D(d_tmp[38]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i37 (.D(d_tmp[37]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i36 (.D(d_tmp[36]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i35 (.D(d_tmp[35]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i34 (.D(d_tmp[34]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i33 (.D(d_tmp[33]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i32 (.D(d_tmp[32]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i31 (.D(d_tmp[31]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i30 (.D(d_tmp[30]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i29 (.D(d_tmp[29]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i28 (.D(d_tmp[28]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i27 (.D(d_tmp[27]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i26 (.D(d_tmp[26]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i25 (.D(d_tmp[25]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i24 (.D(d_tmp[24]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i23 (.D(d_tmp[23]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i22 (.D(d_tmp[22]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i21 (.D(d_tmp[21]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i20 (.D(d_tmp[20]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i19 (.D(d_tmp[19]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i18 (.D(d_tmp[18]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i17 (.D(d_tmp[17]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i16 (.D(d_tmp[16]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i15 (.D(d_tmp[15]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i2 (.D(d5[2]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i2.GSR = "ENABLED";
    LUT4 shift_right_31_i208_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n68_c), .D(n136), .Z(d_out_11__N_1818[7])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i208_3_lut_4_lut.init = 16'hfe10;
    FD1P3AX d_d_tmp_i0_i14 (.D(d_tmp[14]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i13 (.D(d_tmp[13]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i12 (.D(d_tmp[12]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i11 (.D(d_tmp[11]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i10 (.D(d_tmp[10]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i10.GSR = "ENABLED";
    CCU2D add_1033_37 (.A0(d6[71]), .B0(d_d6[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11746), 
          .S0(n5559[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1033_37.INIT0 = 16'h5999;
    defparam add_1033_37.INIT1 = 16'h0000;
    defparam add_1033_37.INJECT1_0 = "NO";
    defparam add_1033_37.INJECT1_1 = "NO";
    CCU2D add_1033_35 (.A0(d6[69]), .B0(d_d6[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[70]), .B1(d_d6[70]), .C1(GND_net), .D1(GND_net), .CIN(n11745), 
          .COUT(n11746), .S0(n5559[33]), .S1(n5559[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1033_35.INIT0 = 16'h5999;
    defparam add_1033_35.INIT1 = 16'h5999;
    defparam add_1033_35.INJECT1_0 = "NO";
    defparam add_1033_35.INJECT1_1 = "NO";
    CCU2D add_1033_33 (.A0(d6[67]), .B0(d_d6[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[68]), .B1(d_d6[68]), .C1(GND_net), .D1(GND_net), .CIN(n11744), 
          .COUT(n11745), .S0(n5559[31]), .S1(n5559[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1033_33.INIT0 = 16'h5999;
    defparam add_1033_33.INIT1 = 16'h5999;
    defparam add_1033_33.INJECT1_0 = "NO";
    defparam add_1033_33.INJECT1_1 = "NO";
    CCU2D add_1033_31 (.A0(d6[65]), .B0(d_d6[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[66]), .B1(d_d6[66]), .C1(GND_net), .D1(GND_net), .CIN(n11743), 
          .COUT(n11744), .S0(n5559[29]), .S1(n5559[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1033_31.INIT0 = 16'h5999;
    defparam add_1033_31.INIT1 = 16'h5999;
    defparam add_1033_31.INJECT1_0 = "NO";
    defparam add_1033_31.INJECT1_1 = "NO";
    CCU2D add_1033_29 (.A0(d6[63]), .B0(d_d6[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[64]), .B1(d_d6[64]), .C1(GND_net), .D1(GND_net), .CIN(n11742), 
          .COUT(n11743), .S0(n5559[27]), .S1(n5559[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1033_29.INIT0 = 16'h5999;
    defparam add_1033_29.INIT1 = 16'h5999;
    defparam add_1033_29.INJECT1_0 = "NO";
    defparam add_1033_29.INJECT1_1 = "NO";
    CCU2D add_1033_27 (.A0(d6[61]), .B0(d_d6[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[62]), .B1(d_d6[62]), .C1(GND_net), .D1(GND_net), .CIN(n11741), 
          .COUT(n11742), .S0(n5559[25]), .S1(n5559[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1033_27.INIT0 = 16'h5999;
    defparam add_1033_27.INIT1 = 16'h5999;
    defparam add_1033_27.INJECT1_0 = "NO";
    defparam add_1033_27.INJECT1_1 = "NO";
    FD1P3AX d_d_tmp_i0_i9 (.D(d_tmp[9]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i9.GSR = "ENABLED";
    CCU2D add_1033_25 (.A0(d6[59]), .B0(d_d6[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[60]), .B1(d_d6[60]), .C1(GND_net), .D1(GND_net), .CIN(n11740), 
          .COUT(n11741), .S0(n5559[23]), .S1(n5559[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1033_25.INIT0 = 16'h5999;
    defparam add_1033_25.INIT1 = 16'h5999;
    defparam add_1033_25.INJECT1_0 = "NO";
    defparam add_1033_25.INJECT1_1 = "NO";
    CCU2D add_1033_23 (.A0(d6[57]), .B0(d_d6[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[58]), .B1(d_d6[58]), .C1(GND_net), .D1(GND_net), .CIN(n11739), 
          .COUT(n11740), .S0(n5559[21]), .S1(n5559[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1033_23.INIT0 = 16'h5999;
    defparam add_1033_23.INIT1 = 16'h5999;
    defparam add_1033_23.INJECT1_0 = "NO";
    defparam add_1033_23.INJECT1_1 = "NO";
    CCU2D add_1033_21 (.A0(d6[55]), .B0(d_d6[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[56]), .B1(d_d6[56]), .C1(GND_net), .D1(GND_net), .CIN(n11738), 
          .COUT(n11739), .S0(n5559[19]), .S1(n5559[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1033_21.INIT0 = 16'h5999;
    defparam add_1033_21.INIT1 = 16'h5999;
    defparam add_1033_21.INJECT1_0 = "NO";
    defparam add_1033_21.INJECT1_1 = "NO";
    FD1P3AX d_d_tmp_i0_i8 (.D(d_tmp[8]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i7 (.D(d_tmp[7]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d_d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i7.GSR = "ENABLED";
    CCU2D add_1033_19 (.A0(d6[53]), .B0(d_d6[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[54]), .B1(d_d6[54]), .C1(GND_net), .D1(GND_net), .CIN(n11737), 
          .COUT(n11738), .S0(n5559[17]), .S1(n5559[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1033_19.INIT0 = 16'h5999;
    defparam add_1033_19.INIT1 = 16'h5999;
    defparam add_1033_19.INJECT1_0 = "NO";
    defparam add_1033_19.INJECT1_1 = "NO";
    FD1P3AX d_tmp_i0_i1 (.D(d5[1]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i1.GSR = "ENABLED";
    CCU2D add_1033_17 (.A0(d6[51]), .B0(d_d6[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[52]), .B1(d_d6[52]), .C1(GND_net), .D1(GND_net), .CIN(n11736), 
          .COUT(n11737), .S0(n5559[15]), .S1(n5559[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1033_17.INIT0 = 16'h5999;
    defparam add_1033_17.INIT1 = 16'h5999;
    defparam add_1033_17.INJECT1_0 = "NO";
    defparam add_1033_17.INJECT1_1 = "NO";
    CCU2D add_1033_15 (.A0(d6[49]), .B0(d_d6[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[50]), .B1(d_d6[50]), .C1(GND_net), .D1(GND_net), .CIN(n11735), 
          .COUT(n11736), .S0(n5559[13]), .S1(n5559[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1033_15.INIT0 = 16'h5999;
    defparam add_1033_15.INIT1 = 16'h5999;
    defparam add_1033_15.INJECT1_0 = "NO";
    defparam add_1033_15.INJECT1_1 = "NO";
    LUT4 i11_3_lut_4_lut_then_3_lut (.A(\CICGain[0] ), .B(d10[67]), .C(d10[68]), 
         .Z(n13778)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam i11_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    CCU2D add_1033_13 (.A0(d6[47]), .B0(d_d6[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[48]), .B1(d_d6[48]), .C1(GND_net), .D1(GND_net), .CIN(n11734), 
          .COUT(n11735), .S0(n5559[11]), .S1(n5559[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1033_13.INIT0 = 16'h5999;
    defparam add_1033_13.INIT1 = 16'h5999;
    defparam add_1033_13.INJECT1_0 = "NO";
    defparam add_1033_13.INJECT1_1 = "NO";
    CCU2D add_1033_11 (.A0(d6[45]), .B0(d_d6[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[46]), .B1(d_d6[46]), .C1(GND_net), .D1(GND_net), .CIN(n11733), 
          .COUT(n11734), .S0(n5559[9]), .S1(n5559[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1033_11.INIT0 = 16'h5999;
    defparam add_1033_11.INIT1 = 16'h5999;
    defparam add_1033_11.INJECT1_0 = "NO";
    defparam add_1033_11.INJECT1_1 = "NO";
    CCU2D add_1033_9 (.A0(d6[43]), .B0(d_d6[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[44]), .B1(d_d6[44]), .C1(GND_net), .D1(GND_net), .CIN(n11732), 
          .COUT(n11733), .S0(n5559[7]), .S1(n5559[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1033_9.INIT0 = 16'h5999;
    defparam add_1033_9.INIT1 = 16'h5999;
    defparam add_1033_9.INJECT1_0 = "NO";
    defparam add_1033_9.INJECT1_1 = "NO";
    CCU2D add_1033_7 (.A0(d6[41]), .B0(d_d6[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[42]), .B1(d_d6[42]), .C1(GND_net), .D1(GND_net), .CIN(n11731), 
          .COUT(n11732), .S0(n5559[5]), .S1(n5559[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1033_7.INIT0 = 16'h5999;
    defparam add_1033_7.INIT1 = 16'h5999;
    defparam add_1033_7.INJECT1_0 = "NO";
    defparam add_1033_7.INJECT1_1 = "NO";
    CCU2D add_1033_5 (.A0(d6[39]), .B0(d_d6[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[40]), .B1(d_d6[40]), .C1(GND_net), .D1(GND_net), .CIN(n11730), 
          .COUT(n11731), .S0(n5559[3]), .S1(n5559[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1033_5.INIT0 = 16'h5999;
    defparam add_1033_5.INIT1 = 16'h5999;
    defparam add_1033_5.INJECT1_0 = "NO";
    defparam add_1033_5.INJECT1_1 = "NO";
    CCU2D add_1033_3 (.A0(d6[37]), .B0(d_d6[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[38]), .B1(d_d6[38]), .C1(GND_net), .D1(GND_net), .CIN(n11729), 
          .COUT(n11730), .S0(n5559[1]), .S1(n5559[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1033_3.INIT0 = 16'h5999;
    defparam add_1033_3.INIT1 = 16'h5999;
    defparam add_1033_3.INJECT1_0 = "NO";
    defparam add_1033_3.INJECT1_1 = "NO";
    CCU2D add_1033_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d6[36]), .B1(d_d6[36]), .C1(GND_net), .D1(GND_net), .COUT(n11729), 
          .S1(n5559[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1033_1.INIT0 = 16'hF000;
    defparam add_1033_1.INIT1 = 16'h5999;
    defparam add_1033_1.INJECT1_0 = "NO";
    defparam add_1033_1.INJECT1_1 = "NO";
    FD1P3AX d_tmp_i0_i0 (.D(d5[0]), .SP(d_clk_tmp_N_1830), .CK(osc_clk), 
            .Q(d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i0.GSR = "ENABLED";
    FD1S3AX d2_i1 (.D(d2_71__N_489[1]), .CK(osc_clk), .Q(d2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i1.GSR = "ENABLED";
    CCU2D add_993_28 (.A0(d2[62]), .B0(d3[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[63]), .B1(d3[63]), .C1(GND_net), .D1(GND_net), .CIN(n12069), 
          .COUT(n12070), .S0(n4343[26]), .S1(n4343[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_993_28.INIT0 = 16'h5666;
    defparam add_993_28.INIT1 = 16'h5666;
    defparam add_993_28.INJECT1_0 = "NO";
    defparam add_993_28.INJECT1_1 = "NO";
    CCU2D add_993_26 (.A0(d2[60]), .B0(d3[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[61]), .B1(d3[61]), .C1(GND_net), .D1(GND_net), .CIN(n12068), 
          .COUT(n12069), .S0(n4343[24]), .S1(n4343[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_993_26.INIT0 = 16'h5666;
    defparam add_993_26.INIT1 = 16'h5666;
    defparam add_993_26.INJECT1_0 = "NO";
    defparam add_993_26.INJECT1_1 = "NO";
    CCU2D add_993_24 (.A0(d2[58]), .B0(d3[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[59]), .B1(d3[59]), .C1(GND_net), .D1(GND_net), .CIN(n12067), 
          .COUT(n12068), .S0(n4343[22]), .S1(n4343[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_993_24.INIT0 = 16'h5666;
    defparam add_993_24.INIT1 = 16'h5666;
    defparam add_993_24.INJECT1_0 = "NO";
    defparam add_993_24.INJECT1_1 = "NO";
    CCU2D add_993_22 (.A0(d2[56]), .B0(d3[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[57]), .B1(d3[57]), .C1(GND_net), .D1(GND_net), .CIN(n12066), 
          .COUT(n12067), .S0(n4343[20]), .S1(n4343[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_993_22.INIT0 = 16'h5666;
    defparam add_993_22.INIT1 = 16'h5666;
    defparam add_993_22.INJECT1_0 = "NO";
    defparam add_993_22.INJECT1_1 = "NO";
    CCU2D add_993_20 (.A0(d2[54]), .B0(d3[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[55]), .B1(d3[55]), .C1(GND_net), .D1(GND_net), .CIN(n12065), 
          .COUT(n12066), .S0(n4343[18]), .S1(n4343[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_993_20.INIT0 = 16'h5666;
    defparam add_993_20.INIT1 = 16'h5666;
    defparam add_993_20.INJECT1_0 = "NO";
    defparam add_993_20.INJECT1_1 = "NO";
    CCU2D add_993_18 (.A0(d2[52]), .B0(d3[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[53]), .B1(d3[53]), .C1(GND_net), .D1(GND_net), .CIN(n12064), 
          .COUT(n12065), .S0(n4343[16]), .S1(n4343[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_993_18.INIT0 = 16'h5666;
    defparam add_993_18.INIT1 = 16'h5666;
    defparam add_993_18.INJECT1_0 = "NO";
    defparam add_993_18.INJECT1_1 = "NO";
    CCU2D add_993_16 (.A0(d2[50]), .B0(d3[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[51]), .B1(d3[51]), .C1(GND_net), .D1(GND_net), .CIN(n12063), 
          .COUT(n12064), .S0(n4343[14]), .S1(n4343[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_993_16.INIT0 = 16'h5666;
    defparam add_993_16.INIT1 = 16'h5666;
    defparam add_993_16.INJECT1_0 = "NO";
    defparam add_993_16.INJECT1_1 = "NO";
    CCU2D add_993_14 (.A0(d2[48]), .B0(d3[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[49]), .B1(d3[49]), .C1(GND_net), .D1(GND_net), .CIN(n12062), 
          .COUT(n12063), .S0(n4343[12]), .S1(n4343[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_993_14.INIT0 = 16'h5666;
    defparam add_993_14.INIT1 = 16'h5666;
    defparam add_993_14.INJECT1_0 = "NO";
    defparam add_993_14.INJECT1_1 = "NO";
    CCU2D add_993_12 (.A0(d2[46]), .B0(d3[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[47]), .B1(d3[47]), .C1(GND_net), .D1(GND_net), .CIN(n12061), 
          .COUT(n12062), .S0(n4343[10]), .S1(n4343[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_993_12.INIT0 = 16'h5666;
    defparam add_993_12.INIT1 = 16'h5666;
    defparam add_993_12.INJECT1_0 = "NO";
    defparam add_993_12.INJECT1_1 = "NO";
    CCU2D add_993_10 (.A0(d2[44]), .B0(d3[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[45]), .B1(d3[45]), .C1(GND_net), .D1(GND_net), .CIN(n12060), 
          .COUT(n12061), .S0(n4343[8]), .S1(n4343[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_993_10.INIT0 = 16'h5666;
    defparam add_993_10.INIT1 = 16'h5666;
    defparam add_993_10.INJECT1_0 = "NO";
    defparam add_993_10.INJECT1_1 = "NO";
    CCU2D add_993_8 (.A0(d2[42]), .B0(d3[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[43]), .B1(d3[43]), .C1(GND_net), .D1(GND_net), .CIN(n12059), 
          .COUT(n12060), .S0(n4343[6]), .S1(n4343[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_993_8.INIT0 = 16'h5666;
    defparam add_993_8.INIT1 = 16'h5666;
    defparam add_993_8.INJECT1_0 = "NO";
    defparam add_993_8.INJECT1_1 = "NO";
    CCU2D add_993_6 (.A0(d2[40]), .B0(d3[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[41]), .B1(d3[41]), .C1(GND_net), .D1(GND_net), .CIN(n12058), 
          .COUT(n12059), .S0(n4343[4]), .S1(n4343[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_993_6.INIT0 = 16'h5666;
    defparam add_993_6.INIT1 = 16'h5666;
    defparam add_993_6.INJECT1_0 = "NO";
    defparam add_993_6.INJECT1_1 = "NO";
    CCU2D add_993_4 (.A0(d2[38]), .B0(d3[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[39]), .B1(d3[39]), .C1(GND_net), .D1(GND_net), .CIN(n12057), 
          .COUT(n12058), .S0(n4343[2]), .S1(n4343[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_993_4.INIT0 = 16'h5666;
    defparam add_993_4.INIT1 = 16'h5666;
    defparam add_993_4.INJECT1_0 = "NO";
    defparam add_993_4.INJECT1_1 = "NO";
    CCU2D add_993_2 (.A0(d2[36]), .B0(d3[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[37]), .B1(d3[37]), .C1(GND_net), .D1(GND_net), .COUT(n12057), 
          .S1(n4343[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_993_2.INIT0 = 16'h7000;
    defparam add_993_2.INIT1 = 16'h5666;
    defparam add_993_2.INJECT1_0 = "NO";
    defparam add_993_2.INJECT1_1 = "NO";
    FD1S3AX d2_i2 (.D(d2_71__N_489[2]), .CK(osc_clk), .Q(d2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i2.GSR = "ENABLED";
    FD1S3AX d2_i3 (.D(d2_71__N_489[3]), .CK(osc_clk), .Q(d2[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i3.GSR = "ENABLED";
    FD1S3AX d2_i4 (.D(d2_71__N_489[4]), .CK(osc_clk), .Q(d2[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i4.GSR = "ENABLED";
    FD1S3AX d2_i5 (.D(d2_71__N_489[5]), .CK(osc_clk), .Q(d2[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i5.GSR = "ENABLED";
    FD1S3AX d2_i6 (.D(d2_71__N_489[6]), .CK(osc_clk), .Q(d2[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i6.GSR = "ENABLED";
    FD1S3AX d2_i7 (.D(d2_71__N_489[7]), .CK(osc_clk), .Q(d2[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i7.GSR = "ENABLED";
    FD1S3AX d2_i8 (.D(d2_71__N_489[8]), .CK(osc_clk), .Q(d2[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i8.GSR = "ENABLED";
    FD1S3AX d2_i9 (.D(d2_71__N_489[9]), .CK(osc_clk), .Q(d2[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i9.GSR = "ENABLED";
    FD1S3AX d2_i10 (.D(d2_71__N_489[10]), .CK(osc_clk), .Q(d2[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i10.GSR = "ENABLED";
    FD1S3AX d2_i11 (.D(d2_71__N_489[11]), .CK(osc_clk), .Q(d2[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i11.GSR = "ENABLED";
    FD1S3AX d2_i12 (.D(d2_71__N_489[12]), .CK(osc_clk), .Q(d2[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i12.GSR = "ENABLED";
    FD1S3AX d2_i13 (.D(d2_71__N_489[13]), .CK(osc_clk), .Q(d2[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i13.GSR = "ENABLED";
    FD1S3AX d2_i14 (.D(d2_71__N_489[14]), .CK(osc_clk), .Q(d2[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i14.GSR = "ENABLED";
    FD1S3AX d2_i15 (.D(d2_71__N_489[15]), .CK(osc_clk), .Q(d2[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i15.GSR = "ENABLED";
    FD1S3AX d2_i16 (.D(d2_71__N_489[16]), .CK(osc_clk), .Q(d2[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i16.GSR = "ENABLED";
    FD1S3AX d2_i17 (.D(d2_71__N_489[17]), .CK(osc_clk), .Q(d2[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i17.GSR = "ENABLED";
    FD1S3AX d2_i18 (.D(d2_71__N_489[18]), .CK(osc_clk), .Q(d2[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i18.GSR = "ENABLED";
    FD1S3AX d2_i19 (.D(d2_71__N_489[19]), .CK(osc_clk), .Q(d2[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i19.GSR = "ENABLED";
    FD1S3AX d2_i20 (.D(d2_71__N_489[20]), .CK(osc_clk), .Q(d2[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i20.GSR = "ENABLED";
    FD1S3AX d2_i21 (.D(d2_71__N_489[21]), .CK(osc_clk), .Q(d2[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i21.GSR = "ENABLED";
    FD1S3AX d2_i22 (.D(d2_71__N_489[22]), .CK(osc_clk), .Q(d2[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i22.GSR = "ENABLED";
    FD1S3AX d2_i23 (.D(d2_71__N_489[23]), .CK(osc_clk), .Q(d2[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i23.GSR = "ENABLED";
    FD1S3AX d2_i24 (.D(d2_71__N_489[24]), .CK(osc_clk), .Q(d2[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i24.GSR = "ENABLED";
    FD1S3AX d2_i25 (.D(d2_71__N_489[25]), .CK(osc_clk), .Q(d2[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i25.GSR = "ENABLED";
    FD1S3AX d2_i26 (.D(d2_71__N_489[26]), .CK(osc_clk), .Q(d2[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i26.GSR = "ENABLED";
    FD1S3AX d2_i27 (.D(d2_71__N_489[27]), .CK(osc_clk), .Q(d2[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i27.GSR = "ENABLED";
    FD1S3AX d2_i28 (.D(d2_71__N_489[28]), .CK(osc_clk), .Q(d2[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i28.GSR = "ENABLED";
    FD1S3AX d2_i29 (.D(d2_71__N_489[29]), .CK(osc_clk), .Q(d2[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i29.GSR = "ENABLED";
    FD1S3AX d2_i30 (.D(d2_71__N_489[30]), .CK(osc_clk), .Q(d2[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i30.GSR = "ENABLED";
    FD1S3AX d2_i31 (.D(d2_71__N_489[31]), .CK(osc_clk), .Q(d2[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i31.GSR = "ENABLED";
    FD1S3AX d2_i32 (.D(d2_71__N_489[32]), .CK(osc_clk), .Q(d2[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i32.GSR = "ENABLED";
    FD1S3AX d2_i33 (.D(d2_71__N_489[33]), .CK(osc_clk), .Q(d2[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i33.GSR = "ENABLED";
    FD1S3AX d2_i34 (.D(d2_71__N_489[34]), .CK(osc_clk), .Q(d2[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i34.GSR = "ENABLED";
    FD1S3AX d2_i35 (.D(d2_71__N_489[35]), .CK(osc_clk), .Q(d2[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i35.GSR = "ENABLED";
    FD1S3AX d2_i36 (.D(d2_71__N_489[36]), .CK(osc_clk), .Q(d2[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i36.GSR = "ENABLED";
    FD1S3AX d2_i37 (.D(d2_71__N_489[37]), .CK(osc_clk), .Q(d2[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i37.GSR = "ENABLED";
    FD1S3AX d2_i38 (.D(d2_71__N_489[38]), .CK(osc_clk), .Q(d2[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i38.GSR = "ENABLED";
    FD1S3AX d2_i39 (.D(d2_71__N_489[39]), .CK(osc_clk), .Q(d2[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i39.GSR = "ENABLED";
    FD1S3AX d2_i40 (.D(d2_71__N_489[40]), .CK(osc_clk), .Q(d2[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i40.GSR = "ENABLED";
    FD1S3AX d2_i41 (.D(d2_71__N_489[41]), .CK(osc_clk), .Q(d2[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i41.GSR = "ENABLED";
    FD1S3AX d2_i42 (.D(d2_71__N_489[42]), .CK(osc_clk), .Q(d2[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i42.GSR = "ENABLED";
    FD1S3AX d2_i43 (.D(d2_71__N_489[43]), .CK(osc_clk), .Q(d2[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i43.GSR = "ENABLED";
    FD1S3AX d2_i44 (.D(d2_71__N_489[44]), .CK(osc_clk), .Q(d2[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i44.GSR = "ENABLED";
    FD1S3AX d2_i45 (.D(d2_71__N_489[45]), .CK(osc_clk), .Q(d2[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i45.GSR = "ENABLED";
    FD1S3AX d2_i46 (.D(d2_71__N_489[46]), .CK(osc_clk), .Q(d2[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i46.GSR = "ENABLED";
    FD1S3AX d2_i47 (.D(d2_71__N_489[47]), .CK(osc_clk), .Q(d2[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i47.GSR = "ENABLED";
    FD1S3AX d2_i48 (.D(d2_71__N_489[48]), .CK(osc_clk), .Q(d2[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i48.GSR = "ENABLED";
    FD1S3AX d2_i49 (.D(d2_71__N_489[49]), .CK(osc_clk), .Q(d2[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i49.GSR = "ENABLED";
    FD1S3AX d2_i50 (.D(d2_71__N_489[50]), .CK(osc_clk), .Q(d2[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i50.GSR = "ENABLED";
    FD1S3AX d2_i51 (.D(d2_71__N_489[51]), .CK(osc_clk), .Q(d2[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i51.GSR = "ENABLED";
    FD1S3AX d2_i52 (.D(d2_71__N_489[52]), .CK(osc_clk), .Q(d2[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i52.GSR = "ENABLED";
    FD1S3AX d2_i53 (.D(d2_71__N_489[53]), .CK(osc_clk), .Q(d2[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i53.GSR = "ENABLED";
    FD1S3AX d2_i54 (.D(d2_71__N_489[54]), .CK(osc_clk), .Q(d2[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i54.GSR = "ENABLED";
    FD1S3AX d2_i55 (.D(d2_71__N_489[55]), .CK(osc_clk), .Q(d2[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i55.GSR = "ENABLED";
    FD1S3AX d2_i56 (.D(d2_71__N_489[56]), .CK(osc_clk), .Q(d2[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i56.GSR = "ENABLED";
    FD1S3AX d2_i57 (.D(d2_71__N_489[57]), .CK(osc_clk), .Q(d2[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i57.GSR = "ENABLED";
    FD1S3AX d2_i58 (.D(d2_71__N_489[58]), .CK(osc_clk), .Q(d2[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i58.GSR = "ENABLED";
    FD1S3AX d2_i59 (.D(d2_71__N_489[59]), .CK(osc_clk), .Q(d2[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i59.GSR = "ENABLED";
    FD1S3AX d2_i60 (.D(d2_71__N_489[60]), .CK(osc_clk), .Q(d2[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i60.GSR = "ENABLED";
    FD1S3AX d2_i61 (.D(d2_71__N_489[61]), .CK(osc_clk), .Q(d2[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i61.GSR = "ENABLED";
    FD1S3AX d2_i62 (.D(d2_71__N_489[62]), .CK(osc_clk), .Q(d2[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i62.GSR = "ENABLED";
    FD1S3AX d2_i63 (.D(d2_71__N_489[63]), .CK(osc_clk), .Q(d2[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i63.GSR = "ENABLED";
    FD1S3AX d2_i64 (.D(d2_71__N_489[64]), .CK(osc_clk), .Q(d2[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i64.GSR = "ENABLED";
    FD1S3AX d2_i65 (.D(d2_71__N_489[65]), .CK(osc_clk), .Q(d2[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i65.GSR = "ENABLED";
    FD1S3AX d2_i66 (.D(d2_71__N_489[66]), .CK(osc_clk), .Q(d2[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i66.GSR = "ENABLED";
    FD1S3AX d2_i67 (.D(d2_71__N_489[67]), .CK(osc_clk), .Q(d2[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i67.GSR = "ENABLED";
    FD1S3AX d2_i68 (.D(d2_71__N_489[68]), .CK(osc_clk), .Q(d2[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i68.GSR = "ENABLED";
    FD1S3AX d2_i69 (.D(d2_71__N_489[69]), .CK(osc_clk), .Q(d2[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i69.GSR = "ENABLED";
    FD1S3AX d2_i70 (.D(d2_71__N_489[70]), .CK(osc_clk), .Q(d2[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i70.GSR = "ENABLED";
    FD1S3AX d2_i71 (.D(d2_71__N_489[71]), .CK(osc_clk), .Q(d2[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i71.GSR = "ENABLED";
    FD1S3AX d3_i1 (.D(d3_71__N_561[1]), .CK(osc_clk), .Q(d3[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i1.GSR = "ENABLED";
    FD1S3AX d3_i2 (.D(d3_71__N_561[2]), .CK(osc_clk), .Q(d3[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i2.GSR = "ENABLED";
    FD1S3AX d3_i3 (.D(d3_71__N_561[3]), .CK(osc_clk), .Q(d3[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i3.GSR = "ENABLED";
    FD1S3AX d3_i4 (.D(d3_71__N_561[4]), .CK(osc_clk), .Q(d3[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i4.GSR = "ENABLED";
    FD1S3AX d3_i5 (.D(d3_71__N_561[5]), .CK(osc_clk), .Q(d3[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i5.GSR = "ENABLED";
    FD1S3AX d3_i6 (.D(d3_71__N_561[6]), .CK(osc_clk), .Q(d3[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i6.GSR = "ENABLED";
    FD1S3AX d3_i7 (.D(d3_71__N_561[7]), .CK(osc_clk), .Q(d3[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i7.GSR = "ENABLED";
    FD1S3AX d3_i8 (.D(d3_71__N_561[8]), .CK(osc_clk), .Q(d3[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i8.GSR = "ENABLED";
    FD1S3AX d3_i9 (.D(d3_71__N_561[9]), .CK(osc_clk), .Q(d3[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i9.GSR = "ENABLED";
    FD1S3AX d3_i10 (.D(d3_71__N_561[10]), .CK(osc_clk), .Q(d3[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i10.GSR = "ENABLED";
    FD1S3AX d3_i11 (.D(d3_71__N_561[11]), .CK(osc_clk), .Q(d3[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i11.GSR = "ENABLED";
    FD1S3AX d3_i12 (.D(d3_71__N_561[12]), .CK(osc_clk), .Q(d3[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i12.GSR = "ENABLED";
    FD1S3AX d3_i13 (.D(d3_71__N_561[13]), .CK(osc_clk), .Q(d3[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i13.GSR = "ENABLED";
    FD1S3AX d3_i14 (.D(d3_71__N_561[14]), .CK(osc_clk), .Q(d3[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i14.GSR = "ENABLED";
    FD1S3AX d3_i15 (.D(d3_71__N_561[15]), .CK(osc_clk), .Q(d3[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i15.GSR = "ENABLED";
    FD1S3AX d3_i16 (.D(d3_71__N_561[16]), .CK(osc_clk), .Q(d3[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i16.GSR = "ENABLED";
    FD1S3AX d3_i17 (.D(d3_71__N_561[17]), .CK(osc_clk), .Q(d3[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i17.GSR = "ENABLED";
    FD1S3AX d3_i18 (.D(d3_71__N_561[18]), .CK(osc_clk), .Q(d3[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i18.GSR = "ENABLED";
    FD1S3AX d3_i19 (.D(d3_71__N_561[19]), .CK(osc_clk), .Q(d3[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i19.GSR = "ENABLED";
    FD1S3AX d3_i20 (.D(d3_71__N_561[20]), .CK(osc_clk), .Q(d3[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i20.GSR = "ENABLED";
    FD1S3AX d3_i21 (.D(d3_71__N_561[21]), .CK(osc_clk), .Q(d3[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i21.GSR = "ENABLED";
    FD1S3AX d3_i22 (.D(d3_71__N_561[22]), .CK(osc_clk), .Q(d3[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i22.GSR = "ENABLED";
    FD1S3AX d3_i23 (.D(d3_71__N_561[23]), .CK(osc_clk), .Q(d3[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i23.GSR = "ENABLED";
    FD1S3AX d3_i24 (.D(d3_71__N_561[24]), .CK(osc_clk), .Q(d3[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i24.GSR = "ENABLED";
    FD1S3AX d3_i25 (.D(d3_71__N_561[25]), .CK(osc_clk), .Q(d3[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i25.GSR = "ENABLED";
    FD1S3AX d3_i26 (.D(d3_71__N_561[26]), .CK(osc_clk), .Q(d3[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i26.GSR = "ENABLED";
    FD1S3AX d3_i27 (.D(d3_71__N_561[27]), .CK(osc_clk), .Q(d3[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i27.GSR = "ENABLED";
    FD1S3AX d3_i28 (.D(d3_71__N_561[28]), .CK(osc_clk), .Q(d3[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i28.GSR = "ENABLED";
    FD1S3AX d3_i29 (.D(d3_71__N_561[29]), .CK(osc_clk), .Q(d3[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i29.GSR = "ENABLED";
    FD1S3AX d3_i30 (.D(d3_71__N_561[30]), .CK(osc_clk), .Q(d3[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i30.GSR = "ENABLED";
    FD1S3AX d3_i31 (.D(d3_71__N_561[31]), .CK(osc_clk), .Q(d3[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i31.GSR = "ENABLED";
    FD1S3AX d3_i32 (.D(d3_71__N_561[32]), .CK(osc_clk), .Q(d3[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i32.GSR = "ENABLED";
    FD1S3AX d3_i33 (.D(d3_71__N_561[33]), .CK(osc_clk), .Q(d3[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i33.GSR = "ENABLED";
    FD1S3AX d3_i34 (.D(d3_71__N_561[34]), .CK(osc_clk), .Q(d3[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i34.GSR = "ENABLED";
    FD1S3AX d3_i35 (.D(d3_71__N_561[35]), .CK(osc_clk), .Q(d3[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i35.GSR = "ENABLED";
    FD1S3AX d3_i36 (.D(d3_71__N_561[36]), .CK(osc_clk), .Q(d3[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i36.GSR = "ENABLED";
    FD1S3AX d3_i37 (.D(d3_71__N_561[37]), .CK(osc_clk), .Q(d3[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i37.GSR = "ENABLED";
    FD1S3AX d3_i38 (.D(d3_71__N_561[38]), .CK(osc_clk), .Q(d3[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i38.GSR = "ENABLED";
    FD1S3AX d3_i39 (.D(d3_71__N_561[39]), .CK(osc_clk), .Q(d3[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i39.GSR = "ENABLED";
    FD1S3AX d3_i40 (.D(d3_71__N_561[40]), .CK(osc_clk), .Q(d3[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i40.GSR = "ENABLED";
    FD1S3AX d3_i41 (.D(d3_71__N_561[41]), .CK(osc_clk), .Q(d3[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i41.GSR = "ENABLED";
    FD1S3AX d3_i42 (.D(d3_71__N_561[42]), .CK(osc_clk), .Q(d3[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i42.GSR = "ENABLED";
    FD1S3AX d3_i43 (.D(d3_71__N_561[43]), .CK(osc_clk), .Q(d3[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i43.GSR = "ENABLED";
    FD1S3AX d3_i44 (.D(d3_71__N_561[44]), .CK(osc_clk), .Q(d3[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i44.GSR = "ENABLED";
    FD1S3AX d3_i45 (.D(d3_71__N_561[45]), .CK(osc_clk), .Q(d3[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i45.GSR = "ENABLED";
    FD1S3AX d3_i46 (.D(d3_71__N_561[46]), .CK(osc_clk), .Q(d3[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i46.GSR = "ENABLED";
    FD1S3AX d3_i47 (.D(d3_71__N_561[47]), .CK(osc_clk), .Q(d3[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i47.GSR = "ENABLED";
    FD1S3AX d3_i48 (.D(d3_71__N_561[48]), .CK(osc_clk), .Q(d3[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i48.GSR = "ENABLED";
    FD1S3AX d3_i49 (.D(d3_71__N_561[49]), .CK(osc_clk), .Q(d3[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i49.GSR = "ENABLED";
    FD1S3AX d3_i50 (.D(d3_71__N_561[50]), .CK(osc_clk), .Q(d3[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i50.GSR = "ENABLED";
    FD1S3AX d3_i51 (.D(d3_71__N_561[51]), .CK(osc_clk), .Q(d3[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i51.GSR = "ENABLED";
    FD1S3AX d3_i52 (.D(d3_71__N_561[52]), .CK(osc_clk), .Q(d3[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i52.GSR = "ENABLED";
    FD1S3AX d3_i53 (.D(d3_71__N_561[53]), .CK(osc_clk), .Q(d3[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i53.GSR = "ENABLED";
    FD1S3AX d3_i54 (.D(d3_71__N_561[54]), .CK(osc_clk), .Q(d3[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i54.GSR = "ENABLED";
    FD1S3AX d3_i55 (.D(d3_71__N_561[55]), .CK(osc_clk), .Q(d3[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i55.GSR = "ENABLED";
    FD1S3AX d3_i56 (.D(d3_71__N_561[56]), .CK(osc_clk), .Q(d3[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i56.GSR = "ENABLED";
    FD1S3AX d3_i57 (.D(d3_71__N_561[57]), .CK(osc_clk), .Q(d3[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i57.GSR = "ENABLED";
    FD1S3AX d3_i58 (.D(d3_71__N_561[58]), .CK(osc_clk), .Q(d3[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i58.GSR = "ENABLED";
    FD1S3AX d3_i59 (.D(d3_71__N_561[59]), .CK(osc_clk), .Q(d3[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i59.GSR = "ENABLED";
    FD1S3AX d3_i60 (.D(d3_71__N_561[60]), .CK(osc_clk), .Q(d3[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i60.GSR = "ENABLED";
    FD1S3AX d3_i61 (.D(d3_71__N_561[61]), .CK(osc_clk), .Q(d3[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i61.GSR = "ENABLED";
    FD1S3AX d3_i62 (.D(d3_71__N_561[62]), .CK(osc_clk), .Q(d3[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i62.GSR = "ENABLED";
    FD1S3AX d3_i63 (.D(d3_71__N_561[63]), .CK(osc_clk), .Q(d3[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i63.GSR = "ENABLED";
    FD1S3AX d3_i64 (.D(d3_71__N_561[64]), .CK(osc_clk), .Q(d3[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i64.GSR = "ENABLED";
    FD1S3AX d3_i65 (.D(d3_71__N_561[65]), .CK(osc_clk), .Q(d3[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i65.GSR = "ENABLED";
    FD1S3AX d3_i66 (.D(d3_71__N_561[66]), .CK(osc_clk), .Q(d3[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i66.GSR = "ENABLED";
    FD1S3AX d3_i67 (.D(d3_71__N_561[67]), .CK(osc_clk), .Q(d3[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i67.GSR = "ENABLED";
    FD1S3AX d3_i68 (.D(d3_71__N_561[68]), .CK(osc_clk), .Q(d3[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i68.GSR = "ENABLED";
    FD1S3AX d3_i69 (.D(d3_71__N_561[69]), .CK(osc_clk), .Q(d3[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i69.GSR = "ENABLED";
    FD1S3AX d3_i70 (.D(d3_71__N_561[70]), .CK(osc_clk), .Q(d3[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i70.GSR = "ENABLED";
    FD1S3AX d3_i71 (.D(d3_71__N_561[71]), .CK(osc_clk), .Q(d3[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i71.GSR = "ENABLED";
    FD1S3AX d4_i1 (.D(d4_71__N_633[1]), .CK(osc_clk), .Q(d4[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i1.GSR = "ENABLED";
    FD1S3AX d4_i2 (.D(d4_71__N_633[2]), .CK(osc_clk), .Q(d4[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i2.GSR = "ENABLED";
    FD1S3AX d4_i3 (.D(d4_71__N_633[3]), .CK(osc_clk), .Q(d4[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i3.GSR = "ENABLED";
    FD1S3AX d4_i4 (.D(d4_71__N_633[4]), .CK(osc_clk), .Q(d4[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i4.GSR = "ENABLED";
    FD1S3AX d4_i5 (.D(d4_71__N_633[5]), .CK(osc_clk), .Q(d4[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i5.GSR = "ENABLED";
    FD1S3AX d4_i6 (.D(d4_71__N_633[6]), .CK(osc_clk), .Q(d4[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i6.GSR = "ENABLED";
    FD1S3AX d4_i7 (.D(d4_71__N_633[7]), .CK(osc_clk), .Q(d4[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i7.GSR = "ENABLED";
    FD1S3AX d4_i8 (.D(d4_71__N_633[8]), .CK(osc_clk), .Q(d4[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i8.GSR = "ENABLED";
    FD1S3AX d4_i9 (.D(d4_71__N_633[9]), .CK(osc_clk), .Q(d4[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i9.GSR = "ENABLED";
    FD1S3AX d4_i10 (.D(d4_71__N_633[10]), .CK(osc_clk), .Q(d4[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i10.GSR = "ENABLED";
    FD1S3AX d4_i11 (.D(d4_71__N_633[11]), .CK(osc_clk), .Q(d4[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i11.GSR = "ENABLED";
    FD1S3AX d4_i12 (.D(d4_71__N_633[12]), .CK(osc_clk), .Q(d4[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i12.GSR = "ENABLED";
    FD1S3AX d4_i13 (.D(d4_71__N_633[13]), .CK(osc_clk), .Q(d4[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i13.GSR = "ENABLED";
    FD1S3AX d4_i14 (.D(d4_71__N_633[14]), .CK(osc_clk), .Q(d4[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i14.GSR = "ENABLED";
    FD1S3AX d4_i15 (.D(d4_71__N_633[15]), .CK(osc_clk), .Q(d4[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i15.GSR = "ENABLED";
    FD1S3AX d4_i16 (.D(d4_71__N_633[16]), .CK(osc_clk), .Q(d4[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i16.GSR = "ENABLED";
    FD1S3AX d4_i17 (.D(d4_71__N_633[17]), .CK(osc_clk), .Q(d4[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i17.GSR = "ENABLED";
    FD1S3AX d4_i18 (.D(d4_71__N_633[18]), .CK(osc_clk), .Q(d4[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i18.GSR = "ENABLED";
    FD1S3AX d4_i19 (.D(d4_71__N_633[19]), .CK(osc_clk), .Q(d4[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i19.GSR = "ENABLED";
    FD1S3AX d4_i20 (.D(d4_71__N_633[20]), .CK(osc_clk), .Q(d4[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i20.GSR = "ENABLED";
    FD1S3AX d4_i21 (.D(d4_71__N_633[21]), .CK(osc_clk), .Q(d4[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i21.GSR = "ENABLED";
    FD1S3AX d4_i22 (.D(d4_71__N_633[22]), .CK(osc_clk), .Q(d4[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i22.GSR = "ENABLED";
    FD1S3AX d4_i23 (.D(d4_71__N_633[23]), .CK(osc_clk), .Q(d4[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i23.GSR = "ENABLED";
    FD1S3AX d4_i24 (.D(d4_71__N_633[24]), .CK(osc_clk), .Q(d4[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i24.GSR = "ENABLED";
    FD1S3AX d4_i25 (.D(d4_71__N_633[25]), .CK(osc_clk), .Q(d4[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i25.GSR = "ENABLED";
    FD1S3AX d4_i26 (.D(d4_71__N_633[26]), .CK(osc_clk), .Q(d4[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i26.GSR = "ENABLED";
    FD1S3AX d4_i27 (.D(d4_71__N_633[27]), .CK(osc_clk), .Q(d4[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i27.GSR = "ENABLED";
    FD1S3AX d4_i28 (.D(d4_71__N_633[28]), .CK(osc_clk), .Q(d4[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i28.GSR = "ENABLED";
    FD1S3AX d4_i29 (.D(d4_71__N_633[29]), .CK(osc_clk), .Q(d4[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i29.GSR = "ENABLED";
    FD1S3AX d4_i30 (.D(d4_71__N_633[30]), .CK(osc_clk), .Q(d4[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i30.GSR = "ENABLED";
    FD1S3AX d4_i31 (.D(d4_71__N_633[31]), .CK(osc_clk), .Q(d4[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i31.GSR = "ENABLED";
    FD1S3AX d4_i32 (.D(d4_71__N_633[32]), .CK(osc_clk), .Q(d4[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i32.GSR = "ENABLED";
    FD1S3AX d4_i33 (.D(d4_71__N_633[33]), .CK(osc_clk), .Q(d4[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i33.GSR = "ENABLED";
    FD1S3AX d4_i34 (.D(d4_71__N_633[34]), .CK(osc_clk), .Q(d4[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i34.GSR = "ENABLED";
    FD1S3AX d4_i35 (.D(d4_71__N_633[35]), .CK(osc_clk), .Q(d4[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i35.GSR = "ENABLED";
    FD1S3AX d4_i36 (.D(d4_71__N_633[36]), .CK(osc_clk), .Q(d4[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i36.GSR = "ENABLED";
    FD1S3AX d4_i37 (.D(d4_71__N_633[37]), .CK(osc_clk), .Q(d4[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i37.GSR = "ENABLED";
    FD1S3AX d4_i38 (.D(d4_71__N_633[38]), .CK(osc_clk), .Q(d4[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i38.GSR = "ENABLED";
    FD1S3AX d4_i39 (.D(d4_71__N_633[39]), .CK(osc_clk), .Q(d4[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i39.GSR = "ENABLED";
    FD1S3AX d4_i40 (.D(d4_71__N_633[40]), .CK(osc_clk), .Q(d4[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i40.GSR = "ENABLED";
    FD1S3AX d4_i41 (.D(d4_71__N_633[41]), .CK(osc_clk), .Q(d4[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i41.GSR = "ENABLED";
    FD1S3AX d4_i42 (.D(d4_71__N_633[42]), .CK(osc_clk), .Q(d4[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i42.GSR = "ENABLED";
    FD1S3AX d4_i43 (.D(d4_71__N_633[43]), .CK(osc_clk), .Q(d4[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i43.GSR = "ENABLED";
    FD1S3AX d4_i44 (.D(d4_71__N_633[44]), .CK(osc_clk), .Q(d4[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i44.GSR = "ENABLED";
    FD1S3AX d4_i45 (.D(d4_71__N_633[45]), .CK(osc_clk), .Q(d4[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i45.GSR = "ENABLED";
    FD1S3AX d4_i46 (.D(d4_71__N_633[46]), .CK(osc_clk), .Q(d4[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i46.GSR = "ENABLED";
    FD1S3AX d4_i47 (.D(d4_71__N_633[47]), .CK(osc_clk), .Q(d4[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i47.GSR = "ENABLED";
    FD1S3AX d4_i48 (.D(d4_71__N_633[48]), .CK(osc_clk), .Q(d4[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i48.GSR = "ENABLED";
    FD1S3AX d4_i49 (.D(d4_71__N_633[49]), .CK(osc_clk), .Q(d4[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i49.GSR = "ENABLED";
    FD1S3AX d4_i50 (.D(d4_71__N_633[50]), .CK(osc_clk), .Q(d4[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i50.GSR = "ENABLED";
    FD1S3AX d4_i51 (.D(d4_71__N_633[51]), .CK(osc_clk), .Q(d4[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i51.GSR = "ENABLED";
    FD1S3AX d4_i52 (.D(d4_71__N_633[52]), .CK(osc_clk), .Q(d4[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i52.GSR = "ENABLED";
    FD1S3AX d4_i53 (.D(d4_71__N_633[53]), .CK(osc_clk), .Q(d4[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i53.GSR = "ENABLED";
    FD1S3AX d4_i54 (.D(d4_71__N_633[54]), .CK(osc_clk), .Q(d4[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i54.GSR = "ENABLED";
    FD1S3AX d4_i55 (.D(d4_71__N_633[55]), .CK(osc_clk), .Q(d4[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i55.GSR = "ENABLED";
    FD1S3AX d4_i56 (.D(d4_71__N_633[56]), .CK(osc_clk), .Q(d4[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i56.GSR = "ENABLED";
    FD1S3AX d4_i57 (.D(d4_71__N_633[57]), .CK(osc_clk), .Q(d4[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i57.GSR = "ENABLED";
    FD1S3AX d4_i58 (.D(d4_71__N_633[58]), .CK(osc_clk), .Q(d4[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i58.GSR = "ENABLED";
    FD1S3AX d4_i59 (.D(d4_71__N_633[59]), .CK(osc_clk), .Q(d4[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i59.GSR = "ENABLED";
    FD1S3AX d4_i60 (.D(d4_71__N_633[60]), .CK(osc_clk), .Q(d4[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i60.GSR = "ENABLED";
    FD1S3AX d4_i61 (.D(d4_71__N_633[61]), .CK(osc_clk), .Q(d4[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i61.GSR = "ENABLED";
    FD1S3AX d4_i62 (.D(d4_71__N_633[62]), .CK(osc_clk), .Q(d4[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i62.GSR = "ENABLED";
    FD1S3AX d4_i63 (.D(d4_71__N_633[63]), .CK(osc_clk), .Q(d4[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i63.GSR = "ENABLED";
    FD1S3AX d4_i64 (.D(d4_71__N_633[64]), .CK(osc_clk), .Q(d4[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i64.GSR = "ENABLED";
    FD1S3AX d4_i65 (.D(d4_71__N_633[65]), .CK(osc_clk), .Q(d4[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i65.GSR = "ENABLED";
    FD1S3AX d4_i66 (.D(d4_71__N_633[66]), .CK(osc_clk), .Q(d4[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i66.GSR = "ENABLED";
    FD1S3AX d4_i67 (.D(d4_71__N_633[67]), .CK(osc_clk), .Q(d4[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i67.GSR = "ENABLED";
    FD1S3AX d4_i68 (.D(d4_71__N_633[68]), .CK(osc_clk), .Q(d4[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i68.GSR = "ENABLED";
    FD1S3AX d4_i69 (.D(d4_71__N_633[69]), .CK(osc_clk), .Q(d4[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i69.GSR = "ENABLED";
    FD1S3AX d4_i70 (.D(d4_71__N_633[70]), .CK(osc_clk), .Q(d4[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i70.GSR = "ENABLED";
    FD1S3AX d4_i71 (.D(d4_71__N_633[71]), .CK(osc_clk), .Q(d4[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i71.GSR = "ENABLED";
    FD1S3AX d5_i1 (.D(d5_71__N_705[1]), .CK(osc_clk), .Q(d5[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i1.GSR = "ENABLED";
    FD1S3AX d5_i2 (.D(d5_71__N_705[2]), .CK(osc_clk), .Q(d5[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i2.GSR = "ENABLED";
    FD1S3AX d5_i3 (.D(d5_71__N_705[3]), .CK(osc_clk), .Q(d5[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i3.GSR = "ENABLED";
    FD1S3AX d5_i4 (.D(d5_71__N_705[4]), .CK(osc_clk), .Q(d5[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i4.GSR = "ENABLED";
    FD1S3AX d5_i5 (.D(d5_71__N_705[5]), .CK(osc_clk), .Q(d5[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i5.GSR = "ENABLED";
    FD1S3AX d5_i6 (.D(d5_71__N_705[6]), .CK(osc_clk), .Q(d5[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i6.GSR = "ENABLED";
    FD1S3AX d5_i7 (.D(d5_71__N_705[7]), .CK(osc_clk), .Q(d5[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i7.GSR = "ENABLED";
    FD1S3AX d5_i8 (.D(d5_71__N_705[8]), .CK(osc_clk), .Q(d5[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i8.GSR = "ENABLED";
    FD1S3AX d5_i9 (.D(d5_71__N_705[9]), .CK(osc_clk), .Q(d5[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i9.GSR = "ENABLED";
    FD1S3AX d5_i10 (.D(d5_71__N_705[10]), .CK(osc_clk), .Q(d5[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i10.GSR = "ENABLED";
    FD1S3AX d5_i11 (.D(d5_71__N_705[11]), .CK(osc_clk), .Q(d5[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i11.GSR = "ENABLED";
    FD1S3AX d5_i12 (.D(d5_71__N_705[12]), .CK(osc_clk), .Q(d5[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i12.GSR = "ENABLED";
    FD1S3AX d5_i13 (.D(d5_71__N_705[13]), .CK(osc_clk), .Q(d5[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i13.GSR = "ENABLED";
    FD1S3AX d5_i14 (.D(d5_71__N_705[14]), .CK(osc_clk), .Q(d5[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i14.GSR = "ENABLED";
    FD1S3AX d5_i15 (.D(d5_71__N_705[15]), .CK(osc_clk), .Q(d5[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i15.GSR = "ENABLED";
    FD1S3AX d5_i16 (.D(d5_71__N_705[16]), .CK(osc_clk), .Q(d5[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i16.GSR = "ENABLED";
    FD1S3AX d5_i17 (.D(d5_71__N_705[17]), .CK(osc_clk), .Q(d5[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i17.GSR = "ENABLED";
    FD1S3AX d5_i18 (.D(d5_71__N_705[18]), .CK(osc_clk), .Q(d5[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i18.GSR = "ENABLED";
    FD1S3AX d5_i19 (.D(d5_71__N_705[19]), .CK(osc_clk), .Q(d5[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i19.GSR = "ENABLED";
    FD1S3AX d5_i20 (.D(d5_71__N_705[20]), .CK(osc_clk), .Q(d5[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i20.GSR = "ENABLED";
    FD1S3AX d5_i21 (.D(d5_71__N_705[21]), .CK(osc_clk), .Q(d5[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i21.GSR = "ENABLED";
    FD1S3AX d5_i22 (.D(d5_71__N_705[22]), .CK(osc_clk), .Q(d5[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i22.GSR = "ENABLED";
    FD1S3AX d5_i23 (.D(d5_71__N_705[23]), .CK(osc_clk), .Q(d5[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i23.GSR = "ENABLED";
    FD1S3AX d5_i24 (.D(d5_71__N_705[24]), .CK(osc_clk), .Q(d5[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i24.GSR = "ENABLED";
    FD1S3AX d5_i25 (.D(d5_71__N_705[25]), .CK(osc_clk), .Q(d5[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i25.GSR = "ENABLED";
    FD1S3AX d5_i26 (.D(d5_71__N_705[26]), .CK(osc_clk), .Q(d5[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i26.GSR = "ENABLED";
    FD1S3AX d5_i27 (.D(d5_71__N_705[27]), .CK(osc_clk), .Q(d5[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i27.GSR = "ENABLED";
    FD1S3AX d5_i28 (.D(d5_71__N_705[28]), .CK(osc_clk), .Q(d5[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i28.GSR = "ENABLED";
    FD1S3AX d5_i29 (.D(d5_71__N_705[29]), .CK(osc_clk), .Q(d5[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i29.GSR = "ENABLED";
    FD1S3AX d5_i30 (.D(d5_71__N_705[30]), .CK(osc_clk), .Q(d5[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i30.GSR = "ENABLED";
    FD1S3AX d5_i31 (.D(d5_71__N_705[31]), .CK(osc_clk), .Q(d5[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i31.GSR = "ENABLED";
    FD1S3AX d5_i32 (.D(d5_71__N_705[32]), .CK(osc_clk), .Q(d5[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i32.GSR = "ENABLED";
    FD1S3AX d5_i33 (.D(d5_71__N_705[33]), .CK(osc_clk), .Q(d5[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i33.GSR = "ENABLED";
    FD1S3AX d5_i34 (.D(d5_71__N_705[34]), .CK(osc_clk), .Q(d5[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i34.GSR = "ENABLED";
    FD1S3AX d5_i35 (.D(d5_71__N_705[35]), .CK(osc_clk), .Q(d5[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i35.GSR = "ENABLED";
    FD1S3AX d5_i36 (.D(d5_71__N_705[36]), .CK(osc_clk), .Q(d5[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i36.GSR = "ENABLED";
    FD1S3AX d5_i37 (.D(d5_71__N_705[37]), .CK(osc_clk), .Q(d5[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i37.GSR = "ENABLED";
    FD1S3AX d5_i38 (.D(d5_71__N_705[38]), .CK(osc_clk), .Q(d5[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i38.GSR = "ENABLED";
    FD1S3AX d5_i39 (.D(d5_71__N_705[39]), .CK(osc_clk), .Q(d5[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i39.GSR = "ENABLED";
    FD1S3AX d5_i40 (.D(d5_71__N_705[40]), .CK(osc_clk), .Q(d5[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i40.GSR = "ENABLED";
    FD1S3AX d5_i41 (.D(d5_71__N_705[41]), .CK(osc_clk), .Q(d5[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i41.GSR = "ENABLED";
    FD1S3AX d5_i42 (.D(d5_71__N_705[42]), .CK(osc_clk), .Q(d5[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i42.GSR = "ENABLED";
    FD1S3AX d5_i43 (.D(d5_71__N_705[43]), .CK(osc_clk), .Q(d5[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i43.GSR = "ENABLED";
    FD1S3AX d5_i44 (.D(d5_71__N_705[44]), .CK(osc_clk), .Q(d5[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i44.GSR = "ENABLED";
    FD1S3AX d5_i45 (.D(d5_71__N_705[45]), .CK(osc_clk), .Q(d5[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i45.GSR = "ENABLED";
    FD1S3AX d5_i46 (.D(d5_71__N_705[46]), .CK(osc_clk), .Q(d5[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i46.GSR = "ENABLED";
    FD1S3AX d5_i47 (.D(d5_71__N_705[47]), .CK(osc_clk), .Q(d5[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i47.GSR = "ENABLED";
    FD1S3AX d5_i48 (.D(d5_71__N_705[48]), .CK(osc_clk), .Q(d5[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i48.GSR = "ENABLED";
    FD1S3AX d5_i49 (.D(d5_71__N_705[49]), .CK(osc_clk), .Q(d5[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i49.GSR = "ENABLED";
    FD1S3AX d5_i50 (.D(d5_71__N_705[50]), .CK(osc_clk), .Q(d5[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i50.GSR = "ENABLED";
    FD1S3AX d5_i51 (.D(d5_71__N_705[51]), .CK(osc_clk), .Q(d5[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i51.GSR = "ENABLED";
    FD1S3AX d5_i52 (.D(d5_71__N_705[52]), .CK(osc_clk), .Q(d5[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i52.GSR = "ENABLED";
    FD1S3AX d5_i53 (.D(d5_71__N_705[53]), .CK(osc_clk), .Q(d5[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i53.GSR = "ENABLED";
    FD1S3AX d5_i54 (.D(d5_71__N_705[54]), .CK(osc_clk), .Q(d5[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i54.GSR = "ENABLED";
    FD1S3AX d5_i55 (.D(d5_71__N_705[55]), .CK(osc_clk), .Q(d5[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i55.GSR = "ENABLED";
    FD1S3AX d5_i56 (.D(d5_71__N_705[56]), .CK(osc_clk), .Q(d5[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i56.GSR = "ENABLED";
    FD1S3AX d5_i57 (.D(d5_71__N_705[57]), .CK(osc_clk), .Q(d5[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i57.GSR = "ENABLED";
    FD1S3AX d5_i58 (.D(d5_71__N_705[58]), .CK(osc_clk), .Q(d5[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i58.GSR = "ENABLED";
    FD1S3AX d5_i59 (.D(d5_71__N_705[59]), .CK(osc_clk), .Q(d5[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i59.GSR = "ENABLED";
    FD1S3AX d5_i60 (.D(d5_71__N_705[60]), .CK(osc_clk), .Q(d5[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i60.GSR = "ENABLED";
    FD1S3AX d5_i61 (.D(d5_71__N_705[61]), .CK(osc_clk), .Q(d5[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i61.GSR = "ENABLED";
    FD1S3AX d5_i62 (.D(d5_71__N_705[62]), .CK(osc_clk), .Q(d5[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i62.GSR = "ENABLED";
    FD1S3AX d5_i63 (.D(d5_71__N_705[63]), .CK(osc_clk), .Q(d5[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i63.GSR = "ENABLED";
    FD1S3AX d5_i64 (.D(d5_71__N_705[64]), .CK(osc_clk), .Q(d5[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i64.GSR = "ENABLED";
    FD1S3AX d5_i65 (.D(d5_71__N_705[65]), .CK(osc_clk), .Q(d5[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i65.GSR = "ENABLED";
    FD1S3AX d5_i66 (.D(d5_71__N_705[66]), .CK(osc_clk), .Q(d5[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i66.GSR = "ENABLED";
    FD1S3AX d5_i67 (.D(d5_71__N_705[67]), .CK(osc_clk), .Q(d5[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i67.GSR = "ENABLED";
    FD1S3AX d5_i68 (.D(d5_71__N_705[68]), .CK(osc_clk), .Q(d5[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i68.GSR = "ENABLED";
    FD1S3AX d5_i69 (.D(d5_71__N_705[69]), .CK(osc_clk), .Q(d5[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i69.GSR = "ENABLED";
    FD1S3AX d5_i70 (.D(d5_71__N_705[70]), .CK(osc_clk), .Q(d5[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i70.GSR = "ENABLED";
    FD1S3AX d5_i71 (.D(d5_71__N_705[71]), .CK(osc_clk), .Q(d5[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i71.GSR = "ENABLED";
    FD1P3AX d6_i0_i1 (.D(d6_71__N_1458[1]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d6_i0_i2 (.D(d6_71__N_1458[2]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d6_i0_i3 (.D(d6_71__N_1458[3]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d6_i0_i4 (.D(d6_71__N_1458[4]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d6_i0_i5 (.D(d6_71__N_1458[5]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d6_i0_i6 (.D(d6_71__N_1458[6]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d6_i0_i7 (.D(d6_71__N_1458[7]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d6_i0_i8 (.D(d6_71__N_1458[8]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d6_i0_i9 (.D(d6_71__N_1458[9]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d6_i0_i10 (.D(d6_71__N_1458[10]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d6_i0_i11 (.D(d6_71__N_1458[11]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d6_i0_i12 (.D(d6_71__N_1458[12]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d6_i0_i13 (.D(d6_71__N_1458[13]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d6_i0_i14 (.D(d6_71__N_1458[14]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d6_i0_i15 (.D(d6_71__N_1458[15]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d6_i0_i16 (.D(d6_71__N_1458[16]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d6_i0_i17 (.D(d6_71__N_1458[17]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d6_i0_i18 (.D(d6_71__N_1458[18]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d6_i0_i19 (.D(d6_71__N_1458[19]), .SP(osc_clk_enable_146), .CK(osc_clk), 
            .Q(d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d6_i0_i20 (.D(d6_71__N_1458[20]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d6_i0_i21 (.D(d6_71__N_1458[21]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d6_i0_i22 (.D(d6_71__N_1458[22]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d6_i0_i23 (.D(d6_71__N_1458[23]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d6_i0_i24 (.D(d6_71__N_1458[24]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d6_i0_i25 (.D(d6_71__N_1458[25]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d6_i0_i26 (.D(d6_71__N_1458[26]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d6_i0_i27 (.D(d6_71__N_1458[27]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d6_i0_i28 (.D(d6_71__N_1458[28]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d6_i0_i29 (.D(d6_71__N_1458[29]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d6_i0_i30 (.D(d6_71__N_1458[30]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d6_i0_i31 (.D(d6_71__N_1458[31]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d6_i0_i32 (.D(d6_71__N_1458[32]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d6_i0_i33 (.D(d6_71__N_1458[33]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d6_i0_i34 (.D(d6_71__N_1458[34]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d6_i0_i35 (.D(d6_71__N_1458[35]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d6_i0_i36 (.D(d6_71__N_1458[36]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d6_i0_i37 (.D(d6_71__N_1458[37]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d6_i0_i38 (.D(d6_71__N_1458[38]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d6_i0_i39 (.D(d6_71__N_1458[39]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d6_i0_i40 (.D(d6_71__N_1458[40]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d6_i0_i41 (.D(d6_71__N_1458[41]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d6_i0_i42 (.D(d6_71__N_1458[42]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d6_i0_i43 (.D(d6_71__N_1458[43]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d6_i0_i44 (.D(d6_71__N_1458[44]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d6_i0_i45 (.D(d6_71__N_1458[45]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d6_i0_i46 (.D(d6_71__N_1458[46]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d6_i0_i47 (.D(d6_71__N_1458[47]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d6_i0_i48 (.D(d6_71__N_1458[48]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d6_i0_i49 (.D(d6_71__N_1458[49]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d6_i0_i50 (.D(d6_71__N_1458[50]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d6_i0_i51 (.D(d6_71__N_1458[51]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d6_i0_i52 (.D(d6_71__N_1458[52]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d6_i0_i53 (.D(d6_71__N_1458[53]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d6_i0_i54 (.D(d6_71__N_1458[54]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d6_i0_i55 (.D(d6_71__N_1458[55]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d6_i0_i56 (.D(d6_71__N_1458[56]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d6_i0_i57 (.D(d6_71__N_1458[57]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d6_i0_i58 (.D(d6_71__N_1458[58]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d6_i0_i59 (.D(d6_71__N_1458[59]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d6_i0_i60 (.D(d6_71__N_1458[60]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d6_i0_i61 (.D(d6_71__N_1458[61]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d6_i0_i62 (.D(d6_71__N_1458[62]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d6_i0_i63 (.D(d6_71__N_1458[63]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d6_i0_i64 (.D(d6_71__N_1458[64]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d6_i0_i65 (.D(d6_71__N_1458[65]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d6_i0_i66 (.D(d6_71__N_1458[66]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d6_i0_i67 (.D(d6_71__N_1458[67]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d6_i0_i68 (.D(d6_71__N_1458[68]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d6_i0_i69 (.D(d6_71__N_1458[69]), .SP(osc_clk_enable_196), .CK(osc_clk), 
            .Q(d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d6_i0_i70 (.D(d6_71__N_1458[70]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d6_i0_i71 (.D(d6_71__N_1458[71]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i1 (.D(d6[1]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i2 (.D(d6[2]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i3 (.D(d6[3]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i4 (.D(d6[4]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i5 (.D(d6[5]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i6 (.D(d6[6]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i7 (.D(d6[7]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i8 (.D(d6[8]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i9 (.D(d6[9]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i10 (.D(d6[10]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i11 (.D(d6[11]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i12 (.D(d6[12]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i13 (.D(d6[13]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i14 (.D(d6[14]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i15 (.D(d6[15]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i16 (.D(d6[16]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i17 (.D(d6[17]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i18 (.D(d6[18]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i19 (.D(d6[19]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i20 (.D(d6[20]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i21 (.D(d6[21]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i22 (.D(d6[22]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i23 (.D(d6[23]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i24 (.D(d6[24]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i25 (.D(d6[25]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i26 (.D(d6[26]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i27 (.D(d6[27]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i28 (.D(d6[28]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i29 (.D(d6[29]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i30 (.D(d6[30]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i31 (.D(d6[31]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i32 (.D(d6[32]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i33 (.D(d6[33]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i34 (.D(d6[34]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i35 (.D(d6[35]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i36 (.D(d6[36]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i37 (.D(d6[37]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i38 (.D(d6[38]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i39 (.D(d6[39]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i40 (.D(d6[40]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i41 (.D(d6[41]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i42 (.D(d6[42]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i43 (.D(d6[43]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i44 (.D(d6[44]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i45 (.D(d6[45]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i46 (.D(d6[46]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i47 (.D(d6[47]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i48 (.D(d6[48]), .SP(osc_clk_enable_246), .CK(osc_clk), 
            .Q(d_d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i49 (.D(d6[49]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d_d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i50 (.D(d6[50]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d_d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i51 (.D(d6[51]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d_d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i52 (.D(d6[52]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d_d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i53 (.D(d6[53]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d_d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i54 (.D(d6[54]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d_d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i55 (.D(d6[55]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d_d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i56 (.D(d6[56]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d_d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i57 (.D(d6[57]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d_d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i58 (.D(d6[58]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d_d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i59 (.D(d6[59]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d_d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i60 (.D(d6[60]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d_d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i61 (.D(d6[61]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d_d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i62 (.D(d6[62]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d_d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i63 (.D(d6[63]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d_d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i64 (.D(d6[64]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d_d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i65 (.D(d6[65]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d_d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i66 (.D(d6[66]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d_d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i67 (.D(d6[67]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d_d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i68 (.D(d6[68]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d_d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i69 (.D(d6[69]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d_d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i70 (.D(d6[70]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d_d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i71 (.D(d6[71]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d_d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d7_i0_i1 (.D(d7_71__N_1530[1]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d7_i0_i2 (.D(d7_71__N_1530[2]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d7_i0_i3 (.D(d7_71__N_1530[3]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d7_i0_i4 (.D(d7_71__N_1530[4]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d7_i0_i5 (.D(d7_71__N_1530[5]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d7_i0_i6 (.D(d7_71__N_1530[6]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d7_i0_i7 (.D(d7_71__N_1530[7]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d7_i0_i8 (.D(d7_71__N_1530[8]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d7_i0_i9 (.D(d7_71__N_1530[9]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d7_i0_i10 (.D(d7_71__N_1530[10]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d7_i0_i11 (.D(d7_71__N_1530[11]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d7_i0_i12 (.D(d7_71__N_1530[12]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d7_i0_i13 (.D(d7_71__N_1530[13]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d7_i0_i14 (.D(d7_71__N_1530[14]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d7_i0_i15 (.D(d7_71__N_1530[15]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d7_i0_i16 (.D(d7_71__N_1530[16]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d7_i0_i17 (.D(d7_71__N_1530[17]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d7_i0_i18 (.D(d7_71__N_1530[18]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d7_i0_i19 (.D(d7_71__N_1530[19]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d7_i0_i20 (.D(d7_71__N_1530[20]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d7_i0_i21 (.D(d7_71__N_1530[21]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d7_i0_i22 (.D(d7_71__N_1530[22]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d7_i0_i23 (.D(d7_71__N_1530[23]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d7_i0_i24 (.D(d7_71__N_1530[24]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d7_i0_i25 (.D(d7_71__N_1530[25]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d7_i0_i26 (.D(d7_71__N_1530[26]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d7_i0_i27 (.D(d7_71__N_1530[27]), .SP(osc_clk_enable_296), .CK(osc_clk), 
            .Q(d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d7_i0_i28 (.D(d7_71__N_1530[28]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d7_i0_i29 (.D(d7_71__N_1530[29]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d7_i0_i30 (.D(d7_71__N_1530[30]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d7_i0_i31 (.D(d7_71__N_1530[31]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d7_i0_i32 (.D(d7_71__N_1530[32]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d7_i0_i33 (.D(d7_71__N_1530[33]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d7_i0_i34 (.D(d7_71__N_1530[34]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d7_i0_i35 (.D(d7_71__N_1530[35]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d7_i0_i36 (.D(d7_71__N_1530[36]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d7_i0_i37 (.D(d7_71__N_1530[37]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d7_i0_i38 (.D(d7_71__N_1530[38]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d7_i0_i39 (.D(d7_71__N_1530[39]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d7_i0_i40 (.D(d7_71__N_1530[40]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d7_i0_i41 (.D(d7_71__N_1530[41]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d7_i0_i42 (.D(d7_71__N_1530[42]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d7_i0_i43 (.D(d7_71__N_1530[43]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d7_i0_i44 (.D(d7_71__N_1530[44]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d7_i0_i45 (.D(d7_71__N_1530[45]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d7_i0_i46 (.D(d7_71__N_1530[46]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d7_i0_i47 (.D(d7_71__N_1530[47]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d7_i0_i48 (.D(d7_71__N_1530[48]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d7_i0_i49 (.D(d7_71__N_1530[49]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d7_i0_i50 (.D(d7_71__N_1530[50]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d7_i0_i51 (.D(d7_71__N_1530[51]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d7_i0_i52 (.D(d7_71__N_1530[52]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d7_i0_i53 (.D(d7_71__N_1530[53]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d7_i0_i54 (.D(d7_71__N_1530[54]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d7_i0_i55 (.D(d7_71__N_1530[55]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d7_i0_i56 (.D(d7_71__N_1530[56]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d7_i0_i57 (.D(d7_71__N_1530[57]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d7_i0_i58 (.D(d7_71__N_1530[58]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d7_i0_i59 (.D(d7_71__N_1530[59]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d7_i0_i60 (.D(d7_71__N_1530[60]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d7_i0_i61 (.D(d7_71__N_1530[61]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d7_i0_i62 (.D(d7_71__N_1530[62]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d7_i0_i63 (.D(d7_71__N_1530[63]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d7_i0_i64 (.D(d7_71__N_1530[64]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d7_i0_i65 (.D(d7_71__N_1530[65]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d7_i0_i66 (.D(d7_71__N_1530[66]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d7_i0_i67 (.D(d7_71__N_1530[67]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d7_i0_i68 (.D(d7_71__N_1530[68]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d7_i0_i69 (.D(d7_71__N_1530[69]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d7_i0_i70 (.D(d7_71__N_1530[70]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d7_i0_i71 (.D(d7_71__N_1530[71]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i1 (.D(d7[1]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d_d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i2 (.D(d7[2]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d_d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i3 (.D(d7[3]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d_d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i4 (.D(d7[4]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d_d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i5 (.D(d7[5]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d_d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i6 (.D(d7[6]), .SP(osc_clk_enable_346), .CK(osc_clk), 
            .Q(d_d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i7 (.D(d7[7]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i8 (.D(d7[8]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i9 (.D(d7[9]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i10 (.D(d7[10]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i11 (.D(d7[11]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i12 (.D(d7[12]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i13 (.D(d7[13]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i14 (.D(d7[14]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i15 (.D(d7[15]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i16 (.D(d7[16]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i17 (.D(d7[17]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i18 (.D(d7[18]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i19 (.D(d7[19]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i20 (.D(d7[20]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i21 (.D(d7[21]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i22 (.D(d7[22]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i23 (.D(d7[23]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i24 (.D(d7[24]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i25 (.D(d7[25]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i26 (.D(d7[26]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i27 (.D(d7[27]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i28 (.D(d7[28]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i29 (.D(d7[29]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i30 (.D(d7[30]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i31 (.D(d7[31]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i32 (.D(d7[32]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i33 (.D(d7[33]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i34 (.D(d7[34]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i35 (.D(d7[35]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i36 (.D(d7[36]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i37 (.D(d7[37]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i38 (.D(d7[38]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i39 (.D(d7[39]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i40 (.D(d7[40]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i41 (.D(d7[41]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i42 (.D(d7[42]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i43 (.D(d7[43]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i44 (.D(d7[44]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i45 (.D(d7[45]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i46 (.D(d7[46]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i47 (.D(d7[47]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i48 (.D(d7[48]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i49 (.D(d7[49]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i50 (.D(d7[50]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i51 (.D(d7[51]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i52 (.D(d7[52]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i53 (.D(d7[53]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i54 (.D(d7[54]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i55 (.D(d7[55]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i56 (.D(d7[56]), .SP(osc_clk_enable_396), .CK(osc_clk), 
            .Q(d_d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i57 (.D(d7[57]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d_d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i58 (.D(d7[58]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d_d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i59 (.D(d7[59]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d_d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i60 (.D(d7[60]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d_d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i61 (.D(d7[61]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d_d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i62 (.D(d7[62]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d_d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i63 (.D(d7[63]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d_d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i64 (.D(d7[64]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d_d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i65 (.D(d7[65]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d_d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i66 (.D(d7[66]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d_d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i67 (.D(d7[67]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d_d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i68 (.D(d7[68]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d_d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i69 (.D(d7[69]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d_d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i70 (.D(d7[70]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d_d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i71 (.D(d7[71]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d_d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d8_i0_i1 (.D(d8_71__N_1602[1]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d8_i0_i2 (.D(d8_71__N_1602[2]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d8_i0_i3 (.D(d8_71__N_1602[3]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d8_i0_i4 (.D(d8_71__N_1602[4]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d8_i0_i5 (.D(d8_71__N_1602[5]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d8_i0_i6 (.D(d8_71__N_1602[6]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d8_i0_i7 (.D(d8_71__N_1602[7]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d8_i0_i8 (.D(d8_71__N_1602[8]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d8_i0_i9 (.D(d8_71__N_1602[9]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d8_i0_i10 (.D(d8_71__N_1602[10]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d8_i0_i11 (.D(d8_71__N_1602[11]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d8_i0_i12 (.D(d8_71__N_1602[12]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d8_i0_i13 (.D(d8_71__N_1602[13]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d8_i0_i14 (.D(d8_71__N_1602[14]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d8_i0_i15 (.D(d8_71__N_1602[15]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d8_i0_i16 (.D(d8_71__N_1602[16]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d8_i0_i17 (.D(d8_71__N_1602[17]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d8_i0_i18 (.D(d8_71__N_1602[18]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d8_i0_i19 (.D(d8_71__N_1602[19]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d8_i0_i20 (.D(d8_71__N_1602[20]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d8_i0_i21 (.D(d8_71__N_1602[21]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d8_i0_i22 (.D(d8_71__N_1602[22]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d8_i0_i23 (.D(d8_71__N_1602[23]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d8_i0_i24 (.D(d8_71__N_1602[24]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d8_i0_i25 (.D(d8_71__N_1602[25]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d8_i0_i26 (.D(d8_71__N_1602[26]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d8_i0_i27 (.D(d8_71__N_1602[27]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d8_i0_i28 (.D(d8_71__N_1602[28]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d8_i0_i29 (.D(d8_71__N_1602[29]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d8_i0_i30 (.D(d8_71__N_1602[30]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d8_i0_i31 (.D(d8_71__N_1602[31]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d8_i0_i32 (.D(d8_71__N_1602[32]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d8_i0_i33 (.D(d8_71__N_1602[33]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d8_i0_i34 (.D(d8_71__N_1602[34]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d8_i0_i35 (.D(d8_71__N_1602[35]), .SP(osc_clk_enable_446), .CK(osc_clk), 
            .Q(d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d8_i0_i36 (.D(d8_71__N_1602[36]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d8_i0_i37 (.D(d8_71__N_1602[37]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d8_i0_i38 (.D(d8_71__N_1602[38]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d8_i0_i39 (.D(d8_71__N_1602[39]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d8_i0_i40 (.D(d8_71__N_1602[40]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d8_i0_i41 (.D(d8_71__N_1602[41]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d8_i0_i42 (.D(d8_71__N_1602[42]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d8_i0_i43 (.D(d8_71__N_1602[43]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d8_i0_i44 (.D(d8_71__N_1602[44]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d8_i0_i45 (.D(d8_71__N_1602[45]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d8_i0_i46 (.D(d8_71__N_1602[46]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d8_i0_i47 (.D(d8_71__N_1602[47]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d8_i0_i48 (.D(d8_71__N_1602[48]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d8_i0_i49 (.D(d8_71__N_1602[49]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d8_i0_i50 (.D(d8_71__N_1602[50]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d8_i0_i51 (.D(d8_71__N_1602[51]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d8_i0_i52 (.D(d8_71__N_1602[52]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d8_i0_i53 (.D(d8_71__N_1602[53]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d8_i0_i54 (.D(d8_71__N_1602[54]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d8_i0_i55 (.D(d8_71__N_1602[55]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d8_i0_i56 (.D(d8_71__N_1602[56]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d8_i0_i57 (.D(d8_71__N_1602[57]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d8_i0_i58 (.D(d8_71__N_1602[58]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d8_i0_i59 (.D(d8_71__N_1602[59]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d8_i0_i60 (.D(d8_71__N_1602[60]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d8_i0_i61 (.D(d8_71__N_1602[61]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d8_i0_i62 (.D(d8_71__N_1602[62]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d8_i0_i63 (.D(d8_71__N_1602[63]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d8_i0_i64 (.D(d8_71__N_1602[64]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d8_i0_i65 (.D(d8_71__N_1602[65]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d8_i0_i66 (.D(d8_71__N_1602[66]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d8_i0_i67 (.D(d8_71__N_1602[67]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d8_i0_i68 (.D(d8_71__N_1602[68]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d8_i0_i69 (.D(d8_71__N_1602[69]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d8_i0_i70 (.D(d8_71__N_1602[70]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d8_i0_i71 (.D(d8_71__N_1602[71]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i1 (.D(d8[1]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d_d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i2 (.D(d8[2]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d_d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i3 (.D(d8[3]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d_d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i4 (.D(d8[4]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d_d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i5 (.D(d8[5]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d_d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i6 (.D(d8[6]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d_d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i7 (.D(d8[7]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d_d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i8 (.D(d8[8]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d_d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i9 (.D(d8[9]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d_d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i10 (.D(d8[10]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d_d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i11 (.D(d8[11]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d_d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i12 (.D(d8[12]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d_d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i13 (.D(d8[13]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d_d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i14 (.D(d8[14]), .SP(osc_clk_enable_496), .CK(osc_clk), 
            .Q(d_d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i15 (.D(d8[15]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i16 (.D(d8[16]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i17 (.D(d8[17]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i18 (.D(d8[18]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i19 (.D(d8[19]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i20 (.D(d8[20]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i21 (.D(d8[21]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i22 (.D(d8[22]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i23 (.D(d8[23]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i24 (.D(d8[24]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i25 (.D(d8[25]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i26 (.D(d8[26]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i27 (.D(d8[27]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i28 (.D(d8[28]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i29 (.D(d8[29]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i30 (.D(d8[30]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i31 (.D(d8[31]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i32 (.D(d8[32]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i33 (.D(d8[33]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i34 (.D(d8[34]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i35 (.D(d8[35]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i36 (.D(d8[36]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i37 (.D(d8[37]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i38 (.D(d8[38]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i39 (.D(d8[39]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i40 (.D(d8[40]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i41 (.D(d8[41]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i42 (.D(d8[42]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i43 (.D(d8[43]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i44 (.D(d8[44]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i45 (.D(d8[45]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i46 (.D(d8[46]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i47 (.D(d8[47]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i48 (.D(d8[48]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i49 (.D(d8[49]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i50 (.D(d8[50]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i51 (.D(d8[51]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i52 (.D(d8[52]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i53 (.D(d8[53]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i54 (.D(d8[54]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i55 (.D(d8[55]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i56 (.D(d8[56]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i57 (.D(d8[57]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i58 (.D(d8[58]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i59 (.D(d8[59]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i60 (.D(d8[60]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i61 (.D(d8[61]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i62 (.D(d8[62]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i63 (.D(d8[63]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i64 (.D(d8[64]), .SP(osc_clk_enable_546), .CK(osc_clk), 
            .Q(d_d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i65 (.D(d8[65]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d_d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i66 (.D(d8[66]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d_d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i67 (.D(d8[67]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d_d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i68 (.D(d8[68]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d_d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i69 (.D(d8[69]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d_d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i70 (.D(d8[70]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d_d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i71 (.D(d8[71]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d_d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d9_i0_i1 (.D(d9_71__N_1674[1]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d9_i0_i2 (.D(d9_71__N_1674[2]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d9_i0_i3 (.D(d9_71__N_1674[3]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d9_i0_i4 (.D(d9_71__N_1674[4]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d9_i0_i5 (.D(d9_71__N_1674[5]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d9_i0_i6 (.D(d9_71__N_1674[6]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d9_i0_i7 (.D(d9_71__N_1674[7]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d9_i0_i8 (.D(d9_71__N_1674[8]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d9_i0_i9 (.D(d9_71__N_1674[9]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d9_i0_i10 (.D(d9_71__N_1674[10]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d9_i0_i11 (.D(d9_71__N_1674[11]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d9_i0_i12 (.D(d9_71__N_1674[12]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d9_i0_i13 (.D(d9_71__N_1674[13]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d9_i0_i14 (.D(d9_71__N_1674[14]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d9_i0_i15 (.D(d9_71__N_1674[15]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d9_i0_i16 (.D(d9_71__N_1674[16]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d9_i0_i17 (.D(d9_71__N_1674[17]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d9_i0_i18 (.D(d9_71__N_1674[18]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d9_i0_i19 (.D(d9_71__N_1674[19]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d9_i0_i20 (.D(d9_71__N_1674[20]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d9_i0_i21 (.D(d9_71__N_1674[21]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d9_i0_i22 (.D(d9_71__N_1674[22]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d9_i0_i23 (.D(d9_71__N_1674[23]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d9_i0_i24 (.D(d9_71__N_1674[24]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d9_i0_i25 (.D(d9_71__N_1674[25]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d9_i0_i26 (.D(d9_71__N_1674[26]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d9_i0_i27 (.D(d9_71__N_1674[27]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d9_i0_i28 (.D(d9_71__N_1674[28]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d9_i0_i29 (.D(d9_71__N_1674[29]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d9_i0_i30 (.D(d9_71__N_1674[30]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d9_i0_i31 (.D(d9_71__N_1674[31]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d9_i0_i32 (.D(d9_71__N_1674[32]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d9_i0_i33 (.D(d9_71__N_1674[33]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d9_i0_i34 (.D(d9_71__N_1674[34]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d9_i0_i35 (.D(d9_71__N_1674[35]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d9_i0_i36 (.D(d9_71__N_1674[36]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d9_i0_i37 (.D(d9_71__N_1674[37]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d9_i0_i38 (.D(d9_71__N_1674[38]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d9_i0_i39 (.D(d9_71__N_1674[39]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d9_i0_i40 (.D(d9_71__N_1674[40]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d9_i0_i41 (.D(d9_71__N_1674[41]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d9_i0_i42 (.D(d9_71__N_1674[42]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d9_i0_i43 (.D(d9_71__N_1674[43]), .SP(osc_clk_enable_596), .CK(osc_clk), 
            .Q(d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d9_i0_i44 (.D(d9_71__N_1674[44]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d9_i0_i45 (.D(d9_71__N_1674[45]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d9_i0_i46 (.D(d9_71__N_1674[46]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d9_i0_i47 (.D(d9_71__N_1674[47]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d9_i0_i48 (.D(d9_71__N_1674[48]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d9_i0_i49 (.D(d9_71__N_1674[49]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d9_i0_i50 (.D(d9_71__N_1674[50]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d9_i0_i51 (.D(d9_71__N_1674[51]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d9_i0_i52 (.D(d9_71__N_1674[52]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d9_i0_i53 (.D(d9_71__N_1674[53]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d9_i0_i54 (.D(d9_71__N_1674[54]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d9_i0_i55 (.D(d9_71__N_1674[55]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d9_i0_i56 (.D(d9_71__N_1674[56]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d9_i0_i57 (.D(d9_71__N_1674[57]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d9_i0_i58 (.D(d9_71__N_1674[58]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d9_i0_i59 (.D(d9_71__N_1674[59]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d9_i0_i60 (.D(d9_71__N_1674[60]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d9_i0_i61 (.D(d9_71__N_1674[61]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d9_i0_i62 (.D(d9_71__N_1674[62]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d9_i0_i63 (.D(d9_71__N_1674[63]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d9_i0_i64 (.D(d9_71__N_1674[64]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d9_i0_i65 (.D(d9_71__N_1674[65]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d9_i0_i66 (.D(d9_71__N_1674[66]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d9_i0_i67 (.D(d9_71__N_1674[67]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d9_i0_i68 (.D(d9_71__N_1674[68]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d9_i0_i69 (.D(d9_71__N_1674[69]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d9_i0_i70 (.D(d9_71__N_1674[70]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d9_i0_i71 (.D(d9_71__N_1674[71]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i1 (.D(d9[1]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d_d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i2 (.D(d9[2]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d_d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i3 (.D(d9[3]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d_d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i4 (.D(d9[4]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d_d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i5 (.D(d9[5]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d_d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i6 (.D(d9[6]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d_d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i7 (.D(d9[7]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d_d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i8 (.D(d9[8]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d_d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i9 (.D(d9[9]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d_d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i10 (.D(d9[10]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d_d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i11 (.D(d9[11]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d_d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i12 (.D(d9[12]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d_d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i13 (.D(d9[13]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d_d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i14 (.D(d9[14]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d_d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i15 (.D(d9[15]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d_d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i16 (.D(d9[16]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d_d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i17 (.D(d9[17]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d_d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i18 (.D(d9[18]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d_d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i19 (.D(d9[19]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d_d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i20 (.D(d9[20]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d_d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i21 (.D(d9[21]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d_d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i22 (.D(d9[22]), .SP(osc_clk_enable_646), .CK(osc_clk), 
            .Q(d_d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i23 (.D(d9[23]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i24 (.D(d9[24]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i25 (.D(d9[25]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i26 (.D(d9[26]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i27 (.D(d9[27]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i28 (.D(d9[28]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i29 (.D(d9[29]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i30 (.D(d9[30]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i31 (.D(d9[31]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i32 (.D(d9[32]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i33 (.D(d9[33]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i34 (.D(d9[34]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i35 (.D(d9[35]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i36 (.D(d9[36]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i37 (.D(d9[37]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i38 (.D(d9[38]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i39 (.D(d9[39]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i40 (.D(d9[40]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i41 (.D(d9[41]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i42 (.D(d9[42]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i43 (.D(d9[43]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i44 (.D(d9[44]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i45 (.D(d9[45]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i46 (.D(d9[46]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i47 (.D(d9[47]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i48 (.D(d9[48]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i49 (.D(d9[49]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i50 (.D(d9[50]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i51 (.D(d9[51]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i52 (.D(d9[52]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i53 (.D(d9[53]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i54 (.D(d9[54]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i55 (.D(d9[55]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i56 (.D(d9[56]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i57 (.D(d9[57]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i58 (.D(d9[58]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i59 (.D(d9[59]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i60 (.D(d9[60]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i61 (.D(d9[61]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i62 (.D(d9[62]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i63 (.D(d9[63]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i64 (.D(d9[64]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i65 (.D(d9[65]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i66 (.D(d9[66]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i67 (.D(d9[67]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i68 (.D(d9[68]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i69 (.D(d9[69]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i70 (.D(d9[70]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i71 (.D(d9[71]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d_d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d10__i2 (.D(d10_71__N_1746[57]), .SP(osc_clk_enable_696), .CK(osc_clk), 
            .Q(d10[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i2.GSR = "ENABLED";
    FD1P3AX d10__i3 (.D(d10_71__N_1746[58]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i3.GSR = "ENABLED";
    FD1P3AX d10__i4 (.D(d10_71__N_1746[59]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i4.GSR = "ENABLED";
    FD1P3AX d10__i5 (.D(d10_71__N_1746[60]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i5.GSR = "ENABLED";
    FD1P3AX d10__i6 (.D(d10_71__N_1746[61]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i6.GSR = "ENABLED";
    FD1P3AX d10__i7 (.D(d10_71__N_1746[62]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i7.GSR = "ENABLED";
    FD1P3AX d10__i8 (.D(d10_71__N_1746[63]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i8.GSR = "ENABLED";
    FD1P3AX d10__i9 (.D(d10_71__N_1746[64]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i9.GSR = "ENABLED";
    FD1P3AX d10__i10 (.D(d10_71__N_1746[65]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i10.GSR = "ENABLED";
    FD1P3AX d10__i11 (.D(d10_71__N_1746[66]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i11.GSR = "ENABLED";
    FD1P3AX d10__i12 (.D(d10_71__N_1746[67]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i12.GSR = "ENABLED";
    FD1P3AX d10__i13 (.D(d10_71__N_1746[68]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i13.GSR = "ENABLED";
    FD1P3AX d10__i14 (.D(d10_71__N_1746[69]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i14.GSR = "ENABLED";
    FD1P3AX d10__i15 (.D(d10_71__N_1746[70]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i15.GSR = "ENABLED";
    FD1P3AX d10__i16 (.D(d10_71__N_1746[71]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i16.GSR = "ENABLED";
    FD1P3AX d_out_i0_i1 (.D(d_out_11__N_1818[1]), .SP(v_comb), .CK(osc_clk), 
            .Q(\CIC1_outSin[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i1.GSR = "ENABLED";
    FD1P3AX d_out_i0_i2 (.D(d_out_11__N_1818[2]), .SP(v_comb), .CK(osc_clk), 
            .Q(\CIC1_outSin[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i2.GSR = "ENABLED";
    FD1P3AX d_out_i0_i3 (.D(d_out_11__N_1818[3]), .SP(v_comb), .CK(osc_clk), 
            .Q(\CIC1_outSin[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i3.GSR = "ENABLED";
    FD1P3AX d_out_i0_i4 (.D(d_out_11__N_1818[4]), .SP(v_comb), .CK(osc_clk), 
            .Q(\CIC1_outSin[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i4.GSR = "ENABLED";
    FD1P3AX d_out_i0_i5 (.D(d_out_11__N_1818[5]), .SP(v_comb), .CK(osc_clk), 
            .Q(\CIC1_outSin[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i5.GSR = "ENABLED";
    FD1P3AX d_out_i0_i6 (.D(d_out_11__N_1818[6]), .SP(v_comb), .CK(osc_clk), 
            .Q(MYLED_c_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i6.GSR = "ENABLED";
    FD1P3AX d_out_i0_i7 (.D(d_out_11__N_1818[7]), .SP(v_comb), .CK(osc_clk), 
            .Q(MYLED_c_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i7.GSR = "ENABLED";
    FD1P3AX d_out_i0_i8 (.D(d_out_11__N_1818[8]), .SP(v_comb), .CK(osc_clk), 
            .Q(MYLED_c_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i8.GSR = "ENABLED";
    FD1P3AX d_out_i0_i9 (.D(d_out_11__N_1818[9]), .SP(v_comb), .CK(osc_clk), 
            .Q(MYLED_c_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i9.GSR = "ENABLED";
    FD1P3AX d_out_i0_i10 (.D(d_out_11__N_1818[10]), .SP(v_comb), .CK(osc_clk), 
            .Q(MYLED_c_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i10.GSR = "ENABLED";
    FD1P3AX d_out_i0_i11 (.D(d_out_11__N_1818[11]), .SP(v_comb), .CK(osc_clk), 
            .Q(MYLED_c_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i11.GSR = "ENABLED";
    FD1S3AX d1_i1 (.D(d1_71__N_417[1]), .CK(osc_clk), .Q(d1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i1.GSR = "ENABLED";
    FD1S3AX d1_i2 (.D(d1_71__N_417[2]), .CK(osc_clk), .Q(d1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i2.GSR = "ENABLED";
    FD1S3AX d1_i3 (.D(d1_71__N_417[3]), .CK(osc_clk), .Q(d1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i3.GSR = "ENABLED";
    FD1S3AX d1_i4 (.D(d1_71__N_417[4]), .CK(osc_clk), .Q(d1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i4.GSR = "ENABLED";
    FD1S3AX d1_i5 (.D(d1_71__N_417[5]), .CK(osc_clk), .Q(d1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i5.GSR = "ENABLED";
    FD1S3AX d1_i6 (.D(d1_71__N_417[6]), .CK(osc_clk), .Q(d1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i6.GSR = "ENABLED";
    FD1S3AX d1_i7 (.D(d1_71__N_417[7]), .CK(osc_clk), .Q(d1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i7.GSR = "ENABLED";
    FD1S3AX d1_i8 (.D(d1_71__N_417[8]), .CK(osc_clk), .Q(d1[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i8.GSR = "ENABLED";
    FD1S3AX d1_i9 (.D(d1_71__N_417[9]), .CK(osc_clk), .Q(d1[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i9.GSR = "ENABLED";
    FD1S3AX d1_i10 (.D(d1_71__N_417[10]), .CK(osc_clk), .Q(d1[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i10.GSR = "ENABLED";
    FD1S3AX d1_i11 (.D(d1_71__N_417[11]), .CK(osc_clk), .Q(d1[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i11.GSR = "ENABLED";
    FD1S3AX d1_i12 (.D(d1_71__N_417[12]), .CK(osc_clk), .Q(d1[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i12.GSR = "ENABLED";
    FD1S3AX d1_i13 (.D(d1_71__N_417[13]), .CK(osc_clk), .Q(d1[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i13.GSR = "ENABLED";
    FD1S3AX d1_i14 (.D(d1_71__N_417[14]), .CK(osc_clk), .Q(d1[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i14.GSR = "ENABLED";
    FD1S3AX d1_i15 (.D(d1_71__N_417[15]), .CK(osc_clk), .Q(d1[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i15.GSR = "ENABLED";
    FD1S3AX d1_i16 (.D(d1_71__N_417[16]), .CK(osc_clk), .Q(d1[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i16.GSR = "ENABLED";
    FD1S3AX d1_i17 (.D(d1_71__N_417[17]), .CK(osc_clk), .Q(d1[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i17.GSR = "ENABLED";
    FD1S3AX d1_i18 (.D(d1_71__N_417[18]), .CK(osc_clk), .Q(d1[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i18.GSR = "ENABLED";
    FD1S3AX d1_i19 (.D(d1_71__N_417[19]), .CK(osc_clk), .Q(d1[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i19.GSR = "ENABLED";
    FD1S3AX d1_i20 (.D(d1_71__N_417[20]), .CK(osc_clk), .Q(d1[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i20.GSR = "ENABLED";
    FD1S3AX d1_i21 (.D(d1_71__N_417[21]), .CK(osc_clk), .Q(d1[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i21.GSR = "ENABLED";
    FD1S3AX d1_i22 (.D(d1_71__N_417[22]), .CK(osc_clk), .Q(d1[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i22.GSR = "ENABLED";
    FD1S3AX d1_i23 (.D(d1_71__N_417[23]), .CK(osc_clk), .Q(d1[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i23.GSR = "ENABLED";
    FD1S3AX d1_i24 (.D(d1_71__N_417[24]), .CK(osc_clk), .Q(d1[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i24.GSR = "ENABLED";
    FD1S3AX d1_i25 (.D(d1_71__N_417[25]), .CK(osc_clk), .Q(d1[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i25.GSR = "ENABLED";
    FD1S3AX d1_i26 (.D(d1_71__N_417[26]), .CK(osc_clk), .Q(d1[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i26.GSR = "ENABLED";
    FD1S3AX d1_i27 (.D(d1_71__N_417[27]), .CK(osc_clk), .Q(d1[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i27.GSR = "ENABLED";
    FD1S3AX d1_i28 (.D(d1_71__N_417[28]), .CK(osc_clk), .Q(d1[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i28.GSR = "ENABLED";
    FD1S3AX d1_i29 (.D(d1_71__N_417[29]), .CK(osc_clk), .Q(d1[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i29.GSR = "ENABLED";
    FD1S3AX d1_i30 (.D(d1_71__N_417[30]), .CK(osc_clk), .Q(d1[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i30.GSR = "ENABLED";
    FD1S3AX d1_i31 (.D(d1_71__N_417[31]), .CK(osc_clk), .Q(d1[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i31.GSR = "ENABLED";
    FD1S3AX d1_i32 (.D(d1_71__N_417[32]), .CK(osc_clk), .Q(d1[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i32.GSR = "ENABLED";
    FD1S3AX d1_i33 (.D(d1_71__N_417[33]), .CK(osc_clk), .Q(d1[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i33.GSR = "ENABLED";
    FD1S3AX d1_i34 (.D(d1_71__N_417[34]), .CK(osc_clk), .Q(d1[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i34.GSR = "ENABLED";
    FD1S3AX d1_i35 (.D(d1_71__N_417[35]), .CK(osc_clk), .Q(d1[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i35.GSR = "ENABLED";
    FD1S3AX d1_i36 (.D(d1_71__N_417[36]), .CK(osc_clk), .Q(d1[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i36.GSR = "ENABLED";
    FD1S3AX d1_i37 (.D(d1_71__N_417[37]), .CK(osc_clk), .Q(d1[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i37.GSR = "ENABLED";
    FD1S3AX d1_i38 (.D(d1_71__N_417[38]), .CK(osc_clk), .Q(d1[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i38.GSR = "ENABLED";
    FD1S3AX d1_i39 (.D(d1_71__N_417[39]), .CK(osc_clk), .Q(d1[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i39.GSR = "ENABLED";
    FD1S3AX d1_i40 (.D(d1_71__N_417[40]), .CK(osc_clk), .Q(d1[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i40.GSR = "ENABLED";
    FD1S3AX d1_i41 (.D(d1_71__N_417[41]), .CK(osc_clk), .Q(d1[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i41.GSR = "ENABLED";
    FD1S3AX d1_i42 (.D(d1_71__N_417[42]), .CK(osc_clk), .Q(d1[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i42.GSR = "ENABLED";
    FD1S3AX d1_i43 (.D(d1_71__N_417[43]), .CK(osc_clk), .Q(d1[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i43.GSR = "ENABLED";
    FD1S3AX d1_i44 (.D(d1_71__N_417[44]), .CK(osc_clk), .Q(d1[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i44.GSR = "ENABLED";
    FD1S3AX d1_i45 (.D(d1_71__N_417[45]), .CK(osc_clk), .Q(d1[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i45.GSR = "ENABLED";
    FD1S3AX d1_i46 (.D(d1_71__N_417[46]), .CK(osc_clk), .Q(d1[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i46.GSR = "ENABLED";
    FD1S3AX d1_i47 (.D(d1_71__N_417[47]), .CK(osc_clk), .Q(d1[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i47.GSR = "ENABLED";
    FD1S3AX d1_i48 (.D(d1_71__N_417[48]), .CK(osc_clk), .Q(d1[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i48.GSR = "ENABLED";
    FD1S3AX d1_i49 (.D(d1_71__N_417[49]), .CK(osc_clk), .Q(d1[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i49.GSR = "ENABLED";
    FD1S3AX d1_i50 (.D(d1_71__N_417[50]), .CK(osc_clk), .Q(d1[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i50.GSR = "ENABLED";
    FD1S3AX d1_i51 (.D(d1_71__N_417[51]), .CK(osc_clk), .Q(d1[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i51.GSR = "ENABLED";
    FD1S3AX d1_i52 (.D(d1_71__N_417[52]), .CK(osc_clk), .Q(d1[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i52.GSR = "ENABLED";
    FD1S3AX d1_i53 (.D(d1_71__N_417[53]), .CK(osc_clk), .Q(d1[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i53.GSR = "ENABLED";
    FD1S3AX d1_i54 (.D(d1_71__N_417[54]), .CK(osc_clk), .Q(d1[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i54.GSR = "ENABLED";
    FD1S3AX d1_i55 (.D(d1_71__N_417[55]), .CK(osc_clk), .Q(d1[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i55.GSR = "ENABLED";
    FD1S3AX d1_i56 (.D(d1_71__N_417[56]), .CK(osc_clk), .Q(d1[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i56.GSR = "ENABLED";
    FD1S3AX d1_i57 (.D(d1_71__N_417[57]), .CK(osc_clk), .Q(d1[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i57.GSR = "ENABLED";
    FD1S3AX d1_i58 (.D(d1_71__N_417[58]), .CK(osc_clk), .Q(d1[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i58.GSR = "ENABLED";
    FD1S3AX d1_i59 (.D(d1_71__N_417[59]), .CK(osc_clk), .Q(d1[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i59.GSR = "ENABLED";
    FD1S3AX d1_i60 (.D(d1_71__N_417[60]), .CK(osc_clk), .Q(d1[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i60.GSR = "ENABLED";
    FD1S3AX d1_i61 (.D(d1_71__N_417[61]), .CK(osc_clk), .Q(d1[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i61.GSR = "ENABLED";
    FD1S3AX d1_i62 (.D(d1_71__N_417[62]), .CK(osc_clk), .Q(d1[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i62.GSR = "ENABLED";
    FD1S3AX d1_i63 (.D(d1_71__N_417[63]), .CK(osc_clk), .Q(d1[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i63.GSR = "ENABLED";
    FD1S3AX d1_i64 (.D(d1_71__N_417[64]), .CK(osc_clk), .Q(d1[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i64.GSR = "ENABLED";
    FD1S3AX d1_i65 (.D(d1_71__N_417[65]), .CK(osc_clk), .Q(d1[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i65.GSR = "ENABLED";
    FD1S3AX d1_i66 (.D(d1_71__N_417[66]), .CK(osc_clk), .Q(d1[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i66.GSR = "ENABLED";
    FD1S3AX d1_i67 (.D(d1_71__N_417[67]), .CK(osc_clk), .Q(d1[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i67.GSR = "ENABLED";
    FD1S3AX d1_i68 (.D(d1_71__N_417[68]), .CK(osc_clk), .Q(d1[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i68.GSR = "ENABLED";
    FD1S3AX d1_i69 (.D(d1_71__N_417[69]), .CK(osc_clk), .Q(d1[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i69.GSR = "ENABLED";
    FD1S3AX d1_i70 (.D(d1_71__N_417[70]), .CK(osc_clk), .Q(d1[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i70.GSR = "ENABLED";
    FD1S3AX d1_i71 (.D(d1_71__N_417[71]), .CK(osc_clk), .Q(d1[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i71.GSR = "ENABLED";
    CCU2D add_994_37 (.A0(d3[70]), .B0(n4342), .C0(n4343[34]), .D0(d2[70]), 
          .A1(d3[71]), .B1(n4342), .C1(n4343[35]), .D1(d2[71]), .CIN(n12054), 
          .S0(d3_71__N_561[70]), .S1(d3_71__N_561[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_994_37.INIT0 = 16'h74b8;
    defparam add_994_37.INIT1 = 16'h74b8;
    defparam add_994_37.INJECT1_0 = "NO";
    defparam add_994_37.INJECT1_1 = "NO";
    CCU2D add_994_35 (.A0(d3[68]), .B0(n4342), .C0(n4343[32]), .D0(d2[68]), 
          .A1(d3[69]), .B1(n4342), .C1(n4343[33]), .D1(d2[69]), .CIN(n12053), 
          .COUT(n12054), .S0(d3_71__N_561[68]), .S1(d3_71__N_561[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_994_35.INIT0 = 16'h74b8;
    defparam add_994_35.INIT1 = 16'h74b8;
    defparam add_994_35.INJECT1_0 = "NO";
    defparam add_994_35.INJECT1_1 = "NO";
    CCU2D add_994_33 (.A0(d3[66]), .B0(n4342), .C0(n4343[30]), .D0(d2[66]), 
          .A1(d3[67]), .B1(n4342), .C1(n4343[31]), .D1(d2[67]), .CIN(n12052), 
          .COUT(n12053), .S0(d3_71__N_561[66]), .S1(d3_71__N_561[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_994_33.INIT0 = 16'h74b8;
    defparam add_994_33.INIT1 = 16'h74b8;
    defparam add_994_33.INJECT1_0 = "NO";
    defparam add_994_33.INJECT1_1 = "NO";
    CCU2D add_994_31 (.A0(d3[64]), .B0(n4342), .C0(n4343[28]), .D0(d2[64]), 
          .A1(d3[65]), .B1(n4342), .C1(n4343[29]), .D1(d2[65]), .CIN(n12051), 
          .COUT(n12052), .S0(d3_71__N_561[64]), .S1(d3_71__N_561[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_994_31.INIT0 = 16'h74b8;
    defparam add_994_31.INIT1 = 16'h74b8;
    defparam add_994_31.INJECT1_0 = "NO";
    defparam add_994_31.INJECT1_1 = "NO";
    CCU2D add_994_29 (.A0(d3[62]), .B0(n4342), .C0(n4343[26]), .D0(d2[62]), 
          .A1(d3[63]), .B1(n4342), .C1(n4343[27]), .D1(d2[63]), .CIN(n12050), 
          .COUT(n12051), .S0(d3_71__N_561[62]), .S1(d3_71__N_561[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_994_29.INIT0 = 16'h74b8;
    defparam add_994_29.INIT1 = 16'h74b8;
    defparam add_994_29.INJECT1_0 = "NO";
    defparam add_994_29.INJECT1_1 = "NO";
    CCU2D add_994_27 (.A0(d3[60]), .B0(n4342), .C0(n4343[24]), .D0(d2[60]), 
          .A1(d3[61]), .B1(n4342), .C1(n4343[25]), .D1(d2[61]), .CIN(n12049), 
          .COUT(n12050), .S0(d3_71__N_561[60]), .S1(d3_71__N_561[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_994_27.INIT0 = 16'h74b8;
    defparam add_994_27.INIT1 = 16'h74b8;
    defparam add_994_27.INJECT1_0 = "NO";
    defparam add_994_27.INJECT1_1 = "NO";
    CCU2D add_994_25 (.A0(d3[58]), .B0(n4342), .C0(n4343[22]), .D0(d2[58]), 
          .A1(d3[59]), .B1(n4342), .C1(n4343[23]), .D1(d2[59]), .CIN(n12048), 
          .COUT(n12049), .S0(d3_71__N_561[58]), .S1(d3_71__N_561[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_994_25.INIT0 = 16'h74b8;
    defparam add_994_25.INIT1 = 16'h74b8;
    defparam add_994_25.INJECT1_0 = "NO";
    defparam add_994_25.INJECT1_1 = "NO";
    CCU2D add_994_23 (.A0(d3[56]), .B0(n4342), .C0(n4343[20]), .D0(d2[56]), 
          .A1(d3[57]), .B1(n4342), .C1(n4343[21]), .D1(d2[57]), .CIN(n12047), 
          .COUT(n12048), .S0(d3_71__N_561[56]), .S1(d3_71__N_561[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_994_23.INIT0 = 16'h74b8;
    defparam add_994_23.INIT1 = 16'h74b8;
    defparam add_994_23.INJECT1_0 = "NO";
    defparam add_994_23.INJECT1_1 = "NO";
    CCU2D add_994_21 (.A0(d3[54]), .B0(n4342), .C0(n4343[18]), .D0(d2[54]), 
          .A1(d3[55]), .B1(n4342), .C1(n4343[19]), .D1(d2[55]), .CIN(n12046), 
          .COUT(n12047), .S0(d3_71__N_561[54]), .S1(d3_71__N_561[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_994_21.INIT0 = 16'h74b8;
    defparam add_994_21.INIT1 = 16'h74b8;
    defparam add_994_21.INJECT1_0 = "NO";
    defparam add_994_21.INJECT1_1 = "NO";
    CCU2D add_994_19 (.A0(d3[52]), .B0(n4342), .C0(n4343[16]), .D0(d2[52]), 
          .A1(d3[53]), .B1(n4342), .C1(n4343[17]), .D1(d2[53]), .CIN(n12045), 
          .COUT(n12046), .S0(d3_71__N_561[52]), .S1(d3_71__N_561[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_994_19.INIT0 = 16'h74b8;
    defparam add_994_19.INIT1 = 16'h74b8;
    defparam add_994_19.INJECT1_0 = "NO";
    defparam add_994_19.INJECT1_1 = "NO";
    CCU2D add_994_17 (.A0(d3[50]), .B0(n4342), .C0(n4343[14]), .D0(d2[50]), 
          .A1(d3[51]), .B1(n4342), .C1(n4343[15]), .D1(d2[51]), .CIN(n12044), 
          .COUT(n12045), .S0(d3_71__N_561[50]), .S1(d3_71__N_561[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_994_17.INIT0 = 16'h74b8;
    defparam add_994_17.INIT1 = 16'h74b8;
    defparam add_994_17.INJECT1_0 = "NO";
    defparam add_994_17.INJECT1_1 = "NO";
    CCU2D add_994_15 (.A0(d3[48]), .B0(n4342), .C0(n4343[12]), .D0(d2[48]), 
          .A1(d3[49]), .B1(n4342), .C1(n4343[13]), .D1(d2[49]), .CIN(n12043), 
          .COUT(n12044), .S0(d3_71__N_561[48]), .S1(d3_71__N_561[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_994_15.INIT0 = 16'h74b8;
    defparam add_994_15.INIT1 = 16'h74b8;
    defparam add_994_15.INJECT1_0 = "NO";
    defparam add_994_15.INJECT1_1 = "NO";
    FD1S3IX count__i2 (.D(n375[2]), .CK(osc_clk), .CD(n8367), .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n375[3]), .CK(osc_clk), .CD(n8367), .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n375[4]), .CK(osc_clk), .CD(n8367), .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n375[5]), .CK(osc_clk), .CD(n8367), .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n375[6]), .CK(osc_clk), .CD(n8367), .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n375[7]), .CK(osc_clk), .CD(n8367), .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n375[8]), .CK(osc_clk), .CD(n8367), .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n375[9]), .CK(osc_clk), .CD(n8367), .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n375[10]), .CK(osc_clk), .CD(n8367), .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_15__N_1441[11]), .CK(osc_clk), .CD(d_clk_tmp_N_1830), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(n375[12]), .CK(osc_clk), .CD(n8367), .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(n375[13]), .CK(osc_clk), .CD(n8367), .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(n375[14]), .CK(osc_clk), .CD(n8367), .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(n375[15]), .CK(osc_clk), .CD(n8367), .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i15.GSR = "ENABLED";
    CCU2D add_982_32 (.A0(MixerOutSin[11]), .B0(d1[30]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12258), .COUT(n12259), .S0(d1_71__N_417[30]), 
          .S1(d1_71__N_417[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_982_32.INIT0 = 16'h5666;
    defparam add_982_32.INIT1 = 16'h5666;
    defparam add_982_32.INJECT1_0 = "NO";
    defparam add_982_32.INJECT1_1 = "NO";
    FD1P3AX d_d_tmp_i0_i5 (.D(d_tmp[5]), .SP(osc_clk_enable_1395), .CK(osc_clk), 
            .Q(d_d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i5.GSR = "ENABLED";
    LUT4 i9_4_lut (.A(count[9]), .B(count[3]), .C(count[4]), .D(count[0]), 
         .Z(n21)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(80[22:52])
    defparam i9_4_lut.init = 16'hfffe;
    CCU2D add_982_30 (.A0(MixerOutSin[11]), .B0(d1[28]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12257), .COUT(n12258), .S0(d1_71__N_417[28]), 
          .S1(d1_71__N_417[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_982_30.INIT0 = 16'h5666;
    defparam add_982_30.INIT1 = 16'h5666;
    defparam add_982_30.INJECT1_0 = "NO";
    defparam add_982_30.INJECT1_1 = "NO";
    CCU2D add_982_28 (.A0(MixerOutSin[11]), .B0(d1[26]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12256), .COUT(n12257), .S0(d1_71__N_417[26]), 
          .S1(d1_71__N_417[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_982_28.INIT0 = 16'h5666;
    defparam add_982_28.INIT1 = 16'h5666;
    defparam add_982_28.INJECT1_0 = "NO";
    defparam add_982_28.INJECT1_1 = "NO";
    CCU2D add_1058_37 (.A0(d9[71]), .B0(d_d9[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11408), 
          .S0(n6319[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1058_37.INIT0 = 16'h5999;
    defparam add_1058_37.INIT1 = 16'h0000;
    defparam add_1058_37.INJECT1_0 = "NO";
    defparam add_1058_37.INJECT1_1 = "NO";
    CCU2D add_1058_35 (.A0(d9[69]), .B0(d_d9[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[70]), .B1(d_d9[70]), .C1(GND_net), .D1(GND_net), .CIN(n11407), 
          .COUT(n11408), .S0(n6319[33]), .S1(n6319[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1058_35.INIT0 = 16'h5999;
    defparam add_1058_35.INIT1 = 16'h5999;
    defparam add_1058_35.INJECT1_0 = "NO";
    defparam add_1058_35.INJECT1_1 = "NO";
    CCU2D add_1058_33 (.A0(d9[67]), .B0(d_d9[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[68]), .B1(d_d9[68]), .C1(GND_net), .D1(GND_net), .CIN(n11406), 
          .COUT(n11407), .S0(n6319[31]), .S1(n6319[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1058_33.INIT0 = 16'h5999;
    defparam add_1058_33.INIT1 = 16'h5999;
    defparam add_1058_33.INJECT1_0 = "NO";
    defparam add_1058_33.INJECT1_1 = "NO";
    CCU2D add_1058_31 (.A0(d9[65]), .B0(d_d9[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[66]), .B1(d_d9[66]), .C1(GND_net), .D1(GND_net), .CIN(n11405), 
          .COUT(n11406), .S0(n6319[29]), .S1(n6319[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1058_31.INIT0 = 16'h5999;
    defparam add_1058_31.INIT1 = 16'h5999;
    defparam add_1058_31.INJECT1_0 = "NO";
    defparam add_1058_31.INJECT1_1 = "NO";
    CCU2D add_1058_29 (.A0(d9[63]), .B0(d_d9[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[64]), .B1(d_d9[64]), .C1(GND_net), .D1(GND_net), .CIN(n11404), 
          .COUT(n11405), .S0(n6319[27]), .S1(n6319[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1058_29.INIT0 = 16'h5999;
    defparam add_1058_29.INIT1 = 16'h5999;
    defparam add_1058_29.INJECT1_0 = "NO";
    defparam add_1058_29.INJECT1_1 = "NO";
    CCU2D add_1058_27 (.A0(d9[61]), .B0(d_d9[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[62]), .B1(d_d9[62]), .C1(GND_net), .D1(GND_net), .CIN(n11403), 
          .COUT(n11404), .S0(n6319[25]), .S1(n6319[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1058_27.INIT0 = 16'h5999;
    defparam add_1058_27.INIT1 = 16'h5999;
    defparam add_1058_27.INJECT1_0 = "NO";
    defparam add_1058_27.INJECT1_1 = "NO";
    CCU2D add_1058_25 (.A0(d9[59]), .B0(d_d9[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[60]), .B1(d_d9[60]), .C1(GND_net), .D1(GND_net), .CIN(n11402), 
          .COUT(n11403), .S0(n6319[23]), .S1(n6319[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1058_25.INIT0 = 16'h5999;
    defparam add_1058_25.INIT1 = 16'h5999;
    defparam add_1058_25.INJECT1_0 = "NO";
    defparam add_1058_25.INJECT1_1 = "NO";
    CCU2D add_1058_23 (.A0(d9[57]), .B0(d_d9[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[58]), .B1(d_d9[58]), .C1(GND_net), .D1(GND_net), .CIN(n11401), 
          .COUT(n11402), .S0(n6319[21]), .S1(n6319[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1058_23.INIT0 = 16'h5999;
    defparam add_1058_23.INIT1 = 16'h5999;
    defparam add_1058_23.INJECT1_0 = "NO";
    defparam add_1058_23.INJECT1_1 = "NO";
    CCU2D add_1058_21 (.A0(d9[55]), .B0(d_d9[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[56]), .B1(d_d9[56]), .C1(GND_net), .D1(GND_net), .CIN(n11400), 
          .COUT(n11401));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1058_21.INIT0 = 16'h5999;
    defparam add_1058_21.INIT1 = 16'h5999;
    defparam add_1058_21.INJECT1_0 = "NO";
    defparam add_1058_21.INJECT1_1 = "NO";
    CCU2D add_1058_19 (.A0(d9[53]), .B0(d_d9[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[54]), .B1(d_d9[54]), .C1(GND_net), .D1(GND_net), .CIN(n11399), 
          .COUT(n11400));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1058_19.INIT0 = 16'h5999;
    defparam add_1058_19.INIT1 = 16'h5999;
    defparam add_1058_19.INJECT1_0 = "NO";
    defparam add_1058_19.INJECT1_1 = "NO";
    CCU2D add_1058_17 (.A0(d9[51]), .B0(d_d9[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[52]), .B1(d_d9[52]), .C1(GND_net), .D1(GND_net), .CIN(n11398), 
          .COUT(n11399));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1058_17.INIT0 = 16'h5999;
    defparam add_1058_17.INIT1 = 16'h5999;
    defparam add_1058_17.INJECT1_0 = "NO";
    defparam add_1058_17.INJECT1_1 = "NO";
    CCU2D add_1058_15 (.A0(d9[49]), .B0(d_d9[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[50]), .B1(d_d9[50]), .C1(GND_net), .D1(GND_net), .CIN(n11397), 
          .COUT(n11398));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1058_15.INIT0 = 16'h5999;
    defparam add_1058_15.INIT1 = 16'h5999;
    defparam add_1058_15.INJECT1_0 = "NO";
    defparam add_1058_15.INJECT1_1 = "NO";
    CCU2D add_1058_13 (.A0(d9[47]), .B0(d_d9[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[48]), .B1(d_d9[48]), .C1(GND_net), .D1(GND_net), .CIN(n11396), 
          .COUT(n11397));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1058_13.INIT0 = 16'h5999;
    defparam add_1058_13.INIT1 = 16'h5999;
    defparam add_1058_13.INJECT1_0 = "NO";
    defparam add_1058_13.INJECT1_1 = "NO";
    CCU2D add_1058_11 (.A0(d9[45]), .B0(d_d9[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[46]), .B1(d_d9[46]), .C1(GND_net), .D1(GND_net), .CIN(n11395), 
          .COUT(n11396));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1058_11.INIT0 = 16'h5999;
    defparam add_1058_11.INIT1 = 16'h5999;
    defparam add_1058_11.INJECT1_0 = "NO";
    defparam add_1058_11.INJECT1_1 = "NO";
    CCU2D add_1058_9 (.A0(d9[43]), .B0(d_d9[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[44]), .B1(d_d9[44]), .C1(GND_net), .D1(GND_net), .CIN(n11394), 
          .COUT(n11395));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1058_9.INIT0 = 16'h5999;
    defparam add_1058_9.INIT1 = 16'h5999;
    defparam add_1058_9.INJECT1_0 = "NO";
    defparam add_1058_9.INJECT1_1 = "NO";
    CCU2D add_1058_7 (.A0(d9[41]), .B0(d_d9[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[42]), .B1(d_d9[42]), .C1(GND_net), .D1(GND_net), .CIN(n11393), 
          .COUT(n11394));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1058_7.INIT0 = 16'h5999;
    defparam add_1058_7.INIT1 = 16'h5999;
    defparam add_1058_7.INJECT1_0 = "NO";
    defparam add_1058_7.INJECT1_1 = "NO";
    CCU2D add_1058_5 (.A0(d9[39]), .B0(d_d9[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[40]), .B1(d_d9[40]), .C1(GND_net), .D1(GND_net), .CIN(n11392), 
          .COUT(n11393));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1058_5.INIT0 = 16'h5999;
    defparam add_1058_5.INIT1 = 16'h5999;
    defparam add_1058_5.INJECT1_0 = "NO";
    defparam add_1058_5.INJECT1_1 = "NO";
    CCU2D add_1058_3 (.A0(d9[37]), .B0(d_d9[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[38]), .B1(d_d9[38]), .C1(GND_net), .D1(GND_net), .CIN(n11391), 
          .COUT(n11392));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1058_3.INIT0 = 16'h5999;
    defparam add_1058_3.INIT1 = 16'h5999;
    defparam add_1058_3.INJECT1_0 = "NO";
    defparam add_1058_3.INJECT1_1 = "NO";
    CCU2D add_1058_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d9[36]), .B1(d_d9[36]), .C1(GND_net), .D1(GND_net), .COUT(n11391));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1058_1.INIT0 = 16'hF000;
    defparam add_1058_1.INIT1 = 16'h5999;
    defparam add_1058_1.INJECT1_0 = "NO";
    defparam add_1058_1.INJECT1_1 = "NO";
    CCU2D add_1059_37 (.A0(d9[71]), .B0(d_d9[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11390), 
          .S0(n6357[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1059_37.INIT0 = 16'h5999;
    defparam add_1059_37.INIT1 = 16'h0000;
    defparam add_1059_37.INJECT1_0 = "NO";
    defparam add_1059_37.INJECT1_1 = "NO";
    CCU2D add_1059_35 (.A0(d9[69]), .B0(d_d9[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[70]), .B1(d_d9[70]), .C1(GND_net), .D1(GND_net), .CIN(n11389), 
          .COUT(n11390), .S0(n6357[33]), .S1(n6357[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1059_35.INIT0 = 16'h5999;
    defparam add_1059_35.INIT1 = 16'h5999;
    defparam add_1059_35.INJECT1_0 = "NO";
    defparam add_1059_35.INJECT1_1 = "NO";
    CCU2D add_1059_33 (.A0(d9[67]), .B0(d_d9[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[68]), .B1(d_d9[68]), .C1(GND_net), .D1(GND_net), .CIN(n11388), 
          .COUT(n11389), .S0(n6357[31]), .S1(n6357[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1059_33.INIT0 = 16'h5999;
    defparam add_1059_33.INIT1 = 16'h5999;
    defparam add_1059_33.INJECT1_0 = "NO";
    defparam add_1059_33.INJECT1_1 = "NO";
    CCU2D add_1059_31 (.A0(d9[65]), .B0(d_d9[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[66]), .B1(d_d9[66]), .C1(GND_net), .D1(GND_net), .CIN(n11387), 
          .COUT(n11388), .S0(n6357[29]), .S1(n6357[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1059_31.INIT0 = 16'h5999;
    defparam add_1059_31.INIT1 = 16'h5999;
    defparam add_1059_31.INJECT1_0 = "NO";
    defparam add_1059_31.INJECT1_1 = "NO";
    CCU2D add_1059_29 (.A0(d9[63]), .B0(d_d9[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[64]), .B1(d_d9[64]), .C1(GND_net), .D1(GND_net), .CIN(n11386), 
          .COUT(n11387), .S0(n6357[27]), .S1(n6357[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1059_29.INIT0 = 16'h5999;
    defparam add_1059_29.INIT1 = 16'h5999;
    defparam add_1059_29.INJECT1_0 = "NO";
    defparam add_1059_29.INJECT1_1 = "NO";
    CCU2D add_1059_27 (.A0(d9[61]), .B0(d_d9[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[62]), .B1(d_d9[62]), .C1(GND_net), .D1(GND_net), .CIN(n11385), 
          .COUT(n11386), .S0(n6357[25]), .S1(n6357[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1059_27.INIT0 = 16'h5999;
    defparam add_1059_27.INIT1 = 16'h5999;
    defparam add_1059_27.INJECT1_0 = "NO";
    defparam add_1059_27.INJECT1_1 = "NO";
    CCU2D add_1059_25 (.A0(d9[59]), .B0(d_d9[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[60]), .B1(d_d9[60]), .C1(GND_net), .D1(GND_net), .CIN(n11384), 
          .COUT(n11385), .S0(n6357[23]), .S1(n6357[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1059_25.INIT0 = 16'h5999;
    defparam add_1059_25.INIT1 = 16'h5999;
    defparam add_1059_25.INJECT1_0 = "NO";
    defparam add_1059_25.INJECT1_1 = "NO";
    CCU2D add_1059_23 (.A0(d9[57]), .B0(d_d9[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[58]), .B1(d_d9[58]), .C1(GND_net), .D1(GND_net), .CIN(n11383), 
          .COUT(n11384), .S0(n6357[21]), .S1(n6357[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1059_23.INIT0 = 16'h5999;
    defparam add_1059_23.INIT1 = 16'h5999;
    defparam add_1059_23.INJECT1_0 = "NO";
    defparam add_1059_23.INJECT1_1 = "NO";
    CCU2D add_1059_21 (.A0(d9[55]), .B0(d_d9[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[56]), .B1(d_d9[56]), .C1(GND_net), .D1(GND_net), .CIN(n11382), 
          .COUT(n11383));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1059_21.INIT0 = 16'h5999;
    defparam add_1059_21.INIT1 = 16'h5999;
    defparam add_1059_21.INJECT1_0 = "NO";
    defparam add_1059_21.INJECT1_1 = "NO";
    CCU2D add_1059_19 (.A0(d9[53]), .B0(d_d9[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[54]), .B1(d_d9[54]), .C1(GND_net), .D1(GND_net), .CIN(n11381), 
          .COUT(n11382));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1059_19.INIT0 = 16'h5999;
    defparam add_1059_19.INIT1 = 16'h5999;
    defparam add_1059_19.INJECT1_0 = "NO";
    defparam add_1059_19.INJECT1_1 = "NO";
    CCU2D add_1059_17 (.A0(d9[51]), .B0(d_d9[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[52]), .B1(d_d9[52]), .C1(GND_net), .D1(GND_net), .CIN(n11380), 
          .COUT(n11381));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1059_17.INIT0 = 16'h5999;
    defparam add_1059_17.INIT1 = 16'h5999;
    defparam add_1059_17.INJECT1_0 = "NO";
    defparam add_1059_17.INJECT1_1 = "NO";
    CCU2D add_1059_15 (.A0(d9[49]), .B0(d_d9[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[50]), .B1(d_d9[50]), .C1(GND_net), .D1(GND_net), .CIN(n11379), 
          .COUT(n11380));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1059_15.INIT0 = 16'h5999;
    defparam add_1059_15.INIT1 = 16'h5999;
    defparam add_1059_15.INJECT1_0 = "NO";
    defparam add_1059_15.INJECT1_1 = "NO";
    CCU2D add_1059_13 (.A0(d9[47]), .B0(d_d9[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[48]), .B1(d_d9[48]), .C1(GND_net), .D1(GND_net), .CIN(n11378), 
          .COUT(n11379));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1059_13.INIT0 = 16'h5999;
    defparam add_1059_13.INIT1 = 16'h5999;
    defparam add_1059_13.INJECT1_0 = "NO";
    defparam add_1059_13.INJECT1_1 = "NO";
    CCU2D add_1059_11 (.A0(d9[45]), .B0(d_d9[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[46]), .B1(d_d9[46]), .C1(GND_net), .D1(GND_net), .CIN(n11377), 
          .COUT(n11378));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1059_11.INIT0 = 16'h5999;
    defparam add_1059_11.INIT1 = 16'h5999;
    defparam add_1059_11.INJECT1_0 = "NO";
    defparam add_1059_11.INJECT1_1 = "NO";
    CCU2D add_1059_9 (.A0(d9[43]), .B0(d_d9[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[44]), .B1(d_d9[44]), .C1(GND_net), .D1(GND_net), .CIN(n11376), 
          .COUT(n11377));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1059_9.INIT0 = 16'h5999;
    defparam add_1059_9.INIT1 = 16'h5999;
    defparam add_1059_9.INJECT1_0 = "NO";
    defparam add_1059_9.INJECT1_1 = "NO";
    CCU2D add_1059_7 (.A0(d9[41]), .B0(d_d9[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[42]), .B1(d_d9[42]), .C1(GND_net), .D1(GND_net), .CIN(n11375), 
          .COUT(n11376));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1059_7.INIT0 = 16'h5999;
    defparam add_1059_7.INIT1 = 16'h5999;
    defparam add_1059_7.INJECT1_0 = "NO";
    defparam add_1059_7.INJECT1_1 = "NO";
    CCU2D add_1059_5 (.A0(d9[39]), .B0(d_d9[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[40]), .B1(d_d9[40]), .C1(GND_net), .D1(GND_net), .CIN(n11374), 
          .COUT(n11375));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1059_5.INIT0 = 16'h5999;
    defparam add_1059_5.INIT1 = 16'h5999;
    defparam add_1059_5.INJECT1_0 = "NO";
    defparam add_1059_5.INJECT1_1 = "NO";
    CCU2D add_1059_3 (.A0(d9[37]), .B0(d_d9[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[38]), .B1(d_d9[38]), .C1(GND_net), .D1(GND_net), .CIN(n11373), 
          .COUT(n11374));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1059_3.INIT0 = 16'h5999;
    defparam add_1059_3.INIT1 = 16'h5999;
    defparam add_1059_3.INJECT1_0 = "NO";
    defparam add_1059_3.INJECT1_1 = "NO";
    CCU2D add_1059_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d9[36]), .B1(d_d9[36]), .C1(GND_net), .D1(GND_net), .COUT(n11373));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1059_1.INIT0 = 16'h0000;
    defparam add_1059_1.INIT1 = 16'h5999;
    defparam add_1059_1.INJECT1_0 = "NO";
    defparam add_1059_1.INJECT1_1 = "NO";
    CCU2D add_1063_37 (.A0(d8[71]), .B0(d_d8[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11372), 
          .S0(n6471[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1063_37.INIT0 = 16'h5999;
    defparam add_1063_37.INIT1 = 16'h0000;
    defparam add_1063_37.INJECT1_0 = "NO";
    defparam add_1063_37.INJECT1_1 = "NO";
    CCU2D add_1063_35 (.A0(d8[69]), .B0(d_d8[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[70]), .B1(d_d8[70]), .C1(GND_net), .D1(GND_net), .CIN(n11371), 
          .COUT(n11372), .S0(n6471[33]), .S1(n6471[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1063_35.INIT0 = 16'h5999;
    defparam add_1063_35.INIT1 = 16'h5999;
    defparam add_1063_35.INJECT1_0 = "NO";
    defparam add_1063_35.INJECT1_1 = "NO";
    CCU2D add_1063_33 (.A0(d8[67]), .B0(d_d8[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[68]), .B1(d_d8[68]), .C1(GND_net), .D1(GND_net), .CIN(n11370), 
          .COUT(n11371), .S0(n6471[31]), .S1(n6471[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1063_33.INIT0 = 16'h5999;
    defparam add_1063_33.INIT1 = 16'h5999;
    defparam add_1063_33.INJECT1_0 = "NO";
    defparam add_1063_33.INJECT1_1 = "NO";
    CCU2D add_1063_31 (.A0(d8[65]), .B0(d_d8[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[66]), .B1(d_d8[66]), .C1(GND_net), .D1(GND_net), .CIN(n11369), 
          .COUT(n11370), .S0(n6471[29]), .S1(n6471[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1063_31.INIT0 = 16'h5999;
    defparam add_1063_31.INIT1 = 16'h5999;
    defparam add_1063_31.INJECT1_0 = "NO";
    defparam add_1063_31.INJECT1_1 = "NO";
    CCU2D add_1063_29 (.A0(d8[63]), .B0(d_d8[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[64]), .B1(d_d8[64]), .C1(GND_net), .D1(GND_net), .CIN(n11368), 
          .COUT(n11369), .S0(n6471[27]), .S1(n6471[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1063_29.INIT0 = 16'h5999;
    defparam add_1063_29.INIT1 = 16'h5999;
    defparam add_1063_29.INJECT1_0 = "NO";
    defparam add_1063_29.INJECT1_1 = "NO";
    CCU2D add_1063_27 (.A0(d8[61]), .B0(d_d8[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[62]), .B1(d_d8[62]), .C1(GND_net), .D1(GND_net), .CIN(n11367), 
          .COUT(n11368), .S0(n6471[25]), .S1(n6471[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1063_27.INIT0 = 16'h5999;
    defparam add_1063_27.INIT1 = 16'h5999;
    defparam add_1063_27.INJECT1_0 = "NO";
    defparam add_1063_27.INJECT1_1 = "NO";
    CCU2D add_1063_25 (.A0(d8[59]), .B0(d_d8[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[60]), .B1(d_d8[60]), .C1(GND_net), .D1(GND_net), .CIN(n11366), 
          .COUT(n11367), .S0(n6471[23]), .S1(n6471[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1063_25.INIT0 = 16'h5999;
    defparam add_1063_25.INIT1 = 16'h5999;
    defparam add_1063_25.INJECT1_0 = "NO";
    defparam add_1063_25.INJECT1_1 = "NO";
    CCU2D add_1063_23 (.A0(d8[57]), .B0(d_d8[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[58]), .B1(d_d8[58]), .C1(GND_net), .D1(GND_net), .CIN(n11365), 
          .COUT(n11366), .S0(n6471[21]), .S1(n6471[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1063_23.INIT0 = 16'h5999;
    defparam add_1063_23.INIT1 = 16'h5999;
    defparam add_1063_23.INJECT1_0 = "NO";
    defparam add_1063_23.INJECT1_1 = "NO";
    CCU2D add_1063_21 (.A0(d8[55]), .B0(d_d8[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[56]), .B1(d_d8[56]), .C1(GND_net), .D1(GND_net), .CIN(n11364), 
          .COUT(n11365), .S0(n6471[19]), .S1(n6471[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1063_21.INIT0 = 16'h5999;
    defparam add_1063_21.INIT1 = 16'h5999;
    defparam add_1063_21.INJECT1_0 = "NO";
    defparam add_1063_21.INJECT1_1 = "NO";
    CCU2D add_1063_19 (.A0(d8[53]), .B0(d_d8[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[54]), .B1(d_d8[54]), .C1(GND_net), .D1(GND_net), .CIN(n11363), 
          .COUT(n11364), .S0(n6471[17]), .S1(n6471[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1063_19.INIT0 = 16'h5999;
    defparam add_1063_19.INIT1 = 16'h5999;
    defparam add_1063_19.INJECT1_0 = "NO";
    defparam add_1063_19.INJECT1_1 = "NO";
    CCU2D add_1063_17 (.A0(d8[51]), .B0(d_d8[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[52]), .B1(d_d8[52]), .C1(GND_net), .D1(GND_net), .CIN(n11362), 
          .COUT(n11363), .S0(n6471[15]), .S1(n6471[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1063_17.INIT0 = 16'h5999;
    defparam add_1063_17.INIT1 = 16'h5999;
    defparam add_1063_17.INJECT1_0 = "NO";
    defparam add_1063_17.INJECT1_1 = "NO";
    CCU2D add_1063_15 (.A0(d8[49]), .B0(d_d8[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[50]), .B1(d_d8[50]), .C1(GND_net), .D1(GND_net), .CIN(n11361), 
          .COUT(n11362), .S0(n6471[13]), .S1(n6471[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1063_15.INIT0 = 16'h5999;
    defparam add_1063_15.INIT1 = 16'h5999;
    defparam add_1063_15.INJECT1_0 = "NO";
    defparam add_1063_15.INJECT1_1 = "NO";
    CCU2D add_1063_13 (.A0(d8[47]), .B0(d_d8[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[48]), .B1(d_d8[48]), .C1(GND_net), .D1(GND_net), .CIN(n11360), 
          .COUT(n11361), .S0(n6471[11]), .S1(n6471[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1063_13.INIT0 = 16'h5999;
    defparam add_1063_13.INIT1 = 16'h5999;
    defparam add_1063_13.INJECT1_0 = "NO";
    defparam add_1063_13.INJECT1_1 = "NO";
    CCU2D add_1063_11 (.A0(d8[45]), .B0(d_d8[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[46]), .B1(d_d8[46]), .C1(GND_net), .D1(GND_net), .CIN(n11359), 
          .COUT(n11360), .S0(n6471[9]), .S1(n6471[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1063_11.INIT0 = 16'h5999;
    defparam add_1063_11.INIT1 = 16'h5999;
    defparam add_1063_11.INJECT1_0 = "NO";
    defparam add_1063_11.INJECT1_1 = "NO";
    CCU2D add_1063_9 (.A0(d8[43]), .B0(d_d8[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[44]), .B1(d_d8[44]), .C1(GND_net), .D1(GND_net), .CIN(n11358), 
          .COUT(n11359), .S0(n6471[7]), .S1(n6471[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1063_9.INIT0 = 16'h5999;
    defparam add_1063_9.INIT1 = 16'h5999;
    defparam add_1063_9.INJECT1_0 = "NO";
    defparam add_1063_9.INJECT1_1 = "NO";
    CCU2D add_1063_7 (.A0(d8[41]), .B0(d_d8[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[42]), .B1(d_d8[42]), .C1(GND_net), .D1(GND_net), .CIN(n11357), 
          .COUT(n11358), .S0(n6471[5]), .S1(n6471[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1063_7.INIT0 = 16'h5999;
    defparam add_1063_7.INIT1 = 16'h5999;
    defparam add_1063_7.INJECT1_0 = "NO";
    defparam add_1063_7.INJECT1_1 = "NO";
    CCU2D add_994_13 (.A0(d3[46]), .B0(n4342), .C0(n4343[10]), .D0(d2[46]), 
          .A1(d3[47]), .B1(n4342), .C1(n4343[11]), .D1(d2[47]), .CIN(n12042), 
          .COUT(n12043), .S0(d3_71__N_561[46]), .S1(d3_71__N_561[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_994_13.INIT0 = 16'h74b8;
    defparam add_994_13.INIT1 = 16'h74b8;
    defparam add_994_13.INJECT1_0 = "NO";
    defparam add_994_13.INJECT1_1 = "NO";
    CCU2D add_982_26 (.A0(MixerOutSin[11]), .B0(d1[24]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12255), .COUT(n12256), .S0(d1_71__N_417[24]), 
          .S1(d1_71__N_417[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_982_26.INIT0 = 16'h5666;
    defparam add_982_26.INIT1 = 16'h5666;
    defparam add_982_26.INJECT1_0 = "NO";
    defparam add_982_26.INJECT1_1 = "NO";
    CCU2D add_1038_5 (.A0(d7[39]), .B0(d_d7[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[40]), .B1(d_d7[40]), .C1(GND_net), .D1(GND_net), .CIN(n11690), 
          .COUT(n11691), .S0(n5711[3]), .S1(n5711[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1038_5.INIT0 = 16'h5999;
    defparam add_1038_5.INIT1 = 16'h5999;
    defparam add_1038_5.INJECT1_0 = "NO";
    defparam add_1038_5.INJECT1_1 = "NO";
    CCU2D add_982_24 (.A0(MixerOutSin[11]), .B0(d1[22]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12254), .COUT(n12255), .S0(d1_71__N_417[22]), 
          .S1(d1_71__N_417[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_982_24.INIT0 = 16'h5666;
    defparam add_982_24.INIT1 = 16'h5666;
    defparam add_982_24.INJECT1_0 = "NO";
    defparam add_982_24.INJECT1_1 = "NO";
    CCU2D add_982_22 (.A0(MixerOutSin[11]), .B0(d1[20]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12253), .COUT(n12254), .S0(d1_71__N_417[20]), 
          .S1(d1_71__N_417[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_982_22.INIT0 = 16'h5666;
    defparam add_982_22.INIT1 = 16'h5666;
    defparam add_982_22.INJECT1_0 = "NO";
    defparam add_982_22.INJECT1_1 = "NO";
    CCU2D add_982_20 (.A0(MixerOutSin[11]), .B0(d1[18]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12252), .COUT(n12253), .S0(d1_71__N_417[18]), 
          .S1(d1_71__N_417[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_982_20.INIT0 = 16'h5666;
    defparam add_982_20.INIT1 = 16'h5666;
    defparam add_982_20.INJECT1_0 = "NO";
    defparam add_982_20.INJECT1_1 = "NO";
    CCU2D add_982_18 (.A0(MixerOutSin[11]), .B0(d1[16]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12251), .COUT(n12252), .S0(d1_71__N_417[16]), 
          .S1(d1_71__N_417[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_982_18.INIT0 = 16'h5666;
    defparam add_982_18.INIT1 = 16'h5666;
    defparam add_982_18.INJECT1_0 = "NO";
    defparam add_982_18.INJECT1_1 = "NO";
    CCU2D add_982_16 (.A0(MixerOutSin[11]), .B0(d1[14]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12250), .COUT(n12251), .S0(d1_71__N_417[14]), 
          .S1(d1_71__N_417[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_982_16.INIT0 = 16'h5666;
    defparam add_982_16.INIT1 = 16'h5666;
    defparam add_982_16.INJECT1_0 = "NO";
    defparam add_982_16.INJECT1_1 = "NO";
    CCU2D add_982_14 (.A0(MixerOutSin[11]), .B0(d1[12]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12249), .COUT(n12250), .S0(d1_71__N_417[12]), 
          .S1(d1_71__N_417[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_982_14.INIT0 = 16'h5666;
    defparam add_982_14.INIT1 = 16'h5666;
    defparam add_982_14.INJECT1_0 = "NO";
    defparam add_982_14.INJECT1_1 = "NO";
    CCU2D add_982_12 (.A0(MixerOutSin[10]), .B0(d1[10]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12248), .COUT(n12249), .S0(d1_71__N_417[10]), 
          .S1(d1_71__N_417[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_982_12.INIT0 = 16'h5666;
    defparam add_982_12.INIT1 = 16'h5666;
    defparam add_982_12.INJECT1_0 = "NO";
    defparam add_982_12.INJECT1_1 = "NO";
    CCU2D add_994_11 (.A0(d3[44]), .B0(n4342), .C0(n4343[8]), .D0(d2[44]), 
          .A1(d3[45]), .B1(n4342), .C1(n4343[9]), .D1(d2[45]), .CIN(n12041), 
          .COUT(n12042), .S0(d3_71__N_561[44]), .S1(d3_71__N_561[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_994_11.INIT0 = 16'h74b8;
    defparam add_994_11.INIT1 = 16'h74b8;
    defparam add_994_11.INJECT1_0 = "NO";
    defparam add_994_11.INJECT1_1 = "NO";
    CCU2D add_994_9 (.A0(d3[42]), .B0(n4342), .C0(n4343[6]), .D0(d2[42]), 
          .A1(d3[43]), .B1(n4342), .C1(n4343[7]), .D1(d2[43]), .CIN(n12040), 
          .COUT(n12041), .S0(d3_71__N_561[42]), .S1(d3_71__N_561[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_994_9.INIT0 = 16'h74b8;
    defparam add_994_9.INIT1 = 16'h74b8;
    defparam add_994_9.INJECT1_0 = "NO";
    defparam add_994_9.INJECT1_1 = "NO";
    CCU2D add_994_7 (.A0(d3[40]), .B0(n4342), .C0(n4343[4]), .D0(d2[40]), 
          .A1(d3[41]), .B1(n4342), .C1(n4343[5]), .D1(d2[41]), .CIN(n12039), 
          .COUT(n12040), .S0(d3_71__N_561[40]), .S1(d3_71__N_561[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_994_7.INIT0 = 16'h74b8;
    defparam add_994_7.INIT1 = 16'h74b8;
    defparam add_994_7.INJECT1_0 = "NO";
    defparam add_994_7.INJECT1_1 = "NO";
    CCU2D add_994_5 (.A0(d3[38]), .B0(n4342), .C0(n4343[2]), .D0(d2[38]), 
          .A1(d3[39]), .B1(n4342), .C1(n4343[3]), .D1(d2[39]), .CIN(n12038), 
          .COUT(n12039), .S0(d3_71__N_561[38]), .S1(d3_71__N_561[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_994_5.INIT0 = 16'h74b8;
    defparam add_994_5.INIT1 = 16'h74b8;
    defparam add_994_5.INJECT1_0 = "NO";
    defparam add_994_5.INJECT1_1 = "NO";
    CCU2D add_994_3 (.A0(d3[36]), .B0(n4342), .C0(n4343[0]), .D0(d2[36]), 
          .A1(d3[37]), .B1(n4342), .C1(n4343[1]), .D1(d2[37]), .CIN(n12037), 
          .COUT(n12038), .S0(d3_71__N_561[36]), .S1(d3_71__N_561[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_994_3.INIT0 = 16'h74b8;
    defparam add_994_3.INIT1 = 16'h74b8;
    defparam add_994_3.INJECT1_0 = "NO";
    defparam add_994_3.INJECT1_1 = "NO";
    CCU2D add_994_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n4342), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n12037));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_994_1.INIT0 = 16'hF000;
    defparam add_994_1.INIT1 = 16'h0555;
    defparam add_994_1.INJECT1_0 = "NO";
    defparam add_994_1.INJECT1_1 = "NO";
    CCU2D add_998_36 (.A0(d3[70]), .B0(d4[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[71]), .B1(d4[71]), .C1(GND_net), .D1(GND_net), .CIN(n12032), 
          .S0(n4495[34]), .S1(n4495[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_998_36.INIT0 = 16'h5666;
    defparam add_998_36.INIT1 = 16'h5666;
    defparam add_998_36.INJECT1_0 = "NO";
    defparam add_998_36.INJECT1_1 = "NO";
    CCU2D add_998_34 (.A0(d3[68]), .B0(d4[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[69]), .B1(d4[69]), .C1(GND_net), .D1(GND_net), .CIN(n12031), 
          .COUT(n12032), .S0(n4495[32]), .S1(n4495[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_998_34.INIT0 = 16'h5666;
    defparam add_998_34.INIT1 = 16'h5666;
    defparam add_998_34.INJECT1_0 = "NO";
    defparam add_998_34.INJECT1_1 = "NO";
    CCU2D add_982_10 (.A0(MixerOutSin[8]), .B0(d1[8]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutSin[9]), .B1(d1[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n12247), .COUT(n12248), .S0(d1_71__N_417[8]), .S1(d1_71__N_417[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_982_10.INIT0 = 16'h5666;
    defparam add_982_10.INIT1 = 16'h5666;
    defparam add_982_10.INJECT1_0 = "NO";
    defparam add_982_10.INJECT1_1 = "NO";
    CCU2D add_982_8 (.A0(MixerOutSin[6]), .B0(d1[6]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutSin[7]), .B1(d1[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n12246), .COUT(n12247), .S0(d1_71__N_417[6]), .S1(d1_71__N_417[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_982_8.INIT0 = 16'h5666;
    defparam add_982_8.INIT1 = 16'h5666;
    defparam add_982_8.INJECT1_0 = "NO";
    defparam add_982_8.INJECT1_1 = "NO";
    LUT4 i11_3_lut_4_lut_else_3_lut (.A(\CICGain[0] ), .B(d10[69]), .C(d10[70]), 
         .Z(n13777)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam i11_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 i2_2_lut (.A(count[13]), .B(count[12]), .Z(n7)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    CCU2D add_982_6 (.A0(MixerOutSin[4]), .B0(d1[4]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutSin[5]), .B1(d1[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n12245), .COUT(n12246), .S0(d1_71__N_417[4]), .S1(d1_71__N_417[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_982_6.INIT0 = 16'h5666;
    defparam add_982_6.INIT1 = 16'h5666;
    defparam add_982_6.INJECT1_0 = "NO";
    defparam add_982_6.INJECT1_1 = "NO";
    CCU2D add_982_4 (.A0(MixerOutSin[2]), .B0(d1[2]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutSin[3]), .B1(d1[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n12244), .COUT(n12245), .S0(d1_71__N_417[2]), .S1(d1_71__N_417[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_982_4.INIT0 = 16'h5666;
    defparam add_982_4.INIT1 = 16'h5666;
    defparam add_982_4.INJECT1_0 = "NO";
    defparam add_982_4.INJECT1_1 = "NO";
    CCU2D add_998_32 (.A0(d3[66]), .B0(d4[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[67]), .B1(d4[67]), .C1(GND_net), .D1(GND_net), .CIN(n12030), 
          .COUT(n12031), .S0(n4495[30]), .S1(n4495[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_998_32.INIT0 = 16'h5666;
    defparam add_998_32.INIT1 = 16'h5666;
    defparam add_998_32.INJECT1_0 = "NO";
    defparam add_998_32.INJECT1_1 = "NO";
    CCU2D add_982_2 (.A0(MixerOutSin[0]), .B0(d1[0]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutSin[1]), .B1(d1[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n12244), .S1(d1_71__N_417[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_982_2.INIT0 = 16'h7000;
    defparam add_982_2.INIT1 = 16'h5666;
    defparam add_982_2.INJECT1_0 = "NO";
    defparam add_982_2.INJECT1_1 = "NO";
    CCU2D add_1038_3 (.A0(d7[37]), .B0(d_d7[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[38]), .B1(d_d7[38]), .C1(GND_net), .D1(GND_net), .CIN(n11689), 
          .COUT(n11690), .S0(n5711[1]), .S1(n5711[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1038_3.INIT0 = 16'h5999;
    defparam add_1038_3.INIT1 = 16'h5999;
    defparam add_1038_3.INJECT1_0 = "NO";
    defparam add_1038_3.INJECT1_1 = "NO";
    CCU2D add_1038_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d7[36]), .B1(d_d7[36]), .C1(GND_net), .D1(GND_net), .COUT(n11689), 
          .S1(n5711[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1038_1.INIT0 = 16'hF000;
    defparam add_1038_1.INIT1 = 16'h5999;
    defparam add_1038_1.INJECT1_0 = "NO";
    defparam add_1038_1.INJECT1_1 = "NO";
    CCU2D add_998_30 (.A0(d3[64]), .B0(d4[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[65]), .B1(d4[65]), .C1(GND_net), .D1(GND_net), .CIN(n12029), 
          .COUT(n12030), .S0(n4495[28]), .S1(n4495[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_998_30.INIT0 = 16'h5666;
    defparam add_998_30.INIT1 = 16'h5666;
    defparam add_998_30.INJECT1_0 = "NO";
    defparam add_998_30.INJECT1_1 = "NO";
    CCU2D add_1039_37 (.A0(d_d7[70]), .B0(n5710), .C0(n5711[34]), .D0(d7[70]), 
          .A1(d_d7[71]), .B1(n5710), .C1(n5711[35]), .D1(d7[71]), .CIN(n11687), 
          .S0(d8_71__N_1602[70]), .S1(d8_71__N_1602[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1039_37.INIT0 = 16'hb874;
    defparam add_1039_37.INIT1 = 16'hb874;
    defparam add_1039_37.INJECT1_0 = "NO";
    defparam add_1039_37.INJECT1_1 = "NO";
    CCU2D add_1039_35 (.A0(d_d7[68]), .B0(n5710), .C0(n5711[32]), .D0(d7[68]), 
          .A1(d_d7[69]), .B1(n5710), .C1(n5711[33]), .D1(d7[69]), .CIN(n11686), 
          .COUT(n11687), .S0(d8_71__N_1602[68]), .S1(d8_71__N_1602[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1039_35.INIT0 = 16'hb874;
    defparam add_1039_35.INIT1 = 16'hb874;
    defparam add_1039_35.INJECT1_0 = "NO";
    defparam add_1039_35.INJECT1_1 = "NO";
    CCU2D add_1039_33 (.A0(d_d7[66]), .B0(n5710), .C0(n5711[30]), .D0(d7[66]), 
          .A1(d_d7[67]), .B1(n5710), .C1(n5711[31]), .D1(d7[67]), .CIN(n11685), 
          .COUT(n11686), .S0(d8_71__N_1602[66]), .S1(d8_71__N_1602[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1039_33.INIT0 = 16'hb874;
    defparam add_1039_33.INIT1 = 16'hb874;
    defparam add_1039_33.INJECT1_0 = "NO";
    defparam add_1039_33.INJECT1_1 = "NO";
    CCU2D add_998_28 (.A0(d3[62]), .B0(d4[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[63]), .B1(d4[63]), .C1(GND_net), .D1(GND_net), .CIN(n12028), 
          .COUT(n12029), .S0(n4495[26]), .S1(n4495[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_998_28.INIT0 = 16'h5666;
    defparam add_998_28.INIT1 = 16'h5666;
    defparam add_998_28.INJECT1_0 = "NO";
    defparam add_998_28.INJECT1_1 = "NO";
    CCU2D add_998_26 (.A0(d3[60]), .B0(d4[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[61]), .B1(d4[61]), .C1(GND_net), .D1(GND_net), .CIN(n12027), 
          .COUT(n12028), .S0(n4495[24]), .S1(n4495[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_998_26.INIT0 = 16'h5666;
    defparam add_998_26.INIT1 = 16'h5666;
    defparam add_998_26.INJECT1_0 = "NO";
    defparam add_998_26.INJECT1_1 = "NO";
    CCU2D add_998_24 (.A0(d3[58]), .B0(d4[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[59]), .B1(d4[59]), .C1(GND_net), .D1(GND_net), .CIN(n12026), 
          .COUT(n12027), .S0(n4495[22]), .S1(n4495[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_998_24.INIT0 = 16'h5666;
    defparam add_998_24.INIT1 = 16'h5666;
    defparam add_998_24.INJECT1_0 = "NO";
    defparam add_998_24.INJECT1_1 = "NO";
    CCU2D add_998_22 (.A0(d3[56]), .B0(d4[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[57]), .B1(d4[57]), .C1(GND_net), .D1(GND_net), .CIN(n12025), 
          .COUT(n12026), .S0(n4495[20]), .S1(n4495[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_998_22.INIT0 = 16'h5666;
    defparam add_998_22.INIT1 = 16'h5666;
    defparam add_998_22.INJECT1_0 = "NO";
    defparam add_998_22.INJECT1_1 = "NO";
    CCU2D add_998_20 (.A0(d3[54]), .B0(d4[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[55]), .B1(d4[55]), .C1(GND_net), .D1(GND_net), .CIN(n12024), 
          .COUT(n12025), .S0(n4495[18]), .S1(n4495[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_998_20.INIT0 = 16'h5666;
    defparam add_998_20.INIT1 = 16'h5666;
    defparam add_998_20.INJECT1_0 = "NO";
    defparam add_998_20.INJECT1_1 = "NO";
    CCU2D add_998_18 (.A0(d3[52]), .B0(d4[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[53]), .B1(d4[53]), .C1(GND_net), .D1(GND_net), .CIN(n12023), 
          .COUT(n12024), .S0(n4495[16]), .S1(n4495[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_998_18.INIT0 = 16'h5666;
    defparam add_998_18.INIT1 = 16'h5666;
    defparam add_998_18.INJECT1_0 = "NO";
    defparam add_998_18.INJECT1_1 = "NO";
    CCU2D add_998_16 (.A0(d3[50]), .B0(d4[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[51]), .B1(d4[51]), .C1(GND_net), .D1(GND_net), .CIN(n12022), 
          .COUT(n12023), .S0(n4495[14]), .S1(n4495[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_998_16.INIT0 = 16'h5666;
    defparam add_998_16.INIT1 = 16'h5666;
    defparam add_998_16.INJECT1_0 = "NO";
    defparam add_998_16.INJECT1_1 = "NO";
    LUT4 i4806_2_lut (.A(d4[36]), .B(d5[36]), .Z(n4647[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4806_2_lut.init = 16'h6666;
    LUT4 shift_right_31_i141_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n137), .D(d10[68]), .Z(d_out_11__N_1818[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i141_3_lut_4_lut.init = 16'hf1e0;
    CCU2D add_998_14 (.A0(d3[48]), .B0(d4[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[49]), .B1(d4[49]), .C1(GND_net), .D1(GND_net), .CIN(n12021), 
          .COUT(n12022), .S0(n4495[12]), .S1(n4495[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_998_14.INIT0 = 16'h5666;
    defparam add_998_14.INIT1 = 16'h5666;
    defparam add_998_14.INJECT1_0 = "NO";
    defparam add_998_14.INJECT1_1 = "NO";
    CCU2D add_998_12 (.A0(d3[46]), .B0(d4[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[47]), .B1(d4[47]), .C1(GND_net), .D1(GND_net), .CIN(n12020), 
          .COUT(n12021), .S0(n4495[10]), .S1(n4495[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_998_12.INIT0 = 16'h5666;
    defparam add_998_12.INIT1 = 16'h5666;
    defparam add_998_12.INJECT1_0 = "NO";
    defparam add_998_12.INJECT1_1 = "NO";
    CCU2D add_1039_31 (.A0(d_d7[64]), .B0(n5710), .C0(n5711[28]), .D0(d7[64]), 
          .A1(d_d7[65]), .B1(n5710), .C1(n5711[29]), .D1(d7[65]), .CIN(n11684), 
          .COUT(n11685), .S0(d8_71__N_1602[64]), .S1(d8_71__N_1602[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1039_31.INIT0 = 16'hb874;
    defparam add_1039_31.INIT1 = 16'hb874;
    defparam add_1039_31.INJECT1_0 = "NO";
    defparam add_1039_31.INJECT1_1 = "NO";
    CCU2D add_1039_29 (.A0(d_d7[62]), .B0(n5710), .C0(n5711[26]), .D0(d7[62]), 
          .A1(d_d7[63]), .B1(n5710), .C1(n5711[27]), .D1(d7[63]), .CIN(n11683), 
          .COUT(n11684), .S0(d8_71__N_1602[62]), .S1(d8_71__N_1602[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1039_29.INIT0 = 16'hb874;
    defparam add_1039_29.INIT1 = 16'hb874;
    defparam add_1039_29.INJECT1_0 = "NO";
    defparam add_1039_29.INJECT1_1 = "NO";
    CCU2D add_1039_27 (.A0(d_d7[60]), .B0(n5710), .C0(n5711[24]), .D0(d7[60]), 
          .A1(d_d7[61]), .B1(n5710), .C1(n5711[25]), .D1(d7[61]), .CIN(n11682), 
          .COUT(n11683), .S0(d8_71__N_1602[60]), .S1(d8_71__N_1602[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1039_27.INIT0 = 16'hb874;
    defparam add_1039_27.INIT1 = 16'hb874;
    defparam add_1039_27.INJECT1_0 = "NO";
    defparam add_1039_27.INJECT1_1 = "NO";
    CCU2D add_998_10 (.A0(d3[44]), .B0(d4[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[45]), .B1(d4[45]), .C1(GND_net), .D1(GND_net), .CIN(n12019), 
          .COUT(n12020), .S0(n4495[8]), .S1(n4495[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_998_10.INIT0 = 16'h5666;
    defparam add_998_10.INIT1 = 16'h5666;
    defparam add_998_10.INJECT1_0 = "NO";
    defparam add_998_10.INJECT1_1 = "NO";
    CCU2D add_1039_25 (.A0(d_d7[58]), .B0(n5710), .C0(n5711[22]), .D0(d7[58]), 
          .A1(d_d7[59]), .B1(n5710), .C1(n5711[23]), .D1(d7[59]), .CIN(n11681), 
          .COUT(n11682), .S0(d8_71__N_1602[58]), .S1(d8_71__N_1602[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1039_25.INIT0 = 16'hb874;
    defparam add_1039_25.INIT1 = 16'hb874;
    defparam add_1039_25.INJECT1_0 = "NO";
    defparam add_1039_25.INJECT1_1 = "NO";
    CCU2D add_1063_5 (.A0(d8[39]), .B0(d_d8[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[40]), .B1(d_d8[40]), .C1(GND_net), .D1(GND_net), .CIN(n11356), 
          .COUT(n11357), .S0(n6471[3]), .S1(n6471[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1063_5.INIT0 = 16'h5999;
    defparam add_1063_5.INIT1 = 16'h5999;
    defparam add_1063_5.INJECT1_0 = "NO";
    defparam add_1063_5.INJECT1_1 = "NO";
    CCU2D add_1063_3 (.A0(d8[37]), .B0(d_d8[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[38]), .B1(d_d8[38]), .C1(GND_net), .D1(GND_net), .CIN(n11355), 
          .COUT(n11356), .S0(n6471[1]), .S1(n6471[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1063_3.INIT0 = 16'h5999;
    defparam add_1063_3.INIT1 = 16'h5999;
    defparam add_1063_3.INJECT1_0 = "NO";
    defparam add_1063_3.INJECT1_1 = "NO";
    CCU2D add_1063_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d8[36]), .B1(d_d8[36]), .C1(GND_net), .D1(GND_net), .COUT(n11355), 
          .S1(n6471[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1063_1.INIT0 = 16'hF000;
    defparam add_1063_1.INIT1 = 16'h5999;
    defparam add_1063_1.INJECT1_0 = "NO";
    defparam add_1063_1.INJECT1_1 = "NO";
    CCU2D add_1064_37 (.A0(d_d8[70]), .B0(n6470), .C0(n6471[34]), .D0(d8[70]), 
          .A1(d_d8[71]), .B1(n6470), .C1(n6471[35]), .D1(d8[71]), .CIN(n11353), 
          .S0(d9_71__N_1674[70]), .S1(d9_71__N_1674[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1064_37.INIT0 = 16'hb874;
    defparam add_1064_37.INIT1 = 16'hb874;
    defparam add_1064_37.INJECT1_0 = "NO";
    defparam add_1064_37.INJECT1_1 = "NO";
    CCU2D add_1064_35 (.A0(d_d8[68]), .B0(n6470), .C0(n6471[32]), .D0(d8[68]), 
          .A1(d_d8[69]), .B1(n6470), .C1(n6471[33]), .D1(d8[69]), .CIN(n11352), 
          .COUT(n11353), .S0(d9_71__N_1674[68]), .S1(d9_71__N_1674[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1064_35.INIT0 = 16'hb874;
    defparam add_1064_35.INIT1 = 16'hb874;
    defparam add_1064_35.INJECT1_0 = "NO";
    defparam add_1064_35.INJECT1_1 = "NO";
    CCU2D add_1064_33 (.A0(d_d8[66]), .B0(n6470), .C0(n6471[30]), .D0(d8[66]), 
          .A1(d_d8[67]), .B1(n6470), .C1(n6471[31]), .D1(d8[67]), .CIN(n11351), 
          .COUT(n11352), .S0(d9_71__N_1674[66]), .S1(d9_71__N_1674[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1064_33.INIT0 = 16'hb874;
    defparam add_1064_33.INIT1 = 16'hb874;
    defparam add_1064_33.INJECT1_0 = "NO";
    defparam add_1064_33.INJECT1_1 = "NO";
    CCU2D add_1064_31 (.A0(d_d8[64]), .B0(n6470), .C0(n6471[28]), .D0(d8[64]), 
          .A1(d_d8[65]), .B1(n6470), .C1(n6471[29]), .D1(d8[65]), .CIN(n11350), 
          .COUT(n11351), .S0(d9_71__N_1674[64]), .S1(d9_71__N_1674[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1064_31.INIT0 = 16'hb874;
    defparam add_1064_31.INIT1 = 16'hb874;
    defparam add_1064_31.INJECT1_0 = "NO";
    defparam add_1064_31.INJECT1_1 = "NO";
    CCU2D add_1064_29 (.A0(d_d8[62]), .B0(n6470), .C0(n6471[26]), .D0(d8[62]), 
          .A1(d_d8[63]), .B1(n6470), .C1(n6471[27]), .D1(d8[63]), .CIN(n11349), 
          .COUT(n11350), .S0(d9_71__N_1674[62]), .S1(d9_71__N_1674[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1064_29.INIT0 = 16'hb874;
    defparam add_1064_29.INIT1 = 16'hb874;
    defparam add_1064_29.INJECT1_0 = "NO";
    defparam add_1064_29.INJECT1_1 = "NO";
    CCU2D add_1064_27 (.A0(d_d8[60]), .B0(n6470), .C0(n6471[24]), .D0(d8[60]), 
          .A1(d_d8[61]), .B1(n6470), .C1(n6471[25]), .D1(d8[61]), .CIN(n11348), 
          .COUT(n11349), .S0(d9_71__N_1674[60]), .S1(d9_71__N_1674[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1064_27.INIT0 = 16'hb874;
    defparam add_1064_27.INIT1 = 16'hb874;
    defparam add_1064_27.INJECT1_0 = "NO";
    defparam add_1064_27.INJECT1_1 = "NO";
    CCU2D add_1064_25 (.A0(d_d8[58]), .B0(n6470), .C0(n6471[22]), .D0(d8[58]), 
          .A1(d_d8[59]), .B1(n6470), .C1(n6471[23]), .D1(d8[59]), .CIN(n11347), 
          .COUT(n11348), .S0(d9_71__N_1674[58]), .S1(d9_71__N_1674[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1064_25.INIT0 = 16'hb874;
    defparam add_1064_25.INIT1 = 16'hb874;
    defparam add_1064_25.INJECT1_0 = "NO";
    defparam add_1064_25.INJECT1_1 = "NO";
    CCU2D add_1064_23 (.A0(d_d8[56]), .B0(n6470), .C0(n6471[20]), .D0(d8[56]), 
          .A1(d_d8[57]), .B1(n6470), .C1(n6471[21]), .D1(d8[57]), .CIN(n11346), 
          .COUT(n11347), .S0(d9_71__N_1674[56]), .S1(d9_71__N_1674[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1064_23.INIT0 = 16'hb874;
    defparam add_1064_23.INIT1 = 16'hb874;
    defparam add_1064_23.INJECT1_0 = "NO";
    defparam add_1064_23.INJECT1_1 = "NO";
    CCU2D add_1064_21 (.A0(d_d8[54]), .B0(n6470), .C0(n6471[18]), .D0(d8[54]), 
          .A1(d_d8[55]), .B1(n6470), .C1(n6471[19]), .D1(d8[55]), .CIN(n11345), 
          .COUT(n11346), .S0(d9_71__N_1674[54]), .S1(d9_71__N_1674[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1064_21.INIT0 = 16'hb874;
    defparam add_1064_21.INIT1 = 16'hb874;
    defparam add_1064_21.INJECT1_0 = "NO";
    defparam add_1064_21.INJECT1_1 = "NO";
    CCU2D add_1064_19 (.A0(d_d8[52]), .B0(n6470), .C0(n6471[16]), .D0(d8[52]), 
          .A1(d_d8[53]), .B1(n6470), .C1(n6471[17]), .D1(d8[53]), .CIN(n11344), 
          .COUT(n11345), .S0(d9_71__N_1674[52]), .S1(d9_71__N_1674[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1064_19.INIT0 = 16'hb874;
    defparam add_1064_19.INIT1 = 16'hb874;
    defparam add_1064_19.INJECT1_0 = "NO";
    defparam add_1064_19.INJECT1_1 = "NO";
    CCU2D add_1064_17 (.A0(d_d8[50]), .B0(n6470), .C0(n6471[14]), .D0(d8[50]), 
          .A1(d_d8[51]), .B1(n6470), .C1(n6471[15]), .D1(d8[51]), .CIN(n11343), 
          .COUT(n11344), .S0(d9_71__N_1674[50]), .S1(d9_71__N_1674[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1064_17.INIT0 = 16'hb874;
    defparam add_1064_17.INIT1 = 16'hb874;
    defparam add_1064_17.INJECT1_0 = "NO";
    defparam add_1064_17.INJECT1_1 = "NO";
    CCU2D add_1064_15 (.A0(d_d8[48]), .B0(n6470), .C0(n6471[12]), .D0(d8[48]), 
          .A1(d_d8[49]), .B1(n6470), .C1(n6471[13]), .D1(d8[49]), .CIN(n11342), 
          .COUT(n11343), .S0(d9_71__N_1674[48]), .S1(d9_71__N_1674[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1064_15.INIT0 = 16'hb874;
    defparam add_1064_15.INIT1 = 16'hb874;
    defparam add_1064_15.INJECT1_0 = "NO";
    defparam add_1064_15.INJECT1_1 = "NO";
    CCU2D add_1064_13 (.A0(d_d8[46]), .B0(n6470), .C0(n6471[10]), .D0(d8[46]), 
          .A1(d_d8[47]), .B1(n6470), .C1(n6471[11]), .D1(d8[47]), .CIN(n11341), 
          .COUT(n11342), .S0(d9_71__N_1674[46]), .S1(d9_71__N_1674[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1064_13.INIT0 = 16'hb874;
    defparam add_1064_13.INIT1 = 16'hb874;
    defparam add_1064_13.INJECT1_0 = "NO";
    defparam add_1064_13.INJECT1_1 = "NO";
    CCU2D add_1064_11 (.A0(d_d8[44]), .B0(n6470), .C0(n6471[8]), .D0(d8[44]), 
          .A1(d_d8[45]), .B1(n6470), .C1(n6471[9]), .D1(d8[45]), .CIN(n11340), 
          .COUT(n11341), .S0(d9_71__N_1674[44]), .S1(d9_71__N_1674[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1064_11.INIT0 = 16'hb874;
    defparam add_1064_11.INIT1 = 16'hb874;
    defparam add_1064_11.INJECT1_0 = "NO";
    defparam add_1064_11.INJECT1_1 = "NO";
    CCU2D add_1064_9 (.A0(d_d8[42]), .B0(n6470), .C0(n6471[6]), .D0(d8[42]), 
          .A1(d_d8[43]), .B1(n6470), .C1(n6471[7]), .D1(d8[43]), .CIN(n11339), 
          .COUT(n11340), .S0(d9_71__N_1674[42]), .S1(d9_71__N_1674[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1064_9.INIT0 = 16'hb874;
    defparam add_1064_9.INIT1 = 16'hb874;
    defparam add_1064_9.INJECT1_0 = "NO";
    defparam add_1064_9.INJECT1_1 = "NO";
    CCU2D add_1064_7 (.A0(d_d8[40]), .B0(n6470), .C0(n6471[4]), .D0(d8[40]), 
          .A1(d_d8[41]), .B1(n6470), .C1(n6471[5]), .D1(d8[41]), .CIN(n11338), 
          .COUT(n11339), .S0(d9_71__N_1674[40]), .S1(d9_71__N_1674[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1064_7.INIT0 = 16'hb874;
    defparam add_1064_7.INIT1 = 16'hb874;
    defparam add_1064_7.INJECT1_0 = "NO";
    defparam add_1064_7.INJECT1_1 = "NO";
    CCU2D add_1064_5 (.A0(d_d8[38]), .B0(n6470), .C0(n6471[2]), .D0(d8[38]), 
          .A1(d_d8[39]), .B1(n6470), .C1(n6471[3]), .D1(d8[39]), .CIN(n11337), 
          .COUT(n11338), .S0(d9_71__N_1674[38]), .S1(d9_71__N_1674[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1064_5.INIT0 = 16'hb874;
    defparam add_1064_5.INIT1 = 16'hb874;
    defparam add_1064_5.INJECT1_0 = "NO";
    defparam add_1064_5.INJECT1_1 = "NO";
    CCU2D add_1064_3 (.A0(d_d8[36]), .B0(n6470), .C0(n6471[0]), .D0(d8[36]), 
          .A1(d_d8[37]), .B1(n6470), .C1(n6471[1]), .D1(d8[37]), .CIN(n11336), 
          .COUT(n11337), .S0(d9_71__N_1674[36]), .S1(d9_71__N_1674[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1064_3.INIT0 = 16'hb874;
    defparam add_1064_3.INIT1 = 16'hb874;
    defparam add_1064_3.INJECT1_0 = "NO";
    defparam add_1064_3.INJECT1_1 = "NO";
    CCU2D add_1064_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n6470), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11336));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1064_1.INIT0 = 16'hF000;
    defparam add_1064_1.INIT1 = 16'h0555;
    defparam add_1064_1.INJECT1_0 = "NO";
    defparam add_1064_1.INJECT1_1 = "NO";
    CCU2D add_1078_37 (.A0(d_tmp[71]), .B0(d_d_tmp[71]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11256), .S0(n6927[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1078_37.INIT0 = 16'h5999;
    defparam add_1078_37.INIT1 = 16'h0000;
    defparam add_1078_37.INJECT1_0 = "NO";
    defparam add_1078_37.INJECT1_1 = "NO";
    CCU2D add_1078_35 (.A0(d_tmp[69]), .B0(d_d_tmp[69]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[70]), .B1(d_d_tmp[70]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11255), .COUT(n11256), .S0(n6927[33]), 
          .S1(n6927[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1078_35.INIT0 = 16'h5999;
    defparam add_1078_35.INIT1 = 16'h5999;
    defparam add_1078_35.INJECT1_0 = "NO";
    defparam add_1078_35.INJECT1_1 = "NO";
    CCU2D add_1078_33 (.A0(d_tmp[67]), .B0(d_d_tmp[67]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[68]), .B1(d_d_tmp[68]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11254), .COUT(n11255), .S0(n6927[31]), 
          .S1(n6927[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1078_33.INIT0 = 16'h5999;
    defparam add_1078_33.INIT1 = 16'h5999;
    defparam add_1078_33.INJECT1_0 = "NO";
    defparam add_1078_33.INJECT1_1 = "NO";
    CCU2D add_1078_31 (.A0(d_tmp[65]), .B0(d_d_tmp[65]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[66]), .B1(d_d_tmp[66]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11253), .COUT(n11254), .S0(n6927[29]), 
          .S1(n6927[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1078_31.INIT0 = 16'h5999;
    defparam add_1078_31.INIT1 = 16'h5999;
    defparam add_1078_31.INJECT1_0 = "NO";
    defparam add_1078_31.INJECT1_1 = "NO";
    CCU2D add_1078_29 (.A0(d_tmp[63]), .B0(d_d_tmp[63]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[64]), .B1(d_d_tmp[64]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11252), .COUT(n11253), .S0(n6927[27]), 
          .S1(n6927[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1078_29.INIT0 = 16'h5999;
    defparam add_1078_29.INIT1 = 16'h5999;
    defparam add_1078_29.INJECT1_0 = "NO";
    defparam add_1078_29.INJECT1_1 = "NO";
    CCU2D add_1078_27 (.A0(d_tmp[61]), .B0(d_d_tmp[61]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[62]), .B1(d_d_tmp[62]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11251), .COUT(n11252), .S0(n6927[25]), 
          .S1(n6927[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1078_27.INIT0 = 16'h5999;
    defparam add_1078_27.INIT1 = 16'h5999;
    defparam add_1078_27.INJECT1_0 = "NO";
    defparam add_1078_27.INJECT1_1 = "NO";
    CCU2D add_1078_25 (.A0(d_tmp[59]), .B0(d_d_tmp[59]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[60]), .B1(d_d_tmp[60]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11250), .COUT(n11251), .S0(n6927[23]), 
          .S1(n6927[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1078_25.INIT0 = 16'h5999;
    defparam add_1078_25.INIT1 = 16'h5999;
    defparam add_1078_25.INJECT1_0 = "NO";
    defparam add_1078_25.INJECT1_1 = "NO";
    CCU2D add_1078_23 (.A0(d_tmp[57]), .B0(d_d_tmp[57]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[58]), .B1(d_d_tmp[58]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11249), .COUT(n11250), .S0(n6927[21]), 
          .S1(n6927[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1078_23.INIT0 = 16'h5999;
    defparam add_1078_23.INIT1 = 16'h5999;
    defparam add_1078_23.INJECT1_0 = "NO";
    defparam add_1078_23.INJECT1_1 = "NO";
    CCU2D add_1078_21 (.A0(d_tmp[55]), .B0(d_d_tmp[55]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[56]), .B1(d_d_tmp[56]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11248), .COUT(n11249), .S0(n6927[19]), 
          .S1(n6927[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1078_21.INIT0 = 16'h5999;
    defparam add_1078_21.INIT1 = 16'h5999;
    defparam add_1078_21.INJECT1_0 = "NO";
    defparam add_1078_21.INJECT1_1 = "NO";
    CCU2D add_1078_19 (.A0(d_tmp[53]), .B0(d_d_tmp[53]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[54]), .B1(d_d_tmp[54]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11247), .COUT(n11248), .S0(n6927[17]), 
          .S1(n6927[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1078_19.INIT0 = 16'h5999;
    defparam add_1078_19.INIT1 = 16'h5999;
    defparam add_1078_19.INJECT1_0 = "NO";
    defparam add_1078_19.INJECT1_1 = "NO";
    CCU2D add_1078_17 (.A0(d_tmp[51]), .B0(d_d_tmp[51]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[52]), .B1(d_d_tmp[52]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11246), .COUT(n11247), .S0(n6927[15]), 
          .S1(n6927[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1078_17.INIT0 = 16'h5999;
    defparam add_1078_17.INIT1 = 16'h5999;
    defparam add_1078_17.INJECT1_0 = "NO";
    defparam add_1078_17.INJECT1_1 = "NO";
    CCU2D add_1078_15 (.A0(d_tmp[49]), .B0(d_d_tmp[49]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[50]), .B1(d_d_tmp[50]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11245), .COUT(n11246), .S0(n6927[13]), 
          .S1(n6927[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1078_15.INIT0 = 16'h5999;
    defparam add_1078_15.INIT1 = 16'h5999;
    defparam add_1078_15.INJECT1_0 = "NO";
    defparam add_1078_15.INJECT1_1 = "NO";
    CCU2D add_1078_13 (.A0(d_tmp[47]), .B0(d_d_tmp[47]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[48]), .B1(d_d_tmp[48]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11244), .COUT(n11245), .S0(n6927[11]), 
          .S1(n6927[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1078_13.INIT0 = 16'h5999;
    defparam add_1078_13.INIT1 = 16'h5999;
    defparam add_1078_13.INJECT1_0 = "NO";
    defparam add_1078_13.INJECT1_1 = "NO";
    CCU2D add_1078_11 (.A0(d_tmp[45]), .B0(d_d_tmp[45]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[46]), .B1(d_d_tmp[46]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11243), .COUT(n11244), .S0(n6927[9]), 
          .S1(n6927[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1078_11.INIT0 = 16'h5999;
    defparam add_1078_11.INIT1 = 16'h5999;
    defparam add_1078_11.INJECT1_0 = "NO";
    defparam add_1078_11.INJECT1_1 = "NO";
    CCU2D add_1078_9 (.A0(d_tmp[43]), .B0(d_d_tmp[43]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[44]), .B1(d_d_tmp[44]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11242), .COUT(n11243), .S0(n6927[7]), 
          .S1(n6927[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1078_9.INIT0 = 16'h5999;
    defparam add_1078_9.INIT1 = 16'h5999;
    defparam add_1078_9.INJECT1_0 = "NO";
    defparam add_1078_9.INJECT1_1 = "NO";
    CCU2D add_1078_7 (.A0(d_tmp[41]), .B0(d_d_tmp[41]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[42]), .B1(d_d_tmp[42]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11241), .COUT(n11242), .S0(n6927[5]), 
          .S1(n6927[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1078_7.INIT0 = 16'h5999;
    defparam add_1078_7.INIT1 = 16'h5999;
    defparam add_1078_7.INJECT1_0 = "NO";
    defparam add_1078_7.INJECT1_1 = "NO";
    CCU2D add_1078_5 (.A0(d_tmp[39]), .B0(d_d_tmp[39]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[40]), .B1(d_d_tmp[40]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11240), .COUT(n11241), .S0(n6927[3]), 
          .S1(n6927[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1078_5.INIT0 = 16'h5999;
    defparam add_1078_5.INIT1 = 16'h5999;
    defparam add_1078_5.INJECT1_0 = "NO";
    defparam add_1078_5.INJECT1_1 = "NO";
    CCU2D add_1078_3 (.A0(d_tmp[37]), .B0(d_d_tmp[37]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[38]), .B1(d_d_tmp[38]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11239), .COUT(n11240), .S0(n6927[1]), 
          .S1(n6927[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1078_3.INIT0 = 16'h5999;
    defparam add_1078_3.INIT1 = 16'h5999;
    defparam add_1078_3.INJECT1_0 = "NO";
    defparam add_1078_3.INJECT1_1 = "NO";
    CCU2D add_1078_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[36]), .B1(d_d_tmp[36]), .C1(GND_net), .D1(GND_net), 
          .COUT(n11239), .S1(n6927[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1078_1.INIT0 = 16'hF000;
    defparam add_1078_1.INIT1 = 16'h5999;
    defparam add_1078_1.INJECT1_0 = "NO";
    defparam add_1078_1.INJECT1_1 = "NO";
    CCU2D add_1079_37 (.A0(d_d_tmp[70]), .B0(n6926), .C0(n6927[34]), .D0(d_tmp[70]), 
          .A1(d_d_tmp[71]), .B1(n6926), .C1(n6927[35]), .D1(d_tmp[71]), 
          .CIN(n11237), .S0(d6_71__N_1458[70]), .S1(d6_71__N_1458[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1079_37.INIT0 = 16'hb874;
    defparam add_1079_37.INIT1 = 16'hb874;
    defparam add_1079_37.INJECT1_0 = "NO";
    defparam add_1079_37.INJECT1_1 = "NO";
    CCU2D add_1079_35 (.A0(d_d_tmp[68]), .B0(n6926), .C0(n6927[32]), .D0(d_tmp[68]), 
          .A1(d_d_tmp[69]), .B1(n6926), .C1(n6927[33]), .D1(d_tmp[69]), 
          .CIN(n11236), .COUT(n11237), .S0(d6_71__N_1458[68]), .S1(d6_71__N_1458[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1079_35.INIT0 = 16'hb874;
    defparam add_1079_35.INIT1 = 16'hb874;
    defparam add_1079_35.INJECT1_0 = "NO";
    defparam add_1079_35.INJECT1_1 = "NO";
    CCU2D add_1079_33 (.A0(d_d_tmp[66]), .B0(n6926), .C0(n6927[30]), .D0(d_tmp[66]), 
          .A1(d_d_tmp[67]), .B1(n6926), .C1(n6927[31]), .D1(d_tmp[67]), 
          .CIN(n11235), .COUT(n11236), .S0(d6_71__N_1458[66]), .S1(d6_71__N_1458[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1079_33.INIT0 = 16'hb874;
    defparam add_1079_33.INIT1 = 16'hb874;
    defparam add_1079_33.INJECT1_0 = "NO";
    defparam add_1079_33.INJECT1_1 = "NO";
    CCU2D add_1079_31 (.A0(d_d_tmp[64]), .B0(n6926), .C0(n6927[28]), .D0(d_tmp[64]), 
          .A1(d_d_tmp[65]), .B1(n6926), .C1(n6927[29]), .D1(d_tmp[65]), 
          .CIN(n11234), .COUT(n11235), .S0(d6_71__N_1458[64]), .S1(d6_71__N_1458[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1079_31.INIT0 = 16'hb874;
    defparam add_1079_31.INIT1 = 16'hb874;
    defparam add_1079_31.INJECT1_0 = "NO";
    defparam add_1079_31.INJECT1_1 = "NO";
    CCU2D add_1079_29 (.A0(d_d_tmp[62]), .B0(n6926), .C0(n6927[26]), .D0(d_tmp[62]), 
          .A1(d_d_tmp[63]), .B1(n6926), .C1(n6927[27]), .D1(d_tmp[63]), 
          .CIN(n11233), .COUT(n11234), .S0(d6_71__N_1458[62]), .S1(d6_71__N_1458[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1079_29.INIT0 = 16'hb874;
    defparam add_1079_29.INIT1 = 16'hb874;
    defparam add_1079_29.INJECT1_0 = "NO";
    defparam add_1079_29.INJECT1_1 = "NO";
    CCU2D add_1079_27 (.A0(d_d_tmp[60]), .B0(n6926), .C0(n6927[24]), .D0(d_tmp[60]), 
          .A1(d_d_tmp[61]), .B1(n6926), .C1(n6927[25]), .D1(d_tmp[61]), 
          .CIN(n11232), .COUT(n11233), .S0(d6_71__N_1458[60]), .S1(d6_71__N_1458[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1079_27.INIT0 = 16'hb874;
    defparam add_1079_27.INIT1 = 16'hb874;
    defparam add_1079_27.INJECT1_0 = "NO";
    defparam add_1079_27.INJECT1_1 = "NO";
    CCU2D add_1079_25 (.A0(d_d_tmp[58]), .B0(n6926), .C0(n6927[22]), .D0(d_tmp[58]), 
          .A1(d_d_tmp[59]), .B1(n6926), .C1(n6927[23]), .D1(d_tmp[59]), 
          .CIN(n11231), .COUT(n11232), .S0(d6_71__N_1458[58]), .S1(d6_71__N_1458[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1079_25.INIT0 = 16'hb874;
    defparam add_1079_25.INIT1 = 16'hb874;
    defparam add_1079_25.INJECT1_0 = "NO";
    defparam add_1079_25.INJECT1_1 = "NO";
    CCU2D add_1079_23 (.A0(d_d_tmp[56]), .B0(n6926), .C0(n6927[20]), .D0(d_tmp[56]), 
          .A1(d_d_tmp[57]), .B1(n6926), .C1(n6927[21]), .D1(d_tmp[57]), 
          .CIN(n11230), .COUT(n11231), .S0(d6_71__N_1458[56]), .S1(d6_71__N_1458[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1079_23.INIT0 = 16'hb874;
    defparam add_1079_23.INIT1 = 16'hb874;
    defparam add_1079_23.INJECT1_0 = "NO";
    defparam add_1079_23.INJECT1_1 = "NO";
    CCU2D add_1079_21 (.A0(d_d_tmp[54]), .B0(n6926), .C0(n6927[18]), .D0(d_tmp[54]), 
          .A1(d_d_tmp[55]), .B1(n6926), .C1(n6927[19]), .D1(d_tmp[55]), 
          .CIN(n11229), .COUT(n11230), .S0(d6_71__N_1458[54]), .S1(d6_71__N_1458[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1079_21.INIT0 = 16'hb874;
    defparam add_1079_21.INIT1 = 16'hb874;
    defparam add_1079_21.INJECT1_0 = "NO";
    defparam add_1079_21.INJECT1_1 = "NO";
    CCU2D add_1079_19 (.A0(d_d_tmp[52]), .B0(n6926), .C0(n6927[16]), .D0(d_tmp[52]), 
          .A1(d_d_tmp[53]), .B1(n6926), .C1(n6927[17]), .D1(d_tmp[53]), 
          .CIN(n11228), .COUT(n11229), .S0(d6_71__N_1458[52]), .S1(d6_71__N_1458[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1079_19.INIT0 = 16'hb874;
    defparam add_1079_19.INIT1 = 16'hb874;
    defparam add_1079_19.INJECT1_0 = "NO";
    defparam add_1079_19.INJECT1_1 = "NO";
    CCU2D add_1079_17 (.A0(d_d_tmp[50]), .B0(n6926), .C0(n6927[14]), .D0(d_tmp[50]), 
          .A1(d_d_tmp[51]), .B1(n6926), .C1(n6927[15]), .D1(d_tmp[51]), 
          .CIN(n11227), .COUT(n11228), .S0(d6_71__N_1458[50]), .S1(d6_71__N_1458[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1079_17.INIT0 = 16'hb874;
    defparam add_1079_17.INIT1 = 16'hb874;
    defparam add_1079_17.INJECT1_0 = "NO";
    defparam add_1079_17.INJECT1_1 = "NO";
    CCU2D add_1079_15 (.A0(d_d_tmp[48]), .B0(n6926), .C0(n6927[12]), .D0(d_tmp[48]), 
          .A1(d_d_tmp[49]), .B1(n6926), .C1(n6927[13]), .D1(d_tmp[49]), 
          .CIN(n11226), .COUT(n11227), .S0(d6_71__N_1458[48]), .S1(d6_71__N_1458[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1079_15.INIT0 = 16'hb874;
    defparam add_1079_15.INIT1 = 16'hb874;
    defparam add_1079_15.INJECT1_0 = "NO";
    defparam add_1079_15.INJECT1_1 = "NO";
    CCU2D add_1079_13 (.A0(d_d_tmp[46]), .B0(n6926), .C0(n6927[10]), .D0(d_tmp[46]), 
          .A1(d_d_tmp[47]), .B1(n6926), .C1(n6927[11]), .D1(d_tmp[47]), 
          .CIN(n11225), .COUT(n11226), .S0(d6_71__N_1458[46]), .S1(d6_71__N_1458[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1079_13.INIT0 = 16'hb874;
    defparam add_1079_13.INIT1 = 16'hb874;
    defparam add_1079_13.INJECT1_0 = "NO";
    defparam add_1079_13.INJECT1_1 = "NO";
    CCU2D add_1079_11 (.A0(d_d_tmp[44]), .B0(n6926), .C0(n6927[8]), .D0(d_tmp[44]), 
          .A1(d_d_tmp[45]), .B1(n6926), .C1(n6927[9]), .D1(d_tmp[45]), 
          .CIN(n11224), .COUT(n11225), .S0(d6_71__N_1458[44]), .S1(d6_71__N_1458[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1079_11.INIT0 = 16'hb874;
    defparam add_1079_11.INIT1 = 16'hb874;
    defparam add_1079_11.INJECT1_0 = "NO";
    defparam add_1079_11.INJECT1_1 = "NO";
    CCU2D add_1079_9 (.A0(d_d_tmp[42]), .B0(n6926), .C0(n6927[6]), .D0(d_tmp[42]), 
          .A1(d_d_tmp[43]), .B1(n6926), .C1(n6927[7]), .D1(d_tmp[43]), 
          .CIN(n11223), .COUT(n11224), .S0(d6_71__N_1458[42]), .S1(d6_71__N_1458[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1079_9.INIT0 = 16'hb874;
    defparam add_1079_9.INIT1 = 16'hb874;
    defparam add_1079_9.INJECT1_0 = "NO";
    defparam add_1079_9.INJECT1_1 = "NO";
    CCU2D add_1079_7 (.A0(d_d_tmp[40]), .B0(n6926), .C0(n6927[4]), .D0(d_tmp[40]), 
          .A1(d_d_tmp[41]), .B1(n6926), .C1(n6927[5]), .D1(d_tmp[41]), 
          .CIN(n11222), .COUT(n11223), .S0(d6_71__N_1458[40]), .S1(d6_71__N_1458[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1079_7.INIT0 = 16'hb874;
    defparam add_1079_7.INIT1 = 16'hb874;
    defparam add_1079_7.INJECT1_0 = "NO";
    defparam add_1079_7.INJECT1_1 = "NO";
    CCU2D add_1079_5 (.A0(d_d_tmp[38]), .B0(n6926), .C0(n6927[2]), .D0(d_tmp[38]), 
          .A1(d_d_tmp[39]), .B1(n6926), .C1(n6927[3]), .D1(d_tmp[39]), 
          .CIN(n11221), .COUT(n11222), .S0(d6_71__N_1458[38]), .S1(d6_71__N_1458[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1079_5.INIT0 = 16'hb874;
    defparam add_1079_5.INIT1 = 16'hb874;
    defparam add_1079_5.INJECT1_0 = "NO";
    defparam add_1079_5.INJECT1_1 = "NO";
    CCU2D add_1079_3 (.A0(d_d_tmp[36]), .B0(n6926), .C0(n6927[0]), .D0(d_tmp[36]), 
          .A1(d_d_tmp[37]), .B1(n6926), .C1(n6927[1]), .D1(d_tmp[37]), 
          .CIN(n11220), .COUT(n11221), .S0(d6_71__N_1458[36]), .S1(d6_71__N_1458[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1079_3.INIT0 = 16'hb874;
    defparam add_1079_3.INIT1 = 16'hb874;
    defparam add_1079_3.INJECT1_0 = "NO";
    defparam add_1079_3.INJECT1_1 = "NO";
    CCU2D add_1079_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n6926), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11220));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1079_1.INIT0 = 16'hF000;
    defparam add_1079_1.INIT1 = 16'h0555;
    defparam add_1079_1.INJECT1_0 = "NO";
    defparam add_1079_1.INJECT1_1 = "NO";
    CCU2D add_983_37 (.A0(d1[70]), .B0(n4038), .C0(n4077[34]), .D0(MixerOutSin[11]), 
          .A1(d1[71]), .B1(n4038), .C1(n4077[35]), .D1(MixerOutSin[11]), 
          .CIN(n11189), .S0(d1_71__N_417[70]), .S1(d1_71__N_417[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_983_37.INIT0 = 16'hd1e2;
    defparam add_983_37.INIT1 = 16'hd1e2;
    defparam add_983_37.INJECT1_0 = "NO";
    defparam add_983_37.INJECT1_1 = "NO";
    CCU2D add_983_35 (.A0(d1[68]), .B0(n4038), .C0(n4077[32]), .D0(MixerOutSin[11]), 
          .A1(d1[69]), .B1(n4038), .C1(n4077[33]), .D1(MixerOutSin[11]), 
          .CIN(n11188), .COUT(n11189), .S0(d1_71__N_417[68]), .S1(d1_71__N_417[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_983_35.INIT0 = 16'hd1e2;
    defparam add_983_35.INIT1 = 16'hd1e2;
    defparam add_983_35.INJECT1_0 = "NO";
    defparam add_983_35.INJECT1_1 = "NO";
    CCU2D add_983_33 (.A0(d1[66]), .B0(n4038), .C0(n4077[30]), .D0(MixerOutSin[11]), 
          .A1(d1[67]), .B1(n4038), .C1(n4077[31]), .D1(MixerOutSin[11]), 
          .CIN(n11187), .COUT(n11188), .S0(d1_71__N_417[66]), .S1(d1_71__N_417[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_983_33.INIT0 = 16'hd1e2;
    defparam add_983_33.INIT1 = 16'hd1e2;
    defparam add_983_33.INJECT1_0 = "NO";
    defparam add_983_33.INJECT1_1 = "NO";
    CCU2D add_983_31 (.A0(d1[64]), .B0(n4038), .C0(n4077[28]), .D0(MixerOutSin[11]), 
          .A1(d1[65]), .B1(n4038), .C1(n4077[29]), .D1(MixerOutSin[11]), 
          .CIN(n11186), .COUT(n11187), .S0(d1_71__N_417[64]), .S1(d1_71__N_417[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_983_31.INIT0 = 16'hd1e2;
    defparam add_983_31.INIT1 = 16'hd1e2;
    defparam add_983_31.INJECT1_0 = "NO";
    defparam add_983_31.INJECT1_1 = "NO";
    CCU2D add_983_29 (.A0(d1[62]), .B0(n4038), .C0(n4077[26]), .D0(MixerOutSin[11]), 
          .A1(d1[63]), .B1(n4038), .C1(n4077[27]), .D1(MixerOutSin[11]), 
          .CIN(n11185), .COUT(n11186), .S0(d1_71__N_417[62]), .S1(d1_71__N_417[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_983_29.INIT0 = 16'hd1e2;
    defparam add_983_29.INIT1 = 16'hd1e2;
    defparam add_983_29.INJECT1_0 = "NO";
    defparam add_983_29.INJECT1_1 = "NO";
    CCU2D add_983_27 (.A0(d1[60]), .B0(n4038), .C0(n4077[24]), .D0(MixerOutSin[11]), 
          .A1(d1[61]), .B1(n4038), .C1(n4077[25]), .D1(MixerOutSin[11]), 
          .CIN(n11184), .COUT(n11185), .S0(d1_71__N_417[60]), .S1(d1_71__N_417[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_983_27.INIT0 = 16'hd1e2;
    defparam add_983_27.INIT1 = 16'hd1e2;
    defparam add_983_27.INJECT1_0 = "NO";
    defparam add_983_27.INJECT1_1 = "NO";
    LUT4 mux_1208_i2_3_lut (.A(n6319[21]), .B(n6357[21]), .C(n6318), .Z(d10_71__N_1746[57])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1208_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1208_i3_3_lut (.A(n6319[22]), .B(n6357[22]), .C(n6318), .Z(d10_71__N_1746[58])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1208_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1208_i4_3_lut (.A(n6319[23]), .B(n6357[23]), .C(n6318), .Z(d10_71__N_1746[59])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1208_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1208_i5_3_lut (.A(n6319[24]), .B(n6357[24]), .C(n6318), .Z(d10_71__N_1746[60])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1208_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1208_i6_3_lut (.A(n6319[25]), .B(n6357[25]), .C(n6318), .Z(d10_71__N_1746[61])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1208_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1208_i7_3_lut (.A(n6319[26]), .B(n6357[26]), .C(n6318), .Z(d10_71__N_1746[62])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1208_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1208_i8_3_lut (.A(n6319[27]), .B(n6357[27]), .C(n6318), .Z(d10_71__N_1746[63])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1208_i8_3_lut.init = 16'hcaca;
    LUT4 i4749_2_lut (.A(d1[0]), .B(d2[0]), .Z(d2_71__N_489[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4749_2_lut.init = 16'h6666;
    LUT4 i5855_4_lut_rep_196 (.A(n13252), .B(n13), .C(n13254), .D(n13238), 
         .Z(osc_clk_enable_62)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i5855_4_lut_rep_196.init = 16'h2000;
    LUT4 mux_1208_i9_3_lut (.A(n6319[28]), .B(n6357[28]), .C(n6318), .Z(d10_71__N_1746[64])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1208_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1208_i10_3_lut (.A(n6319[29]), .B(n6357[29]), .C(n6318), 
         .Z(d10_71__N_1746[65])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1208_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1208_i11_3_lut (.A(n6319[30]), .B(n6357[30]), .C(n6318), 
         .Z(d10_71__N_1746[66])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1208_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1208_i12_3_lut (.A(n6319[31]), .B(n6357[31]), .C(n6318), 
         .Z(d10_71__N_1746[67])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1208_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1208_i13_3_lut (.A(n6319[32]), .B(n6357[32]), .C(n6318), 
         .Z(d10_71__N_1746[68])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1208_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1208_i14_3_lut (.A(n6319[33]), .B(n6357[33]), .C(n6318), 
         .Z(d10_71__N_1746[69])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1208_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1208_i15_3_lut (.A(n6319[34]), .B(n6357[34]), .C(n6318), 
         .Z(d10_71__N_1746[70])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1208_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1208_i16_3_lut (.A(n6319[35]), .B(n6357[35]), .C(n6318), 
         .Z(d10_71__N_1746[71])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1208_i16_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i62_3_lut (.A(d10[61]), .B(d10[62]), .C(\CICGain[0] ), 
         .Z(n62_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i62_3_lut.init = 16'hcaca;
    CCU2D add_1034_37 (.A0(d_d6[70]), .B0(n5558), .C0(n5559[34]), .D0(d6[70]), 
          .A1(d_d6[71]), .B1(n5558), .C1(n5559[35]), .D1(d6[71]), .CIN(n11727), 
          .S0(d7_71__N_1530[70]), .S1(d7_71__N_1530[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1034_37.INIT0 = 16'hb874;
    defparam add_1034_37.INIT1 = 16'hb874;
    defparam add_1034_37.INJECT1_0 = "NO";
    defparam add_1034_37.INJECT1_1 = "NO";
    CCU2D add_998_8 (.A0(d3[42]), .B0(d4[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[43]), .B1(d4[43]), .C1(GND_net), .D1(GND_net), .CIN(n12018), 
          .COUT(n12019), .S0(n4495[6]), .S1(n4495[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_998_8.INIT0 = 16'h5666;
    defparam add_998_8.INIT1 = 16'h5666;
    defparam add_998_8.INJECT1_0 = "NO";
    defparam add_998_8.INJECT1_1 = "NO";
    CCU2D add_998_6 (.A0(d3[40]), .B0(d4[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[41]), .B1(d4[41]), .C1(GND_net), .D1(GND_net), .CIN(n12017), 
          .COUT(n12018), .S0(n4495[4]), .S1(n4495[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_998_6.INIT0 = 16'h5666;
    defparam add_998_6.INIT1 = 16'h5666;
    defparam add_998_6.INJECT1_0 = "NO";
    defparam add_998_6.INJECT1_1 = "NO";
    CCU2D add_998_4 (.A0(d3[38]), .B0(d4[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[39]), .B1(d4[39]), .C1(GND_net), .D1(GND_net), .CIN(n12016), 
          .COUT(n12017), .S0(n4495[2]), .S1(n4495[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_998_4.INIT0 = 16'h5666;
    defparam add_998_4.INIT1 = 16'h5666;
    defparam add_998_4.INJECT1_0 = "NO";
    defparam add_998_4.INJECT1_1 = "NO";
    CCU2D add_998_2 (.A0(d3[36]), .B0(d4[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[37]), .B1(d4[37]), .C1(GND_net), .D1(GND_net), .COUT(n12016), 
          .S1(n4495[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_998_2.INIT0 = 16'h7000;
    defparam add_998_2.INIT1 = 16'h5666;
    defparam add_998_2.INJECT1_0 = "NO";
    defparam add_998_2.INJECT1_1 = "NO";
    LUT4 shift_right_31_i63_3_lut (.A(d10[62]), .B(d10[63]), .C(\CICGain[0] ), 
         .Z(n63_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i63_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i64_3_lut (.A(d10[63]), .B(d10[64]), .C(\CICGain[0] ), 
         .Z(n64_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i64_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i65_3_lut (.A(d10[64]), .B(d10[65]), .C(\CICGain[0] ), 
         .Z(n65_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i65_3_lut.init = 16'hcaca;
    LUT4 i5948_then_3_lut (.A(\CICGain[1] ), .B(d10[59]), .C(d10[57]), 
         .Z(n13799)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i5948_then_3_lut.init = 16'he4e4;
    LUT4 i5948_else_3_lut (.A(n61_c), .B(\CICGain[1] ), .C(d10[58]), .Z(n13798)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i5948_else_3_lut.init = 16'he2e2;
    CCU2D add_999_37 (.A0(d4[70]), .B0(n4494), .C0(n4495[34]), .D0(d3[70]), 
          .A1(d4[71]), .B1(n4494), .C1(n4495[35]), .D1(d3[71]), .CIN(n12013), 
          .S0(d4_71__N_633[70]), .S1(d4_71__N_633[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_999_37.INIT0 = 16'h74b8;
    defparam add_999_37.INIT1 = 16'h74b8;
    defparam add_999_37.INJECT1_0 = "NO";
    defparam add_999_37.INJECT1_1 = "NO";
    LUT4 shift_right_31_i66_3_lut (.A(d10[65]), .B(d10[66]), .C(\CICGain[0] ), 
         .Z(n66_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i66_3_lut.init = 16'hcaca;
    LUT4 i4816_2_lut (.A(MixerOutSin[11]), .B(d1[36]), .Z(n12116)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i4816_2_lut.init = 16'h9999;
    CCU2D add_999_35 (.A0(d4[68]), .B0(n4494), .C0(n4495[32]), .D0(d3[68]), 
          .A1(d4[69]), .B1(n4494), .C1(n4495[33]), .D1(d3[69]), .CIN(n12012), 
          .COUT(n12013), .S0(d4_71__N_633[68]), .S1(d4_71__N_633[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_999_35.INIT0 = 16'h74b8;
    defparam add_999_35.INIT1 = 16'h74b8;
    defparam add_999_35.INJECT1_0 = "NO";
    defparam add_999_35.INJECT1_1 = "NO";
    CCU2D add_999_33 (.A0(d4[66]), .B0(n4494), .C0(n4495[30]), .D0(d3[66]), 
          .A1(d4[67]), .B1(n4494), .C1(n4495[31]), .D1(d3[67]), .CIN(n12011), 
          .COUT(n12012), .S0(d4_71__N_633[66]), .S1(d4_71__N_633[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_999_33.INIT0 = 16'h74b8;
    defparam add_999_33.INIT1 = 16'h74b8;
    defparam add_999_33.INJECT1_0 = "NO";
    defparam add_999_33.INJECT1_1 = "NO";
    CCU2D add_999_31 (.A0(d4[64]), .B0(n4494), .C0(n4495[28]), .D0(d3[64]), 
          .A1(d4[65]), .B1(n4494), .C1(n4495[29]), .D1(d3[65]), .CIN(n12010), 
          .COUT(n12011), .S0(d4_71__N_633[64]), .S1(d4_71__N_633[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_999_31.INIT0 = 16'h74b8;
    defparam add_999_31.INIT1 = 16'h74b8;
    defparam add_999_31.INJECT1_0 = "NO";
    defparam add_999_31.INJECT1_1 = "NO";
    CCU2D add_999_29 (.A0(d4[62]), .B0(n4494), .C0(n4495[26]), .D0(d3[62]), 
          .A1(d4[63]), .B1(n4494), .C1(n4495[27]), .D1(d3[63]), .CIN(n12009), 
          .COUT(n12010), .S0(d4_71__N_633[62]), .S1(d4_71__N_633[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_999_29.INIT0 = 16'h74b8;
    defparam add_999_29.INIT1 = 16'h74b8;
    defparam add_999_29.INJECT1_0 = "NO";
    defparam add_999_29.INJECT1_1 = "NO";
    LUT4 shift_right_31_i67_3_lut (.A(d10[66]), .B(d10[67]), .C(\CICGain[0] ), 
         .Z(n67_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i67_3_lut.init = 16'hcaca;
    CCU2D add_999_27 (.A0(d4[60]), .B0(n4494), .C0(n4495[24]), .D0(d3[60]), 
          .A1(d4[61]), .B1(n4494), .C1(n4495[25]), .D1(d3[61]), .CIN(n12008), 
          .COUT(n12009), .S0(d4_71__N_633[60]), .S1(d4_71__N_633[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_999_27.INIT0 = 16'h74b8;
    defparam add_999_27.INIT1 = 16'h74b8;
    defparam add_999_27.INJECT1_0 = "NO";
    defparam add_999_27.INJECT1_1 = "NO";
    LUT4 shift_right_31_i68_3_lut (.A(d10[67]), .B(d10[68]), .C(\CICGain[0] ), 
         .Z(n68_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i68_3_lut.init = 16'hcaca;
    CCU2D add_999_25 (.A0(d4[58]), .B0(n4494), .C0(n4495[22]), .D0(d3[58]), 
          .A1(d4[59]), .B1(n4494), .C1(n4495[23]), .D1(d3[59]), .CIN(n12007), 
          .COUT(n12008), .S0(d4_71__N_633[58]), .S1(d4_71__N_633[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_999_25.INIT0 = 16'h74b8;
    defparam add_999_25.INIT1 = 16'h74b8;
    defparam add_999_25.INJECT1_0 = "NO";
    defparam add_999_25.INJECT1_1 = "NO";
    CCU2D add_999_23 (.A0(d4[56]), .B0(n4494), .C0(n4495[20]), .D0(d3[56]), 
          .A1(d4[57]), .B1(n4494), .C1(n4495[21]), .D1(d3[57]), .CIN(n12006), 
          .COUT(n12007), .S0(d4_71__N_633[56]), .S1(d4_71__N_633[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_999_23.INIT0 = 16'h74b8;
    defparam add_999_23.INIT1 = 16'h74b8;
    defparam add_999_23.INJECT1_0 = "NO";
    defparam add_999_23.INJECT1_1 = "NO";
    CCU2D add_999_21 (.A0(d4[54]), .B0(n4494), .C0(n4495[18]), .D0(d3[54]), 
          .A1(d4[55]), .B1(n4494), .C1(n4495[19]), .D1(d3[55]), .CIN(n12005), 
          .COUT(n12006), .S0(d4_71__N_633[54]), .S1(d4_71__N_633[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_999_21.INIT0 = 16'h74b8;
    defparam add_999_21.INIT1 = 16'h74b8;
    defparam add_999_21.INJECT1_0 = "NO";
    defparam add_999_21.INJECT1_1 = "NO";
    CCU2D add_999_19 (.A0(d4[52]), .B0(n4494), .C0(n4495[16]), .D0(d3[52]), 
          .A1(d4[53]), .B1(n4494), .C1(n4495[17]), .D1(d3[53]), .CIN(n12004), 
          .COUT(n12005), .S0(d4_71__N_633[52]), .S1(d4_71__N_633[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_999_19.INIT0 = 16'h74b8;
    defparam add_999_19.INIT1 = 16'h74b8;
    defparam add_999_19.INJECT1_0 = "NO";
    defparam add_999_19.INJECT1_1 = "NO";
    FD1S3AX v_comb_66_rep_194 (.D(osc_clk_enable_62), .CK(osc_clk), .Q(osc_clk_enable_696)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_194.GSR = "ENABLED";
    CCU2D add_1039_23 (.A0(d_d7[56]), .B0(n5710), .C0(n5711[20]), .D0(d7[56]), 
          .A1(d_d7[57]), .B1(n5710), .C1(n5711[21]), .D1(d7[57]), .CIN(n11680), 
          .COUT(n11681), .S0(d8_71__N_1602[56]), .S1(d8_71__N_1602[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1039_23.INIT0 = 16'hb874;
    defparam add_1039_23.INIT1 = 16'hb874;
    defparam add_1039_23.INJECT1_0 = "NO";
    defparam add_1039_23.INJECT1_1 = "NO";
    CCU2D add_1039_21 (.A0(d_d7[54]), .B0(n5710), .C0(n5711[18]), .D0(d7[54]), 
          .A1(d_d7[55]), .B1(n5710), .C1(n5711[19]), .D1(d7[55]), .CIN(n11679), 
          .COUT(n11680), .S0(d8_71__N_1602[54]), .S1(d8_71__N_1602[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1039_21.INIT0 = 16'hb874;
    defparam add_1039_21.INIT1 = 16'hb874;
    defparam add_1039_21.INJECT1_0 = "NO";
    defparam add_1039_21.INJECT1_1 = "NO";
    CCU2D add_1039_19 (.A0(d_d7[52]), .B0(n5710), .C0(n5711[16]), .D0(d7[52]), 
          .A1(d_d7[53]), .B1(n5710), .C1(n5711[17]), .D1(d7[53]), .CIN(n11678), 
          .COUT(n11679), .S0(d8_71__N_1602[52]), .S1(d8_71__N_1602[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1039_19.INIT0 = 16'hb874;
    defparam add_1039_19.INIT1 = 16'hb874;
    defparam add_1039_19.INJECT1_0 = "NO";
    defparam add_1039_19.INJECT1_1 = "NO";
    CCU2D add_1039_17 (.A0(d_d7[50]), .B0(n5710), .C0(n5711[14]), .D0(d7[50]), 
          .A1(d_d7[51]), .B1(n5710), .C1(n5711[15]), .D1(d7[51]), .CIN(n11677), 
          .COUT(n11678), .S0(d8_71__N_1602[50]), .S1(d8_71__N_1602[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1039_17.INIT0 = 16'hb874;
    defparam add_1039_17.INIT1 = 16'hb874;
    defparam add_1039_17.INJECT1_0 = "NO";
    defparam add_1039_17.INJECT1_1 = "NO";
    CCU2D add_1039_15 (.A0(d_d7[48]), .B0(n5710), .C0(n5711[12]), .D0(d7[48]), 
          .A1(d_d7[49]), .B1(n5710), .C1(n5711[13]), .D1(d7[49]), .CIN(n11676), 
          .COUT(n11677), .S0(d8_71__N_1602[48]), .S1(d8_71__N_1602[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1039_15.INIT0 = 16'hb874;
    defparam add_1039_15.INIT1 = 16'hb874;
    defparam add_1039_15.INJECT1_0 = "NO";
    defparam add_1039_15.INJECT1_1 = "NO";
    CCU2D add_1039_13 (.A0(d_d7[46]), .B0(n5710), .C0(n5711[10]), .D0(d7[46]), 
          .A1(d_d7[47]), .B1(n5710), .C1(n5711[11]), .D1(d7[47]), .CIN(n11675), 
          .COUT(n11676), .S0(d8_71__N_1602[46]), .S1(d8_71__N_1602[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1039_13.INIT0 = 16'hb874;
    defparam add_1039_13.INIT1 = 16'hb874;
    defparam add_1039_13.INJECT1_0 = "NO";
    defparam add_1039_13.INJECT1_1 = "NO";
    CCU2D add_1039_11 (.A0(d_d7[44]), .B0(n5710), .C0(n5711[8]), .D0(d7[44]), 
          .A1(d_d7[45]), .B1(n5710), .C1(n5711[9]), .D1(d7[45]), .CIN(n11674), 
          .COUT(n11675), .S0(d8_71__N_1602[44]), .S1(d8_71__N_1602[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1039_11.INIT0 = 16'hb874;
    defparam add_1039_11.INIT1 = 16'hb874;
    defparam add_1039_11.INJECT1_0 = "NO";
    defparam add_1039_11.INJECT1_1 = "NO";
    CCU2D add_1039_9 (.A0(d_d7[42]), .B0(n5710), .C0(n5711[6]), .D0(d7[42]), 
          .A1(d_d7[43]), .B1(n5710), .C1(n5711[7]), .D1(d7[43]), .CIN(n11673), 
          .COUT(n11674), .S0(d8_71__N_1602[42]), .S1(d8_71__N_1602[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1039_9.INIT0 = 16'hb874;
    defparam add_1039_9.INIT1 = 16'hb874;
    defparam add_1039_9.INJECT1_0 = "NO";
    defparam add_1039_9.INJECT1_1 = "NO";
    CCU2D add_1039_7 (.A0(d_d7[40]), .B0(n5710), .C0(n5711[4]), .D0(d7[40]), 
          .A1(d_d7[41]), .B1(n5710), .C1(n5711[5]), .D1(d7[41]), .CIN(n11672), 
          .COUT(n11673), .S0(d8_71__N_1602[40]), .S1(d8_71__N_1602[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1039_7.INIT0 = 16'hb874;
    defparam add_1039_7.INIT1 = 16'hb874;
    defparam add_1039_7.INJECT1_0 = "NO";
    defparam add_1039_7.INJECT1_1 = "NO";
    CCU2D add_1039_5 (.A0(d_d7[38]), .B0(n5710), .C0(n5711[2]), .D0(d7[38]), 
          .A1(d_d7[39]), .B1(n5710), .C1(n5711[3]), .D1(d7[39]), .CIN(n11671), 
          .COUT(n11672), .S0(d8_71__N_1602[38]), .S1(d8_71__N_1602[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1039_5.INIT0 = 16'hb874;
    defparam add_1039_5.INIT1 = 16'hb874;
    defparam add_1039_5.INJECT1_0 = "NO";
    defparam add_1039_5.INJECT1_1 = "NO";
    CCU2D add_1039_3 (.A0(d_d7[36]), .B0(n5710), .C0(n5711[0]), .D0(d7[36]), 
          .A1(d_d7[37]), .B1(n5710), .C1(n5711[1]), .D1(d7[37]), .CIN(n11670), 
          .COUT(n11671), .S0(d8_71__N_1602[36]), .S1(d8_71__N_1602[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1039_3.INIT0 = 16'hb874;
    defparam add_1039_3.INIT1 = 16'hb874;
    defparam add_1039_3.INJECT1_0 = "NO";
    defparam add_1039_3.INJECT1_1 = "NO";
    CCU2D add_1039_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5710), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11670));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1039_1.INIT0 = 16'hF000;
    defparam add_1039_1.INIT1 = 16'h0555;
    defparam add_1039_1.INJECT1_0 = "NO";
    defparam add_1039_1.INJECT1_1 = "NO";
    LUT4 shift_right_31_i70_3_lut (.A(d10[69]), .B(d10[70]), .C(\CICGain[0] ), 
         .Z(n70_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i70_3_lut.init = 16'hcaca;
    LUT4 i11_3_lut_4_lut_then_3_lut_adj_35 (.A(\CICGain[0] ), .B(\d10[67] ), 
         .C(\d10[68] ), .Z(n13808)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam i11_3_lut_4_lut_then_3_lut_adj_35.init = 16'hd8d8;
    LUT4 i11_3_lut_4_lut_else_3_lut_adj_36 (.A(\CICGain[0] ), .B(\d10[69] ), 
         .C(\d10[70] ), .Z(n13807)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam i11_3_lut_4_lut_else_3_lut_adj_36.init = 16'hd8d8;
    LUT4 i4812_2_lut (.A(d2[36]), .B(d3[36]), .Z(n4343[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4812_2_lut.init = 16'h6666;
    FD1S3AX v_comb_66_rep_193 (.D(osc_clk_enable_62), .CK(osc_clk), .Q(osc_clk_enable_646)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_193.GSR = "ENABLED";
    CCU2D add_983_25 (.A0(d1[58]), .B0(n4038), .C0(n4077[22]), .D0(MixerOutSin[11]), 
          .A1(d1[59]), .B1(n4038), .C1(n4077[23]), .D1(MixerOutSin[11]), 
          .CIN(n11183), .COUT(n11184), .S0(d1_71__N_417[58]), .S1(d1_71__N_417[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_983_25.INIT0 = 16'hd1e2;
    defparam add_983_25.INIT1 = 16'hd1e2;
    defparam add_983_25.INJECT1_0 = "NO";
    defparam add_983_25.INJECT1_1 = "NO";
    CCU2D add_983_23 (.A0(d1[56]), .B0(n4038), .C0(n4077[20]), .D0(MixerOutSin[11]), 
          .A1(d1[57]), .B1(n4038), .C1(n4077[21]), .D1(MixerOutSin[11]), 
          .CIN(n11182), .COUT(n11183), .S0(d1_71__N_417[56]), .S1(d1_71__N_417[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_983_23.INIT0 = 16'hd1e2;
    defparam add_983_23.INIT1 = 16'hd1e2;
    defparam add_983_23.INJECT1_0 = "NO";
    defparam add_983_23.INJECT1_1 = "NO";
    CCU2D add_983_21 (.A0(d1[54]), .B0(n4038), .C0(n4077[18]), .D0(MixerOutSin[11]), 
          .A1(d1[55]), .B1(n4038), .C1(n4077[19]), .D1(MixerOutSin[11]), 
          .CIN(n11181), .COUT(n11182), .S0(d1_71__N_417[54]), .S1(d1_71__N_417[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_983_21.INIT0 = 16'hd1e2;
    defparam add_983_21.INIT1 = 16'hd1e2;
    defparam add_983_21.INJECT1_0 = "NO";
    defparam add_983_21.INJECT1_1 = "NO";
    CCU2D add_983_19 (.A0(d1[52]), .B0(n4038), .C0(n4077[16]), .D0(MixerOutSin[11]), 
          .A1(d1[53]), .B1(n4038), .C1(n4077[17]), .D1(MixerOutSin[11]), 
          .CIN(n11180), .COUT(n11181), .S0(d1_71__N_417[52]), .S1(d1_71__N_417[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_983_19.INIT0 = 16'hd1e2;
    defparam add_983_19.INIT1 = 16'hd1e2;
    defparam add_983_19.INJECT1_0 = "NO";
    defparam add_983_19.INJECT1_1 = "NO";
    CCU2D add_983_17 (.A0(d1[50]), .B0(n4038), .C0(n4077[14]), .D0(MixerOutSin[11]), 
          .A1(d1[51]), .B1(n4038), .C1(n4077[15]), .D1(MixerOutSin[11]), 
          .CIN(n11179), .COUT(n11180), .S0(d1_71__N_417[50]), .S1(d1_71__N_417[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_983_17.INIT0 = 16'hd1e2;
    defparam add_983_17.INIT1 = 16'hd1e2;
    defparam add_983_17.INJECT1_0 = "NO";
    defparam add_983_17.INJECT1_1 = "NO";
    CCU2D add_983_15 (.A0(d1[48]), .B0(n4038), .C0(n4077[12]), .D0(MixerOutSin[11]), 
          .A1(d1[49]), .B1(n4038), .C1(n4077[13]), .D1(MixerOutSin[11]), 
          .CIN(n11178), .COUT(n11179), .S0(d1_71__N_417[48]), .S1(d1_71__N_417[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_983_15.INIT0 = 16'hd1e2;
    defparam add_983_15.INIT1 = 16'hd1e2;
    defparam add_983_15.INJECT1_0 = "NO";
    defparam add_983_15.INJECT1_1 = "NO";
    CCU2D add_983_13 (.A0(d1[46]), .B0(n4038), .C0(n4077[10]), .D0(MixerOutSin[11]), 
          .A1(d1[47]), .B1(n4038), .C1(n4077[11]), .D1(MixerOutSin[11]), 
          .CIN(n11177), .COUT(n11178), .S0(d1_71__N_417[46]), .S1(d1_71__N_417[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_983_13.INIT0 = 16'hd1e2;
    defparam add_983_13.INIT1 = 16'hd1e2;
    defparam add_983_13.INJECT1_0 = "NO";
    defparam add_983_13.INJECT1_1 = "NO";
    CCU2D add_983_11 (.A0(d1[44]), .B0(n4038), .C0(n4077[8]), .D0(MixerOutSin[11]), 
          .A1(d1[45]), .B1(n4038), .C1(n4077[9]), .D1(MixerOutSin[11]), 
          .CIN(n11176), .COUT(n11177), .S0(d1_71__N_417[44]), .S1(d1_71__N_417[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_983_11.INIT0 = 16'hd1e2;
    defparam add_983_11.INIT1 = 16'hd1e2;
    defparam add_983_11.INJECT1_0 = "NO";
    defparam add_983_11.INJECT1_1 = "NO";
    CCU2D add_983_9 (.A0(d1[42]), .B0(n4038), .C0(n4077[6]), .D0(MixerOutSin[11]), 
          .A1(d1[43]), .B1(n4038), .C1(n4077[7]), .D1(MixerOutSin[11]), 
          .CIN(n11175), .COUT(n11176), .S0(d1_71__N_417[42]), .S1(d1_71__N_417[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_983_9.INIT0 = 16'hd1e2;
    defparam add_983_9.INIT1 = 16'hd1e2;
    defparam add_983_9.INJECT1_0 = "NO";
    defparam add_983_9.INJECT1_1 = "NO";
    CCU2D add_983_7 (.A0(d1[40]), .B0(n4038), .C0(n4077[4]), .D0(MixerOutSin[11]), 
          .A1(d1[41]), .B1(n4038), .C1(n4077[5]), .D1(MixerOutSin[11]), 
          .CIN(n11174), .COUT(n11175), .S0(d1_71__N_417[40]), .S1(d1_71__N_417[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_983_7.INIT0 = 16'hd1e2;
    defparam add_983_7.INIT1 = 16'hd1e2;
    defparam add_983_7.INJECT1_0 = "NO";
    defparam add_983_7.INJECT1_1 = "NO";
    CCU2D add_983_5 (.A0(d1[38]), .B0(n4038), .C0(n4077[2]), .D0(MixerOutSin[11]), 
          .A1(d1[39]), .B1(n4038), .C1(n4077[3]), .D1(MixerOutSin[11]), 
          .CIN(n11173), .COUT(n11174), .S0(d1_71__N_417[38]), .S1(d1_71__N_417[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_983_5.INIT0 = 16'hd1e2;
    defparam add_983_5.INIT1 = 16'hd1e2;
    defparam add_983_5.INJECT1_0 = "NO";
    defparam add_983_5.INJECT1_1 = "NO";
    CCU2D add_983_3 (.A0(d1[36]), .B0(n4038), .C0(n12116), .D0(MixerOutSin[11]), 
          .A1(d1[37]), .B1(n4038), .C1(n4077[1]), .D1(MixerOutSin[11]), 
          .CIN(n11172), .COUT(n11173), .S0(d1_71__N_417[36]), .S1(d1_71__N_417[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_983_3.INIT0 = 16'hd1e2;
    defparam add_983_3.INIT1 = 16'hd1e2;
    defparam add_983_3.INJECT1_0 = "NO";
    defparam add_983_3.INJECT1_1 = "NO";
    CCU2D add_983_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n4038), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11172));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_983_1.INIT0 = 16'hF000;
    defparam add_983_1.INIT1 = 16'h0fff;
    defparam add_983_1.INJECT1_0 = "NO";
    defparam add_983_1.INJECT1_1 = "NO";
    CCU2D add_1077_37 (.A0(d_tmp[35]), .B0(d_d_tmp[35]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11168), .S0(d6_71__N_1458[35]), .S1(n6926));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1077_37.INIT0 = 16'h5999;
    defparam add_1077_37.INIT1 = 16'h0000;
    defparam add_1077_37.INJECT1_0 = "NO";
    defparam add_1077_37.INJECT1_1 = "NO";
    CCU2D add_1077_35 (.A0(d_tmp[33]), .B0(d_d_tmp[33]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[34]), .B1(d_d_tmp[34]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11167), .COUT(n11168), .S0(d6_71__N_1458[33]), 
          .S1(d6_71__N_1458[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1077_35.INIT0 = 16'h5999;
    defparam add_1077_35.INIT1 = 16'h5999;
    defparam add_1077_35.INJECT1_0 = "NO";
    defparam add_1077_35.INJECT1_1 = "NO";
    CCU2D add_1077_33 (.A0(d_tmp[31]), .B0(d_d_tmp[31]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[32]), .B1(d_d_tmp[32]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11166), .COUT(n11167), .S0(d6_71__N_1458[31]), 
          .S1(d6_71__N_1458[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1077_33.INIT0 = 16'h5999;
    defparam add_1077_33.INIT1 = 16'h5999;
    defparam add_1077_33.INJECT1_0 = "NO";
    defparam add_1077_33.INJECT1_1 = "NO";
    CCU2D add_1077_31 (.A0(d_tmp[29]), .B0(d_d_tmp[29]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[30]), .B1(d_d_tmp[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11165), .COUT(n11166), .S0(d6_71__N_1458[29]), 
          .S1(d6_71__N_1458[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1077_31.INIT0 = 16'h5999;
    defparam add_1077_31.INIT1 = 16'h5999;
    defparam add_1077_31.INJECT1_0 = "NO";
    defparam add_1077_31.INJECT1_1 = "NO";
    CCU2D add_1077_29 (.A0(d_tmp[27]), .B0(d_d_tmp[27]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[28]), .B1(d_d_tmp[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11164), .COUT(n11165), .S0(d6_71__N_1458[27]), 
          .S1(d6_71__N_1458[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1077_29.INIT0 = 16'h5999;
    defparam add_1077_29.INIT1 = 16'h5999;
    defparam add_1077_29.INJECT1_0 = "NO";
    defparam add_1077_29.INJECT1_1 = "NO";
    CCU2D add_1077_27 (.A0(d_tmp[25]), .B0(d_d_tmp[25]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[26]), .B1(d_d_tmp[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11163), .COUT(n11164), .S0(d6_71__N_1458[25]), 
          .S1(d6_71__N_1458[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1077_27.INIT0 = 16'h5999;
    defparam add_1077_27.INIT1 = 16'h5999;
    defparam add_1077_27.INJECT1_0 = "NO";
    defparam add_1077_27.INJECT1_1 = "NO";
    CCU2D add_1077_25 (.A0(d_tmp[23]), .B0(d_d_tmp[23]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[24]), .B1(d_d_tmp[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11162), .COUT(n11163), .S0(d6_71__N_1458[23]), 
          .S1(d6_71__N_1458[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1077_25.INIT0 = 16'h5999;
    defparam add_1077_25.INIT1 = 16'h5999;
    defparam add_1077_25.INJECT1_0 = "NO";
    defparam add_1077_25.INJECT1_1 = "NO";
    CCU2D add_1077_23 (.A0(d_tmp[21]), .B0(d_d_tmp[21]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[22]), .B1(d_d_tmp[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11161), .COUT(n11162), .S0(d6_71__N_1458[21]), 
          .S1(d6_71__N_1458[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1077_23.INIT0 = 16'h5999;
    defparam add_1077_23.INIT1 = 16'h5999;
    defparam add_1077_23.INJECT1_0 = "NO";
    defparam add_1077_23.INJECT1_1 = "NO";
    CCU2D add_1077_21 (.A0(d_tmp[19]), .B0(d_d_tmp[19]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[20]), .B1(d_d_tmp[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11160), .COUT(n11161), .S0(d6_71__N_1458[19]), 
          .S1(d6_71__N_1458[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1077_21.INIT0 = 16'h5999;
    defparam add_1077_21.INIT1 = 16'h5999;
    defparam add_1077_21.INJECT1_0 = "NO";
    defparam add_1077_21.INJECT1_1 = "NO";
    CCU2D add_1077_19 (.A0(d_tmp[17]), .B0(d_d_tmp[17]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[18]), .B1(d_d_tmp[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11159), .COUT(n11160), .S0(d6_71__N_1458[17]), 
          .S1(d6_71__N_1458[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1077_19.INIT0 = 16'h5999;
    defparam add_1077_19.INIT1 = 16'h5999;
    defparam add_1077_19.INJECT1_0 = "NO";
    defparam add_1077_19.INJECT1_1 = "NO";
    CCU2D add_1077_17 (.A0(d_tmp[15]), .B0(d_d_tmp[15]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[16]), .B1(d_d_tmp[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11158), .COUT(n11159), .S0(d6_71__N_1458[15]), 
          .S1(d6_71__N_1458[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1077_17.INIT0 = 16'h5999;
    defparam add_1077_17.INIT1 = 16'h5999;
    defparam add_1077_17.INJECT1_0 = "NO";
    defparam add_1077_17.INJECT1_1 = "NO";
    CCU2D add_1077_15 (.A0(d_tmp[13]), .B0(d_d_tmp[13]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[14]), .B1(d_d_tmp[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11157), .COUT(n11158), .S0(d6_71__N_1458[13]), 
          .S1(d6_71__N_1458[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1077_15.INIT0 = 16'h5999;
    defparam add_1077_15.INIT1 = 16'h5999;
    defparam add_1077_15.INJECT1_0 = "NO";
    defparam add_1077_15.INJECT1_1 = "NO";
    CCU2D add_1077_13 (.A0(d_tmp[11]), .B0(d_d_tmp[11]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[12]), .B1(d_d_tmp[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11156), .COUT(n11157), .S0(d6_71__N_1458[11]), 
          .S1(d6_71__N_1458[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1077_13.INIT0 = 16'h5999;
    defparam add_1077_13.INIT1 = 16'h5999;
    defparam add_1077_13.INJECT1_0 = "NO";
    defparam add_1077_13.INJECT1_1 = "NO";
    CCU2D add_1077_11 (.A0(d_tmp[9]), .B0(d_d_tmp[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[10]), .B1(d_d_tmp[10]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11155), .COUT(n11156), .S0(d6_71__N_1458[9]), .S1(d6_71__N_1458[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1077_11.INIT0 = 16'h5999;
    defparam add_1077_11.INIT1 = 16'h5999;
    defparam add_1077_11.INJECT1_0 = "NO";
    defparam add_1077_11.INJECT1_1 = "NO";
    CCU2D add_1077_9 (.A0(d_tmp[7]), .B0(d_d_tmp[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[8]), .B1(d_d_tmp[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11154), .COUT(n11155), .S0(d6_71__N_1458[7]), .S1(d6_71__N_1458[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1077_9.INIT0 = 16'h5999;
    defparam add_1077_9.INIT1 = 16'h5999;
    defparam add_1077_9.INJECT1_0 = "NO";
    defparam add_1077_9.INJECT1_1 = "NO";
    CCU2D add_1077_7 (.A0(d_tmp[5]), .B0(d_d_tmp[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[6]), .B1(d_d_tmp[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11153), .COUT(n11154), .S0(d6_71__N_1458[5]), .S1(d6_71__N_1458[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1077_7.INIT0 = 16'h5999;
    defparam add_1077_7.INIT1 = 16'h5999;
    defparam add_1077_7.INJECT1_0 = "NO";
    defparam add_1077_7.INJECT1_1 = "NO";
    CCU2D add_1077_5 (.A0(d_tmp[3]), .B0(d_d_tmp[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[4]), .B1(d_d_tmp[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11152), .COUT(n11153), .S0(d6_71__N_1458[3]), .S1(d6_71__N_1458[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1077_5.INIT0 = 16'h5999;
    defparam add_1077_5.INIT1 = 16'h5999;
    defparam add_1077_5.INJECT1_0 = "NO";
    defparam add_1077_5.INJECT1_1 = "NO";
    CCU2D add_1077_3 (.A0(d_tmp[1]), .B0(d_d_tmp[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[2]), .B1(d_d_tmp[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11151), .COUT(n11152), .S0(d6_71__N_1458[1]), .S1(d6_71__N_1458[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1077_3.INIT0 = 16'h5999;
    defparam add_1077_3.INIT1 = 16'h5999;
    defparam add_1077_3.INJECT1_0 = "NO";
    defparam add_1077_3.INJECT1_1 = "NO";
    CCU2D add_1077_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[0]), .B1(d_d_tmp[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n11151), .S1(d6_71__N_1458[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1077_1.INIT0 = 16'h0000;
    defparam add_1077_1.INIT1 = 16'h5999;
    defparam add_1077_1.INJECT1_0 = "NO";
    defparam add_1077_1.INJECT1_1 = "NO";
    CCU2D add_1062_37 (.A0(d8[35]), .B0(d_d8[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11109), 
          .S0(d9_71__N_1674[35]), .S1(n6470));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1062_37.INIT0 = 16'h5999;
    defparam add_1062_37.INIT1 = 16'h0000;
    defparam add_1062_37.INJECT1_0 = "NO";
    defparam add_1062_37.INJECT1_1 = "NO";
    CCU2D add_1062_35 (.A0(d8[33]), .B0(d_d8[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[34]), .B1(d_d8[34]), .C1(GND_net), .D1(GND_net), .CIN(n11108), 
          .COUT(n11109), .S0(d9_71__N_1674[33]), .S1(d9_71__N_1674[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1062_35.INIT0 = 16'h5999;
    defparam add_1062_35.INIT1 = 16'h5999;
    defparam add_1062_35.INJECT1_0 = "NO";
    defparam add_1062_35.INJECT1_1 = "NO";
    CCU2D add_1062_33 (.A0(d8[31]), .B0(d_d8[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[32]), .B1(d_d8[32]), .C1(GND_net), .D1(GND_net), .CIN(n11107), 
          .COUT(n11108), .S0(d9_71__N_1674[31]), .S1(d9_71__N_1674[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1062_33.INIT0 = 16'h5999;
    defparam add_1062_33.INIT1 = 16'h5999;
    defparam add_1062_33.INJECT1_0 = "NO";
    defparam add_1062_33.INJECT1_1 = "NO";
    CCU2D add_1062_31 (.A0(d8[29]), .B0(d_d8[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[30]), .B1(d_d8[30]), .C1(GND_net), .D1(GND_net), .CIN(n11106), 
          .COUT(n11107), .S0(d9_71__N_1674[29]), .S1(d9_71__N_1674[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1062_31.INIT0 = 16'h5999;
    defparam add_1062_31.INIT1 = 16'h5999;
    defparam add_1062_31.INJECT1_0 = "NO";
    defparam add_1062_31.INJECT1_1 = "NO";
    CCU2D add_1062_29 (.A0(d8[27]), .B0(d_d8[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[28]), .B1(d_d8[28]), .C1(GND_net), .D1(GND_net), .CIN(n11105), 
          .COUT(n11106), .S0(d9_71__N_1674[27]), .S1(d9_71__N_1674[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1062_29.INIT0 = 16'h5999;
    defparam add_1062_29.INIT1 = 16'h5999;
    defparam add_1062_29.INJECT1_0 = "NO";
    defparam add_1062_29.INJECT1_1 = "NO";
    CCU2D add_1062_27 (.A0(d8[25]), .B0(d_d8[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[26]), .B1(d_d8[26]), .C1(GND_net), .D1(GND_net), .CIN(n11104), 
          .COUT(n11105), .S0(d9_71__N_1674[25]), .S1(d9_71__N_1674[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1062_27.INIT0 = 16'h5999;
    defparam add_1062_27.INIT1 = 16'h5999;
    defparam add_1062_27.INJECT1_0 = "NO";
    defparam add_1062_27.INJECT1_1 = "NO";
    CCU2D add_1062_25 (.A0(d8[23]), .B0(d_d8[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[24]), .B1(d_d8[24]), .C1(GND_net), .D1(GND_net), .CIN(n11103), 
          .COUT(n11104), .S0(d9_71__N_1674[23]), .S1(d9_71__N_1674[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1062_25.INIT0 = 16'h5999;
    defparam add_1062_25.INIT1 = 16'h5999;
    defparam add_1062_25.INJECT1_0 = "NO";
    defparam add_1062_25.INJECT1_1 = "NO";
    CCU2D add_1062_23 (.A0(d8[21]), .B0(d_d8[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[22]), .B1(d_d8[22]), .C1(GND_net), .D1(GND_net), .CIN(n11102), 
          .COUT(n11103), .S0(d9_71__N_1674[21]), .S1(d9_71__N_1674[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1062_23.INIT0 = 16'h5999;
    defparam add_1062_23.INIT1 = 16'h5999;
    defparam add_1062_23.INJECT1_0 = "NO";
    defparam add_1062_23.INJECT1_1 = "NO";
    CCU2D add_1062_21 (.A0(d8[19]), .B0(d_d8[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[20]), .B1(d_d8[20]), .C1(GND_net), .D1(GND_net), .CIN(n11101), 
          .COUT(n11102), .S0(d9_71__N_1674[19]), .S1(d9_71__N_1674[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1062_21.INIT0 = 16'h5999;
    defparam add_1062_21.INIT1 = 16'h5999;
    defparam add_1062_21.INJECT1_0 = "NO";
    defparam add_1062_21.INJECT1_1 = "NO";
    CCU2D add_1062_19 (.A0(d8[17]), .B0(d_d8[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[18]), .B1(d_d8[18]), .C1(GND_net), .D1(GND_net), .CIN(n11100), 
          .COUT(n11101), .S0(d9_71__N_1674[17]), .S1(d9_71__N_1674[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1062_19.INIT0 = 16'h5999;
    defparam add_1062_19.INIT1 = 16'h5999;
    defparam add_1062_19.INJECT1_0 = "NO";
    defparam add_1062_19.INJECT1_1 = "NO";
    CCU2D add_1062_17 (.A0(d8[15]), .B0(d_d8[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[16]), .B1(d_d8[16]), .C1(GND_net), .D1(GND_net), .CIN(n11099), 
          .COUT(n11100), .S0(d9_71__N_1674[15]), .S1(d9_71__N_1674[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1062_17.INIT0 = 16'h5999;
    defparam add_1062_17.INIT1 = 16'h5999;
    defparam add_1062_17.INJECT1_0 = "NO";
    defparam add_1062_17.INJECT1_1 = "NO";
    CCU2D add_1062_15 (.A0(d8[13]), .B0(d_d8[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[14]), .B1(d_d8[14]), .C1(GND_net), .D1(GND_net), .CIN(n11098), 
          .COUT(n11099), .S0(d9_71__N_1674[13]), .S1(d9_71__N_1674[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1062_15.INIT0 = 16'h5999;
    defparam add_1062_15.INIT1 = 16'h5999;
    defparam add_1062_15.INJECT1_0 = "NO";
    defparam add_1062_15.INJECT1_1 = "NO";
    CCU2D add_1062_13 (.A0(d8[11]), .B0(d_d8[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[12]), .B1(d_d8[12]), .C1(GND_net), .D1(GND_net), .CIN(n11097), 
          .COUT(n11098), .S0(d9_71__N_1674[11]), .S1(d9_71__N_1674[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1062_13.INIT0 = 16'h5999;
    defparam add_1062_13.INIT1 = 16'h5999;
    defparam add_1062_13.INJECT1_0 = "NO";
    defparam add_1062_13.INJECT1_1 = "NO";
    CCU2D add_1062_11 (.A0(d8[9]), .B0(d_d8[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[10]), .B1(d_d8[10]), .C1(GND_net), .D1(GND_net), .CIN(n11096), 
          .COUT(n11097), .S0(d9_71__N_1674[9]), .S1(d9_71__N_1674[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1062_11.INIT0 = 16'h5999;
    defparam add_1062_11.INIT1 = 16'h5999;
    defparam add_1062_11.INJECT1_0 = "NO";
    defparam add_1062_11.INJECT1_1 = "NO";
    CCU2D add_1062_9 (.A0(d8[7]), .B0(d_d8[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[8]), .B1(d_d8[8]), .C1(GND_net), .D1(GND_net), .CIN(n11095), 
          .COUT(n11096), .S0(d9_71__N_1674[7]), .S1(d9_71__N_1674[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1062_9.INIT0 = 16'h5999;
    defparam add_1062_9.INIT1 = 16'h5999;
    defparam add_1062_9.INJECT1_0 = "NO";
    defparam add_1062_9.INJECT1_1 = "NO";
    CCU2D add_1062_7 (.A0(d8[5]), .B0(d_d8[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[6]), .B1(d_d8[6]), .C1(GND_net), .D1(GND_net), .CIN(n11094), 
          .COUT(n11095), .S0(d9_71__N_1674[5]), .S1(d9_71__N_1674[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1062_7.INIT0 = 16'h5999;
    defparam add_1062_7.INIT1 = 16'h5999;
    defparam add_1062_7.INJECT1_0 = "NO";
    defparam add_1062_7.INJECT1_1 = "NO";
    CCU2D add_1062_5 (.A0(d8[3]), .B0(d_d8[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[4]), .B1(d_d8[4]), .C1(GND_net), .D1(GND_net), .CIN(n11093), 
          .COUT(n11094), .S0(d9_71__N_1674[3]), .S1(d9_71__N_1674[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1062_5.INIT0 = 16'h5999;
    defparam add_1062_5.INIT1 = 16'h5999;
    defparam add_1062_5.INJECT1_0 = "NO";
    defparam add_1062_5.INJECT1_1 = "NO";
    CCU2D add_1062_3 (.A0(d8[1]), .B0(d_d8[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[2]), .B1(d_d8[2]), .C1(GND_net), .D1(GND_net), .CIN(n11092), 
          .COUT(n11093), .S0(d9_71__N_1674[1]), .S1(d9_71__N_1674[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1062_3.INIT0 = 16'h5999;
    defparam add_1062_3.INIT1 = 16'h5999;
    defparam add_1062_3.INJECT1_0 = "NO";
    defparam add_1062_3.INJECT1_1 = "NO";
    CCU2D add_1062_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d8[0]), .B1(d_d8[0]), .C1(GND_net), .D1(GND_net), .COUT(n11092), 
          .S1(d9_71__N_1674[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1062_1.INIT0 = 16'h0000;
    defparam add_1062_1.INIT1 = 16'h5999;
    defparam add_1062_1.INJECT1_0 = "NO";
    defparam add_1062_1.INJECT1_1 = "NO";
    CCU2D add_1057_37 (.A0(d9[35]), .B0(d_d9[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11091), 
          .S1(n6318));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1057_37.INIT0 = 16'h5999;
    defparam add_1057_37.INIT1 = 16'h0000;
    defparam add_1057_37.INJECT1_0 = "NO";
    defparam add_1057_37.INJECT1_1 = "NO";
    CCU2D add_1057_35 (.A0(d9[33]), .B0(d_d9[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[34]), .B1(d_d9[34]), .C1(GND_net), .D1(GND_net), .CIN(n11090), 
          .COUT(n11091));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1057_35.INIT0 = 16'h5999;
    defparam add_1057_35.INIT1 = 16'h5999;
    defparam add_1057_35.INJECT1_0 = "NO";
    defparam add_1057_35.INJECT1_1 = "NO";
    CCU2D add_1057_33 (.A0(d9[31]), .B0(d_d9[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[32]), .B1(d_d9[32]), .C1(GND_net), .D1(GND_net), .CIN(n11089), 
          .COUT(n11090));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1057_33.INIT0 = 16'h5999;
    defparam add_1057_33.INIT1 = 16'h5999;
    defparam add_1057_33.INJECT1_0 = "NO";
    defparam add_1057_33.INJECT1_1 = "NO";
    CCU2D add_1057_31 (.A0(d9[29]), .B0(d_d9[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[30]), .B1(d_d9[30]), .C1(GND_net), .D1(GND_net), .CIN(n11088), 
          .COUT(n11089));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1057_31.INIT0 = 16'h5999;
    defparam add_1057_31.INIT1 = 16'h5999;
    defparam add_1057_31.INJECT1_0 = "NO";
    defparam add_1057_31.INJECT1_1 = "NO";
    CCU2D add_1057_29 (.A0(d9[27]), .B0(d_d9[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[28]), .B1(d_d9[28]), .C1(GND_net), .D1(GND_net), .CIN(n11087), 
          .COUT(n11088));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1057_29.INIT0 = 16'h5999;
    defparam add_1057_29.INIT1 = 16'h5999;
    defparam add_1057_29.INJECT1_0 = "NO";
    defparam add_1057_29.INJECT1_1 = "NO";
    CCU2D add_1057_27 (.A0(d9[25]), .B0(d_d9[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[26]), .B1(d_d9[26]), .C1(GND_net), .D1(GND_net), .CIN(n11086), 
          .COUT(n11087));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1057_27.INIT0 = 16'h5999;
    defparam add_1057_27.INIT1 = 16'h5999;
    defparam add_1057_27.INJECT1_0 = "NO";
    defparam add_1057_27.INJECT1_1 = "NO";
    CCU2D add_1057_25 (.A0(d9[23]), .B0(d_d9[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[24]), .B1(d_d9[24]), .C1(GND_net), .D1(GND_net), .CIN(n11085), 
          .COUT(n11086));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1057_25.INIT0 = 16'h5999;
    defparam add_1057_25.INIT1 = 16'h5999;
    defparam add_1057_25.INJECT1_0 = "NO";
    defparam add_1057_25.INJECT1_1 = "NO";
    CCU2D add_1057_23 (.A0(d9[21]), .B0(d_d9[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[22]), .B1(d_d9[22]), .C1(GND_net), .D1(GND_net), .CIN(n11084), 
          .COUT(n11085));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1057_23.INIT0 = 16'h5999;
    defparam add_1057_23.INIT1 = 16'h5999;
    defparam add_1057_23.INJECT1_0 = "NO";
    defparam add_1057_23.INJECT1_1 = "NO";
    CCU2D add_1057_21 (.A0(d9[19]), .B0(d_d9[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[20]), .B1(d_d9[20]), .C1(GND_net), .D1(GND_net), .CIN(n11083), 
          .COUT(n11084));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1057_21.INIT0 = 16'h5999;
    defparam add_1057_21.INIT1 = 16'h5999;
    defparam add_1057_21.INJECT1_0 = "NO";
    defparam add_1057_21.INJECT1_1 = "NO";
    CCU2D add_1057_19 (.A0(d9[17]), .B0(d_d9[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[18]), .B1(d_d9[18]), .C1(GND_net), .D1(GND_net), .CIN(n11082), 
          .COUT(n11083));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1057_19.INIT0 = 16'h5999;
    defparam add_1057_19.INIT1 = 16'h5999;
    defparam add_1057_19.INJECT1_0 = "NO";
    defparam add_1057_19.INJECT1_1 = "NO";
    CCU2D add_1057_17 (.A0(d9[15]), .B0(d_d9[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[16]), .B1(d_d9[16]), .C1(GND_net), .D1(GND_net), .CIN(n11081), 
          .COUT(n11082));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1057_17.INIT0 = 16'h5999;
    defparam add_1057_17.INIT1 = 16'h5999;
    defparam add_1057_17.INJECT1_0 = "NO";
    defparam add_1057_17.INJECT1_1 = "NO";
    CCU2D add_1057_15 (.A0(d9[13]), .B0(d_d9[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[14]), .B1(d_d9[14]), .C1(GND_net), .D1(GND_net), .CIN(n11080), 
          .COUT(n11081));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1057_15.INIT0 = 16'h5999;
    defparam add_1057_15.INIT1 = 16'h5999;
    defparam add_1057_15.INJECT1_0 = "NO";
    defparam add_1057_15.INJECT1_1 = "NO";
    CCU2D add_1057_13 (.A0(d9[11]), .B0(d_d9[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[12]), .B1(d_d9[12]), .C1(GND_net), .D1(GND_net), .CIN(n11079), 
          .COUT(n11080));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1057_13.INIT0 = 16'h5999;
    defparam add_1057_13.INIT1 = 16'h5999;
    defparam add_1057_13.INJECT1_0 = "NO";
    defparam add_1057_13.INJECT1_1 = "NO";
    CCU2D add_1057_11 (.A0(d9[9]), .B0(d_d9[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[10]), .B1(d_d9[10]), .C1(GND_net), .D1(GND_net), .CIN(n11078), 
          .COUT(n11079));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1057_11.INIT0 = 16'h5999;
    defparam add_1057_11.INIT1 = 16'h5999;
    defparam add_1057_11.INJECT1_0 = "NO";
    defparam add_1057_11.INJECT1_1 = "NO";
    CCU2D add_1057_9 (.A0(d9[7]), .B0(d_d9[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[8]), .B1(d_d9[8]), .C1(GND_net), .D1(GND_net), .CIN(n11077), 
          .COUT(n11078));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1057_9.INIT0 = 16'h5999;
    defparam add_1057_9.INIT1 = 16'h5999;
    defparam add_1057_9.INJECT1_0 = "NO";
    defparam add_1057_9.INJECT1_1 = "NO";
    CCU2D add_1057_7 (.A0(d9[5]), .B0(d_d9[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[6]), .B1(d_d9[6]), .C1(GND_net), .D1(GND_net), .CIN(n11076), 
          .COUT(n11077));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1057_7.INIT0 = 16'h5999;
    defparam add_1057_7.INIT1 = 16'h5999;
    defparam add_1057_7.INJECT1_0 = "NO";
    defparam add_1057_7.INJECT1_1 = "NO";
    CCU2D add_1057_5 (.A0(d9[3]), .B0(d_d9[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[4]), .B1(d_d9[4]), .C1(GND_net), .D1(GND_net), .CIN(n11075), 
          .COUT(n11076));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1057_5.INIT0 = 16'h5999;
    defparam add_1057_5.INIT1 = 16'h5999;
    defparam add_1057_5.INJECT1_0 = "NO";
    defparam add_1057_5.INJECT1_1 = "NO";
    CCU2D add_1057_3 (.A0(d9[1]), .B0(d_d9[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[2]), .B1(d_d9[2]), .C1(GND_net), .D1(GND_net), .CIN(n11074), 
          .COUT(n11075));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1057_3.INIT0 = 16'h5999;
    defparam add_1057_3.INIT1 = 16'h5999;
    defparam add_1057_3.INJECT1_0 = "NO";
    defparam add_1057_3.INJECT1_1 = "NO";
    CCU2D add_1057_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d9[0]), .B1(d_d9[0]), .C1(GND_net), .D1(GND_net), .COUT(n11074));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1057_1.INIT0 = 16'h0000;
    defparam add_1057_1.INIT1 = 16'h5999;
    defparam add_1057_1.INJECT1_0 = "NO";
    defparam add_1057_1.INJECT1_1 = "NO";
    CCU2D add_1037_37 (.A0(d7[35]), .B0(d_d7[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11019), 
          .S0(d8_71__N_1602[35]), .S1(n5710));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1037_37.INIT0 = 16'h5999;
    defparam add_1037_37.INIT1 = 16'h0000;
    defparam add_1037_37.INJECT1_0 = "NO";
    defparam add_1037_37.INJECT1_1 = "NO";
    CCU2D add_1037_35 (.A0(d7[33]), .B0(d_d7[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[34]), .B1(d_d7[34]), .C1(GND_net), .D1(GND_net), .CIN(n11018), 
          .COUT(n11019), .S0(d8_71__N_1602[33]), .S1(d8_71__N_1602[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1037_35.INIT0 = 16'h5999;
    defparam add_1037_35.INIT1 = 16'h5999;
    defparam add_1037_35.INJECT1_0 = "NO";
    defparam add_1037_35.INJECT1_1 = "NO";
    CCU2D add_1037_33 (.A0(d7[31]), .B0(d_d7[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[32]), .B1(d_d7[32]), .C1(GND_net), .D1(GND_net), .CIN(n11017), 
          .COUT(n11018), .S0(d8_71__N_1602[31]), .S1(d8_71__N_1602[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1037_33.INIT0 = 16'h5999;
    defparam add_1037_33.INIT1 = 16'h5999;
    defparam add_1037_33.INJECT1_0 = "NO";
    defparam add_1037_33.INJECT1_1 = "NO";
    CCU2D add_1037_31 (.A0(d7[29]), .B0(d_d7[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[30]), .B1(d_d7[30]), .C1(GND_net), .D1(GND_net), .CIN(n11016), 
          .COUT(n11017), .S0(d8_71__N_1602[29]), .S1(d8_71__N_1602[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1037_31.INIT0 = 16'h5999;
    defparam add_1037_31.INIT1 = 16'h5999;
    defparam add_1037_31.INJECT1_0 = "NO";
    defparam add_1037_31.INJECT1_1 = "NO";
    CCU2D add_1037_29 (.A0(d7[27]), .B0(d_d7[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[28]), .B1(d_d7[28]), .C1(GND_net), .D1(GND_net), .CIN(n11015), 
          .COUT(n11016), .S0(d8_71__N_1602[27]), .S1(d8_71__N_1602[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1037_29.INIT0 = 16'h5999;
    defparam add_1037_29.INIT1 = 16'h5999;
    defparam add_1037_29.INJECT1_0 = "NO";
    defparam add_1037_29.INJECT1_1 = "NO";
    CCU2D add_1037_27 (.A0(d7[25]), .B0(d_d7[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[26]), .B1(d_d7[26]), .C1(GND_net), .D1(GND_net), .CIN(n11014), 
          .COUT(n11015), .S0(d8_71__N_1602[25]), .S1(d8_71__N_1602[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1037_27.INIT0 = 16'h5999;
    defparam add_1037_27.INIT1 = 16'h5999;
    defparam add_1037_27.INJECT1_0 = "NO";
    defparam add_1037_27.INJECT1_1 = "NO";
    CCU2D add_1037_25 (.A0(d7[23]), .B0(d_d7[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[24]), .B1(d_d7[24]), .C1(GND_net), .D1(GND_net), .CIN(n11013), 
          .COUT(n11014), .S0(d8_71__N_1602[23]), .S1(d8_71__N_1602[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1037_25.INIT0 = 16'h5999;
    defparam add_1037_25.INIT1 = 16'h5999;
    defparam add_1037_25.INJECT1_0 = "NO";
    defparam add_1037_25.INJECT1_1 = "NO";
    CCU2D add_1037_23 (.A0(d7[21]), .B0(d_d7[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[22]), .B1(d_d7[22]), .C1(GND_net), .D1(GND_net), .CIN(n11012), 
          .COUT(n11013), .S0(d8_71__N_1602[21]), .S1(d8_71__N_1602[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1037_23.INIT0 = 16'h5999;
    defparam add_1037_23.INIT1 = 16'h5999;
    defparam add_1037_23.INJECT1_0 = "NO";
    defparam add_1037_23.INJECT1_1 = "NO";
    CCU2D add_1037_21 (.A0(d7[19]), .B0(d_d7[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[20]), .B1(d_d7[20]), .C1(GND_net), .D1(GND_net), .CIN(n11011), 
          .COUT(n11012), .S0(d8_71__N_1602[19]), .S1(d8_71__N_1602[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1037_21.INIT0 = 16'h5999;
    defparam add_1037_21.INIT1 = 16'h5999;
    defparam add_1037_21.INJECT1_0 = "NO";
    defparam add_1037_21.INJECT1_1 = "NO";
    CCU2D add_1037_19 (.A0(d7[17]), .B0(d_d7[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[18]), .B1(d_d7[18]), .C1(GND_net), .D1(GND_net), .CIN(n11010), 
          .COUT(n11011), .S0(d8_71__N_1602[17]), .S1(d8_71__N_1602[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1037_19.INIT0 = 16'h5999;
    defparam add_1037_19.INIT1 = 16'h5999;
    defparam add_1037_19.INJECT1_0 = "NO";
    defparam add_1037_19.INJECT1_1 = "NO";
    CCU2D add_1037_17 (.A0(d7[15]), .B0(d_d7[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[16]), .B1(d_d7[16]), .C1(GND_net), .D1(GND_net), .CIN(n11009), 
          .COUT(n11010), .S0(d8_71__N_1602[15]), .S1(d8_71__N_1602[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1037_17.INIT0 = 16'h5999;
    defparam add_1037_17.INIT1 = 16'h5999;
    defparam add_1037_17.INJECT1_0 = "NO";
    defparam add_1037_17.INJECT1_1 = "NO";
    CCU2D add_1037_15 (.A0(d7[13]), .B0(d_d7[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[14]), .B1(d_d7[14]), .C1(GND_net), .D1(GND_net), .CIN(n11008), 
          .COUT(n11009), .S0(d8_71__N_1602[13]), .S1(d8_71__N_1602[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1037_15.INIT0 = 16'h5999;
    defparam add_1037_15.INIT1 = 16'h5999;
    defparam add_1037_15.INJECT1_0 = "NO";
    defparam add_1037_15.INJECT1_1 = "NO";
    CCU2D add_1037_13 (.A0(d7[11]), .B0(d_d7[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[12]), .B1(d_d7[12]), .C1(GND_net), .D1(GND_net), .CIN(n11007), 
          .COUT(n11008), .S0(d8_71__N_1602[11]), .S1(d8_71__N_1602[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1037_13.INIT0 = 16'h5999;
    defparam add_1037_13.INIT1 = 16'h5999;
    defparam add_1037_13.INJECT1_0 = "NO";
    defparam add_1037_13.INJECT1_1 = "NO";
    CCU2D add_1037_11 (.A0(d7[9]), .B0(d_d7[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[10]), .B1(d_d7[10]), .C1(GND_net), .D1(GND_net), .CIN(n11006), 
          .COUT(n11007), .S0(d8_71__N_1602[9]), .S1(d8_71__N_1602[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1037_11.INIT0 = 16'h5999;
    defparam add_1037_11.INIT1 = 16'h5999;
    defparam add_1037_11.INJECT1_0 = "NO";
    defparam add_1037_11.INJECT1_1 = "NO";
    CCU2D add_1037_9 (.A0(d7[7]), .B0(d_d7[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[8]), .B1(d_d7[8]), .C1(GND_net), .D1(GND_net), .CIN(n11005), 
          .COUT(n11006), .S0(d8_71__N_1602[7]), .S1(d8_71__N_1602[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1037_9.INIT0 = 16'h5999;
    defparam add_1037_9.INIT1 = 16'h5999;
    defparam add_1037_9.INJECT1_0 = "NO";
    defparam add_1037_9.INJECT1_1 = "NO";
    CCU2D add_1037_7 (.A0(d7[5]), .B0(d_d7[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[6]), .B1(d_d7[6]), .C1(GND_net), .D1(GND_net), .CIN(n11004), 
          .COUT(n11005), .S0(d8_71__N_1602[5]), .S1(d8_71__N_1602[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1037_7.INIT0 = 16'h5999;
    defparam add_1037_7.INIT1 = 16'h5999;
    defparam add_1037_7.INJECT1_0 = "NO";
    defparam add_1037_7.INJECT1_1 = "NO";
    CCU2D add_1037_5 (.A0(d7[3]), .B0(d_d7[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[4]), .B1(d_d7[4]), .C1(GND_net), .D1(GND_net), .CIN(n11003), 
          .COUT(n11004), .S0(d8_71__N_1602[3]), .S1(d8_71__N_1602[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1037_5.INIT0 = 16'h5999;
    defparam add_1037_5.INIT1 = 16'h5999;
    defparam add_1037_5.INJECT1_0 = "NO";
    defparam add_1037_5.INJECT1_1 = "NO";
    CCU2D add_1037_3 (.A0(d7[1]), .B0(d_d7[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[2]), .B1(d_d7[2]), .C1(GND_net), .D1(GND_net), .CIN(n11002), 
          .COUT(n11003), .S0(d8_71__N_1602[1]), .S1(d8_71__N_1602[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1037_3.INIT0 = 16'h5999;
    defparam add_1037_3.INIT1 = 16'h5999;
    defparam add_1037_3.INJECT1_0 = "NO";
    defparam add_1037_3.INJECT1_1 = "NO";
    CCU2D add_1037_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d7[0]), .B1(d_d7[0]), .C1(GND_net), .D1(GND_net), .COUT(n11002), 
          .S1(d8_71__N_1602[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1037_1.INIT0 = 16'h0000;
    defparam add_1037_1.INIT1 = 16'h5999;
    defparam add_1037_1.INJECT1_0 = "NO";
    defparam add_1037_1.INJECT1_1 = "NO";
    CCU2D add_1032_37 (.A0(d6[35]), .B0(d_d6[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10980), 
          .S0(d7_71__N_1530[35]), .S1(n5558));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1032_37.INIT0 = 16'h5999;
    defparam add_1032_37.INIT1 = 16'h0000;
    defparam add_1032_37.INJECT1_0 = "NO";
    defparam add_1032_37.INJECT1_1 = "NO";
    CCU2D add_1032_35 (.A0(d6[33]), .B0(d_d6[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[34]), .B1(d_d6[34]), .C1(GND_net), .D1(GND_net), .CIN(n10979), 
          .COUT(n10980), .S0(d7_71__N_1530[33]), .S1(d7_71__N_1530[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1032_35.INIT0 = 16'h5999;
    defparam add_1032_35.INIT1 = 16'h5999;
    defparam add_1032_35.INJECT1_0 = "NO";
    defparam add_1032_35.INJECT1_1 = "NO";
    CCU2D add_1032_33 (.A0(d6[31]), .B0(d_d6[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[32]), .B1(d_d6[32]), .C1(GND_net), .D1(GND_net), .CIN(n10978), 
          .COUT(n10979), .S0(d7_71__N_1530[31]), .S1(d7_71__N_1530[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1032_33.INIT0 = 16'h5999;
    defparam add_1032_33.INIT1 = 16'h5999;
    defparam add_1032_33.INJECT1_0 = "NO";
    defparam add_1032_33.INJECT1_1 = "NO";
    CCU2D add_1032_31 (.A0(d6[29]), .B0(d_d6[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[30]), .B1(d_d6[30]), .C1(GND_net), .D1(GND_net), .CIN(n10977), 
          .COUT(n10978), .S0(d7_71__N_1530[29]), .S1(d7_71__N_1530[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1032_31.INIT0 = 16'h5999;
    defparam add_1032_31.INIT1 = 16'h5999;
    defparam add_1032_31.INJECT1_0 = "NO";
    defparam add_1032_31.INJECT1_1 = "NO";
    CCU2D add_1032_29 (.A0(d6[27]), .B0(d_d6[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[28]), .B1(d_d6[28]), .C1(GND_net), .D1(GND_net), .CIN(n10976), 
          .COUT(n10977), .S0(d7_71__N_1530[27]), .S1(d7_71__N_1530[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1032_29.INIT0 = 16'h5999;
    defparam add_1032_29.INIT1 = 16'h5999;
    defparam add_1032_29.INJECT1_0 = "NO";
    defparam add_1032_29.INJECT1_1 = "NO";
    CCU2D add_1032_27 (.A0(d6[25]), .B0(d_d6[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[26]), .B1(d_d6[26]), .C1(GND_net), .D1(GND_net), .CIN(n10975), 
          .COUT(n10976), .S0(d7_71__N_1530[25]), .S1(d7_71__N_1530[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1032_27.INIT0 = 16'h5999;
    defparam add_1032_27.INIT1 = 16'h5999;
    defparam add_1032_27.INJECT1_0 = "NO";
    defparam add_1032_27.INJECT1_1 = "NO";
    CCU2D add_1032_25 (.A0(d6[23]), .B0(d_d6[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[24]), .B1(d_d6[24]), .C1(GND_net), .D1(GND_net), .CIN(n10974), 
          .COUT(n10975), .S0(d7_71__N_1530[23]), .S1(d7_71__N_1530[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1032_25.INIT0 = 16'h5999;
    defparam add_1032_25.INIT1 = 16'h5999;
    defparam add_1032_25.INJECT1_0 = "NO";
    defparam add_1032_25.INJECT1_1 = "NO";
    CCU2D add_1032_23 (.A0(d6[21]), .B0(d_d6[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[22]), .B1(d_d6[22]), .C1(GND_net), .D1(GND_net), .CIN(n10973), 
          .COUT(n10974), .S0(d7_71__N_1530[21]), .S1(d7_71__N_1530[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1032_23.INIT0 = 16'h5999;
    defparam add_1032_23.INIT1 = 16'h5999;
    defparam add_1032_23.INJECT1_0 = "NO";
    defparam add_1032_23.INJECT1_1 = "NO";
    CCU2D add_1032_21 (.A0(d6[19]), .B0(d_d6[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[20]), .B1(d_d6[20]), .C1(GND_net), .D1(GND_net), .CIN(n10972), 
          .COUT(n10973), .S0(d7_71__N_1530[19]), .S1(d7_71__N_1530[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1032_21.INIT0 = 16'h5999;
    defparam add_1032_21.INIT1 = 16'h5999;
    defparam add_1032_21.INJECT1_0 = "NO";
    defparam add_1032_21.INJECT1_1 = "NO";
    CCU2D add_1032_19 (.A0(d6[17]), .B0(d_d6[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[18]), .B1(d_d6[18]), .C1(GND_net), .D1(GND_net), .CIN(n10971), 
          .COUT(n10972), .S0(d7_71__N_1530[17]), .S1(d7_71__N_1530[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1032_19.INIT0 = 16'h5999;
    defparam add_1032_19.INIT1 = 16'h5999;
    defparam add_1032_19.INJECT1_0 = "NO";
    defparam add_1032_19.INJECT1_1 = "NO";
    CCU2D add_1032_17 (.A0(d6[15]), .B0(d_d6[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[16]), .B1(d_d6[16]), .C1(GND_net), .D1(GND_net), .CIN(n10970), 
          .COUT(n10971), .S0(d7_71__N_1530[15]), .S1(d7_71__N_1530[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1032_17.INIT0 = 16'h5999;
    defparam add_1032_17.INIT1 = 16'h5999;
    defparam add_1032_17.INJECT1_0 = "NO";
    defparam add_1032_17.INJECT1_1 = "NO";
    CCU2D add_1032_15 (.A0(d6[13]), .B0(d_d6[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[14]), .B1(d_d6[14]), .C1(GND_net), .D1(GND_net), .CIN(n10969), 
          .COUT(n10970), .S0(d7_71__N_1530[13]), .S1(d7_71__N_1530[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1032_15.INIT0 = 16'h5999;
    defparam add_1032_15.INIT1 = 16'h5999;
    defparam add_1032_15.INJECT1_0 = "NO";
    defparam add_1032_15.INJECT1_1 = "NO";
    CCU2D add_1032_13 (.A0(d6[11]), .B0(d_d6[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[12]), .B1(d_d6[12]), .C1(GND_net), .D1(GND_net), .CIN(n10968), 
          .COUT(n10969), .S0(d7_71__N_1530[11]), .S1(d7_71__N_1530[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1032_13.INIT0 = 16'h5999;
    defparam add_1032_13.INIT1 = 16'h5999;
    defparam add_1032_13.INJECT1_0 = "NO";
    defparam add_1032_13.INJECT1_1 = "NO";
    CCU2D add_1032_11 (.A0(d6[9]), .B0(d_d6[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[10]), .B1(d_d6[10]), .C1(GND_net), .D1(GND_net), .CIN(n10967), 
          .COUT(n10968), .S0(d7_71__N_1530[9]), .S1(d7_71__N_1530[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1032_11.INIT0 = 16'h5999;
    defparam add_1032_11.INIT1 = 16'h5999;
    defparam add_1032_11.INJECT1_0 = "NO";
    defparam add_1032_11.INJECT1_1 = "NO";
    CCU2D add_1032_9 (.A0(d6[7]), .B0(d_d6[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[8]), .B1(d_d6[8]), .C1(GND_net), .D1(GND_net), .CIN(n10966), 
          .COUT(n10967), .S0(d7_71__N_1530[7]), .S1(d7_71__N_1530[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1032_9.INIT0 = 16'h5999;
    defparam add_1032_9.INIT1 = 16'h5999;
    defparam add_1032_9.INJECT1_0 = "NO";
    defparam add_1032_9.INJECT1_1 = "NO";
    CCU2D add_1032_7 (.A0(d6[5]), .B0(d_d6[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[6]), .B1(d_d6[6]), .C1(GND_net), .D1(GND_net), .CIN(n10965), 
          .COUT(n10966), .S0(d7_71__N_1530[5]), .S1(d7_71__N_1530[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1032_7.INIT0 = 16'h5999;
    defparam add_1032_7.INIT1 = 16'h5999;
    defparam add_1032_7.INJECT1_0 = "NO";
    defparam add_1032_7.INJECT1_1 = "NO";
    CCU2D add_1032_5 (.A0(d6[3]), .B0(d_d6[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[4]), .B1(d_d6[4]), .C1(GND_net), .D1(GND_net), .CIN(n10964), 
          .COUT(n10965), .S0(d7_71__N_1530[3]), .S1(d7_71__N_1530[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1032_5.INIT0 = 16'h5999;
    defparam add_1032_5.INIT1 = 16'h5999;
    defparam add_1032_5.INJECT1_0 = "NO";
    defparam add_1032_5.INJECT1_1 = "NO";
    CCU2D add_1032_3 (.A0(d6[1]), .B0(d_d6[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[2]), .B1(d_d6[2]), .C1(GND_net), .D1(GND_net), .CIN(n10963), 
          .COUT(n10964), .S0(d7_71__N_1530[1]), .S1(d7_71__N_1530[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1032_3.INIT0 = 16'h5999;
    defparam add_1032_3.INIT1 = 16'h5999;
    defparam add_1032_3.INJECT1_0 = "NO";
    defparam add_1032_3.INJECT1_1 = "NO";
    CCU2D add_1032_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d6[0]), .B1(d_d6[0]), .C1(GND_net), .D1(GND_net), .COUT(n10963), 
          .S1(d7_71__N_1530[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1032_1.INIT0 = 16'h0000;
    defparam add_1032_1.INIT1 = 16'h5999;
    defparam add_1032_1.INJECT1_0 = "NO";
    defparam add_1032_1.INJECT1_1 = "NO";
    CCU2D add_10_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10886), 
          .S0(n375[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_17.INIT0 = 16'h5aaa;
    defparam add_10_17.INIT1 = 16'h0000;
    defparam add_10_17.INJECT1_0 = "NO";
    defparam add_10_17.INJECT1_1 = "NO";
    CCU2D add_10_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n10885), .COUT(n10886), .S0(n375[13]), .S1(n375[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_15.INIT0 = 16'h5aaa;
    defparam add_10_15.INIT1 = 16'h5aaa;
    defparam add_10_15.INJECT1_0 = "NO";
    defparam add_10_15.INJECT1_1 = "NO";
    CCU2D add_10_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n10884), .COUT(n10885), .S0(n375[11]), .S1(n375[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_13.INIT0 = 16'h5aaa;
    defparam add_10_13.INIT1 = 16'h5aaa;
    defparam add_10_13.INJECT1_0 = "NO";
    defparam add_10_13.INJECT1_1 = "NO";
    CCU2D add_10_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n10883), .COUT(n10884), .S0(n375[9]), .S1(n375[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_11.INIT0 = 16'h5aaa;
    defparam add_10_11.INIT1 = 16'h5aaa;
    defparam add_10_11.INJECT1_0 = "NO";
    defparam add_10_11.INJECT1_1 = "NO";
    CCU2D add_10_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10882), 
          .COUT(n10883), .S0(n375[7]), .S1(n375[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_9.INIT0 = 16'h5aaa;
    defparam add_10_9.INIT1 = 16'h5aaa;
    defparam add_10_9.INJECT1_0 = "NO";
    defparam add_10_9.INJECT1_1 = "NO";
    CCU2D add_10_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10881), 
          .COUT(n10882), .S0(n375[5]), .S1(n375[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_7.INIT0 = 16'h5aaa;
    defparam add_10_7.INIT1 = 16'h5aaa;
    defparam add_10_7.INJECT1_0 = "NO";
    defparam add_10_7.INJECT1_1 = "NO";
    CCU2D add_10_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10880), 
          .COUT(n10881), .S0(n375[3]), .S1(n375[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_5.INIT0 = 16'h5aaa;
    defparam add_10_5.INIT1 = 16'h5aaa;
    defparam add_10_5.INJECT1_0 = "NO";
    defparam add_10_5.INJECT1_1 = "NO";
    CCU2D add_10_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10879), 
          .COUT(n10880), .S0(n375[1]), .S1(n375[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_3.INIT0 = 16'h5aaa;
    defparam add_10_3.INIT1 = 16'h5aaa;
    defparam add_10_3.INJECT1_0 = "NO";
    defparam add_10_3.INJECT1_1 = "NO";
    CCU2D add_10_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n10879), 
          .S1(n375[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_1.INIT0 = 16'hF000;
    defparam add_10_1.INIT1 = 16'h5555;
    defparam add_10_1.INJECT1_0 = "NO";
    defparam add_10_1.INJECT1_1 = "NO";
    CCU2D add_1002_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10859), 
          .S0(n4646));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1002_cout.INIT0 = 16'h0000;
    defparam add_1002_cout.INIT1 = 16'h0000;
    defparam add_1002_cout.INJECT1_0 = "NO";
    defparam add_1002_cout.INJECT1_1 = "NO";
    CCU2D add_1002_36 (.A0(d4[34]), .B0(d5[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[35]), .B1(d5[35]), .C1(GND_net), .D1(GND_net), .CIN(n10858), 
          .COUT(n10859), .S0(d5_71__N_705[34]), .S1(d5_71__N_705[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1002_36.INIT0 = 16'h5666;
    defparam add_1002_36.INIT1 = 16'h5666;
    defparam add_1002_36.INJECT1_0 = "NO";
    defparam add_1002_36.INJECT1_1 = "NO";
    CCU2D add_1002_34 (.A0(d4[32]), .B0(d5[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[33]), .B1(d5[33]), .C1(GND_net), .D1(GND_net), .CIN(n10857), 
          .COUT(n10858), .S0(d5_71__N_705[32]), .S1(d5_71__N_705[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1002_34.INIT0 = 16'h5666;
    defparam add_1002_34.INIT1 = 16'h5666;
    defparam add_1002_34.INJECT1_0 = "NO";
    defparam add_1002_34.INJECT1_1 = "NO";
    CCU2D add_1002_32 (.A0(d4[30]), .B0(d5[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[31]), .B1(d5[31]), .C1(GND_net), .D1(GND_net), .CIN(n10856), 
          .COUT(n10857), .S0(d5_71__N_705[30]), .S1(d5_71__N_705[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1002_32.INIT0 = 16'h5666;
    defparam add_1002_32.INIT1 = 16'h5666;
    defparam add_1002_32.INJECT1_0 = "NO";
    defparam add_1002_32.INJECT1_1 = "NO";
    CCU2D add_1002_30 (.A0(d4[28]), .B0(d5[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[29]), .B1(d5[29]), .C1(GND_net), .D1(GND_net), .CIN(n10855), 
          .COUT(n10856), .S0(d5_71__N_705[28]), .S1(d5_71__N_705[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1002_30.INIT0 = 16'h5666;
    defparam add_1002_30.INIT1 = 16'h5666;
    defparam add_1002_30.INJECT1_0 = "NO";
    defparam add_1002_30.INJECT1_1 = "NO";
    CCU2D add_1002_28 (.A0(d4[26]), .B0(d5[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[27]), .B1(d5[27]), .C1(GND_net), .D1(GND_net), .CIN(n10854), 
          .COUT(n10855), .S0(d5_71__N_705[26]), .S1(d5_71__N_705[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1002_28.INIT0 = 16'h5666;
    defparam add_1002_28.INIT1 = 16'h5666;
    defparam add_1002_28.INJECT1_0 = "NO";
    defparam add_1002_28.INJECT1_1 = "NO";
    CCU2D add_1002_26 (.A0(d4[24]), .B0(d5[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[25]), .B1(d5[25]), .C1(GND_net), .D1(GND_net), .CIN(n10853), 
          .COUT(n10854), .S0(d5_71__N_705[24]), .S1(d5_71__N_705[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1002_26.INIT0 = 16'h5666;
    defparam add_1002_26.INIT1 = 16'h5666;
    defparam add_1002_26.INJECT1_0 = "NO";
    defparam add_1002_26.INJECT1_1 = "NO";
    CCU2D add_1002_24 (.A0(d4[22]), .B0(d5[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[23]), .B1(d5[23]), .C1(GND_net), .D1(GND_net), .CIN(n10852), 
          .COUT(n10853), .S0(d5_71__N_705[22]), .S1(d5_71__N_705[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1002_24.INIT0 = 16'h5666;
    defparam add_1002_24.INIT1 = 16'h5666;
    defparam add_1002_24.INJECT1_0 = "NO";
    defparam add_1002_24.INJECT1_1 = "NO";
    CCU2D add_1002_22 (.A0(d4[20]), .B0(d5[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[21]), .B1(d5[21]), .C1(GND_net), .D1(GND_net), .CIN(n10851), 
          .COUT(n10852), .S0(d5_71__N_705[20]), .S1(d5_71__N_705[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1002_22.INIT0 = 16'h5666;
    defparam add_1002_22.INIT1 = 16'h5666;
    defparam add_1002_22.INJECT1_0 = "NO";
    defparam add_1002_22.INJECT1_1 = "NO";
    CCU2D add_1002_20 (.A0(d4[18]), .B0(d5[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[19]), .B1(d5[19]), .C1(GND_net), .D1(GND_net), .CIN(n10850), 
          .COUT(n10851), .S0(d5_71__N_705[18]), .S1(d5_71__N_705[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1002_20.INIT0 = 16'h5666;
    defparam add_1002_20.INIT1 = 16'h5666;
    defparam add_1002_20.INJECT1_0 = "NO";
    defparam add_1002_20.INJECT1_1 = "NO";
    CCU2D add_1002_18 (.A0(d4[16]), .B0(d5[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[17]), .B1(d5[17]), .C1(GND_net), .D1(GND_net), .CIN(n10849), 
          .COUT(n10850), .S0(d5_71__N_705[16]), .S1(d5_71__N_705[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1002_18.INIT0 = 16'h5666;
    defparam add_1002_18.INIT1 = 16'h5666;
    defparam add_1002_18.INJECT1_0 = "NO";
    defparam add_1002_18.INJECT1_1 = "NO";
    CCU2D add_1002_16 (.A0(d4[14]), .B0(d5[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[15]), .B1(d5[15]), .C1(GND_net), .D1(GND_net), .CIN(n10848), 
          .COUT(n10849), .S0(d5_71__N_705[14]), .S1(d5_71__N_705[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1002_16.INIT0 = 16'h5666;
    defparam add_1002_16.INIT1 = 16'h5666;
    defparam add_1002_16.INJECT1_0 = "NO";
    defparam add_1002_16.INJECT1_1 = "NO";
    CCU2D add_1002_14 (.A0(d4[12]), .B0(d5[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[13]), .B1(d5[13]), .C1(GND_net), .D1(GND_net), .CIN(n10847), 
          .COUT(n10848), .S0(d5_71__N_705[12]), .S1(d5_71__N_705[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1002_14.INIT0 = 16'h5666;
    defparam add_1002_14.INIT1 = 16'h5666;
    defparam add_1002_14.INJECT1_0 = "NO";
    defparam add_1002_14.INJECT1_1 = "NO";
    CCU2D add_1002_12 (.A0(d4[10]), .B0(d5[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[11]), .B1(d5[11]), .C1(GND_net), .D1(GND_net), .CIN(n10846), 
          .COUT(n10847), .S0(d5_71__N_705[10]), .S1(d5_71__N_705[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1002_12.INIT0 = 16'h5666;
    defparam add_1002_12.INIT1 = 16'h5666;
    defparam add_1002_12.INJECT1_0 = "NO";
    defparam add_1002_12.INJECT1_1 = "NO";
    CCU2D add_1002_10 (.A0(d4[8]), .B0(d5[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[9]), .B1(d5[9]), .C1(GND_net), .D1(GND_net), .CIN(n10845), 
          .COUT(n10846), .S0(d5_71__N_705[8]), .S1(d5_71__N_705[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1002_10.INIT0 = 16'h5666;
    defparam add_1002_10.INIT1 = 16'h5666;
    defparam add_1002_10.INJECT1_0 = "NO";
    defparam add_1002_10.INJECT1_1 = "NO";
    CCU2D add_1002_8 (.A0(d4[6]), .B0(d5[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[7]), .B1(d5[7]), .C1(GND_net), .D1(GND_net), .CIN(n10844), 
          .COUT(n10845), .S0(d5_71__N_705[6]), .S1(d5_71__N_705[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1002_8.INIT0 = 16'h5666;
    defparam add_1002_8.INIT1 = 16'h5666;
    defparam add_1002_8.INJECT1_0 = "NO";
    defparam add_1002_8.INJECT1_1 = "NO";
    CCU2D add_1002_6 (.A0(d4[4]), .B0(d5[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[5]), .B1(d5[5]), .C1(GND_net), .D1(GND_net), .CIN(n10843), 
          .COUT(n10844), .S0(d5_71__N_705[4]), .S1(d5_71__N_705[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1002_6.INIT0 = 16'h5666;
    defparam add_1002_6.INIT1 = 16'h5666;
    defparam add_1002_6.INJECT1_0 = "NO";
    defparam add_1002_6.INJECT1_1 = "NO";
    CCU2D add_1002_4 (.A0(d4[2]), .B0(d5[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[3]), .B1(d5[3]), .C1(GND_net), .D1(GND_net), .CIN(n10842), 
          .COUT(n10843), .S0(d5_71__N_705[2]), .S1(d5_71__N_705[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1002_4.INIT0 = 16'h5666;
    defparam add_1002_4.INIT1 = 16'h5666;
    defparam add_1002_4.INJECT1_0 = "NO";
    defparam add_1002_4.INJECT1_1 = "NO";
    CCU2D add_1002_2 (.A0(d4[0]), .B0(d5[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[1]), .B1(d5[1]), .C1(GND_net), .D1(GND_net), .COUT(n10842), 
          .S1(d5_71__N_705[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1002_2.INIT0 = 16'h7000;
    defparam add_1002_2.INIT1 = 16'h5666;
    defparam add_1002_2.INJECT1_0 = "NO";
    defparam add_1002_2.INJECT1_1 = "NO";
    CCU2D add_997_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10840), 
          .S0(n4494));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_997_cout.INIT0 = 16'h0000;
    defparam add_997_cout.INIT1 = 16'h0000;
    defparam add_997_cout.INJECT1_0 = "NO";
    defparam add_997_cout.INJECT1_1 = "NO";
    CCU2D add_997_36 (.A0(d3[34]), .B0(d4[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[35]), .B1(d4[35]), .C1(GND_net), .D1(GND_net), .CIN(n10839), 
          .COUT(n10840), .S0(d4_71__N_633[34]), .S1(d4_71__N_633[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_997_36.INIT0 = 16'h5666;
    defparam add_997_36.INIT1 = 16'h5666;
    defparam add_997_36.INJECT1_0 = "NO";
    defparam add_997_36.INJECT1_1 = "NO";
    CCU2D add_997_34 (.A0(d3[32]), .B0(d4[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[33]), .B1(d4[33]), .C1(GND_net), .D1(GND_net), .CIN(n10838), 
          .COUT(n10839), .S0(d4_71__N_633[32]), .S1(d4_71__N_633[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_997_34.INIT0 = 16'h5666;
    defparam add_997_34.INIT1 = 16'h5666;
    defparam add_997_34.INJECT1_0 = "NO";
    defparam add_997_34.INJECT1_1 = "NO";
    CCU2D add_997_32 (.A0(d3[30]), .B0(d4[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[31]), .B1(d4[31]), .C1(GND_net), .D1(GND_net), .CIN(n10837), 
          .COUT(n10838), .S0(d4_71__N_633[30]), .S1(d4_71__N_633[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_997_32.INIT0 = 16'h5666;
    defparam add_997_32.INIT1 = 16'h5666;
    defparam add_997_32.INJECT1_0 = "NO";
    defparam add_997_32.INJECT1_1 = "NO";
    CCU2D add_997_30 (.A0(d3[28]), .B0(d4[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[29]), .B1(d4[29]), .C1(GND_net), .D1(GND_net), .CIN(n10836), 
          .COUT(n10837), .S0(d4_71__N_633[28]), .S1(d4_71__N_633[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_997_30.INIT0 = 16'h5666;
    defparam add_997_30.INIT1 = 16'h5666;
    defparam add_997_30.INJECT1_0 = "NO";
    defparam add_997_30.INJECT1_1 = "NO";
    CCU2D add_997_28 (.A0(d3[26]), .B0(d4[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[27]), .B1(d4[27]), .C1(GND_net), .D1(GND_net), .CIN(n10835), 
          .COUT(n10836), .S0(d4_71__N_633[26]), .S1(d4_71__N_633[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_997_28.INIT0 = 16'h5666;
    defparam add_997_28.INIT1 = 16'h5666;
    defparam add_997_28.INJECT1_0 = "NO";
    defparam add_997_28.INJECT1_1 = "NO";
    CCU2D add_997_26 (.A0(d3[24]), .B0(d4[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[25]), .B1(d4[25]), .C1(GND_net), .D1(GND_net), .CIN(n10834), 
          .COUT(n10835), .S0(d4_71__N_633[24]), .S1(d4_71__N_633[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_997_26.INIT0 = 16'h5666;
    defparam add_997_26.INIT1 = 16'h5666;
    defparam add_997_26.INJECT1_0 = "NO";
    defparam add_997_26.INJECT1_1 = "NO";
    CCU2D add_997_24 (.A0(d3[22]), .B0(d4[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[23]), .B1(d4[23]), .C1(GND_net), .D1(GND_net), .CIN(n10833), 
          .COUT(n10834), .S0(d4_71__N_633[22]), .S1(d4_71__N_633[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_997_24.INIT0 = 16'h5666;
    defparam add_997_24.INIT1 = 16'h5666;
    defparam add_997_24.INJECT1_0 = "NO";
    defparam add_997_24.INJECT1_1 = "NO";
    CCU2D add_997_22 (.A0(d3[20]), .B0(d4[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[21]), .B1(d4[21]), .C1(GND_net), .D1(GND_net), .CIN(n10832), 
          .COUT(n10833), .S0(d4_71__N_633[20]), .S1(d4_71__N_633[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_997_22.INIT0 = 16'h5666;
    defparam add_997_22.INIT1 = 16'h5666;
    defparam add_997_22.INJECT1_0 = "NO";
    defparam add_997_22.INJECT1_1 = "NO";
    CCU2D add_997_20 (.A0(d3[18]), .B0(d4[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[19]), .B1(d4[19]), .C1(GND_net), .D1(GND_net), .CIN(n10831), 
          .COUT(n10832), .S0(d4_71__N_633[18]), .S1(d4_71__N_633[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_997_20.INIT0 = 16'h5666;
    defparam add_997_20.INIT1 = 16'h5666;
    defparam add_997_20.INJECT1_0 = "NO";
    defparam add_997_20.INJECT1_1 = "NO";
    CCU2D add_997_18 (.A0(d3[16]), .B0(d4[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[17]), .B1(d4[17]), .C1(GND_net), .D1(GND_net), .CIN(n10830), 
          .COUT(n10831), .S0(d4_71__N_633[16]), .S1(d4_71__N_633[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_997_18.INIT0 = 16'h5666;
    defparam add_997_18.INIT1 = 16'h5666;
    defparam add_997_18.INJECT1_0 = "NO";
    defparam add_997_18.INJECT1_1 = "NO";
    CCU2D add_997_16 (.A0(d3[14]), .B0(d4[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[15]), .B1(d4[15]), .C1(GND_net), .D1(GND_net), .CIN(n10829), 
          .COUT(n10830), .S0(d4_71__N_633[14]), .S1(d4_71__N_633[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_997_16.INIT0 = 16'h5666;
    defparam add_997_16.INIT1 = 16'h5666;
    defparam add_997_16.INJECT1_0 = "NO";
    defparam add_997_16.INJECT1_1 = "NO";
    CCU2D add_997_14 (.A0(d3[12]), .B0(d4[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[13]), .B1(d4[13]), .C1(GND_net), .D1(GND_net), .CIN(n10828), 
          .COUT(n10829), .S0(d4_71__N_633[12]), .S1(d4_71__N_633[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_997_14.INIT0 = 16'h5666;
    defparam add_997_14.INIT1 = 16'h5666;
    defparam add_997_14.INJECT1_0 = "NO";
    defparam add_997_14.INJECT1_1 = "NO";
    CCU2D add_997_12 (.A0(d3[10]), .B0(d4[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[11]), .B1(d4[11]), .C1(GND_net), .D1(GND_net), .CIN(n10827), 
          .COUT(n10828), .S0(d4_71__N_633[10]), .S1(d4_71__N_633[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_997_12.INIT0 = 16'h5666;
    defparam add_997_12.INIT1 = 16'h5666;
    defparam add_997_12.INJECT1_0 = "NO";
    defparam add_997_12.INJECT1_1 = "NO";
    CCU2D add_997_10 (.A0(d3[8]), .B0(d4[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[9]), .B1(d4[9]), .C1(GND_net), .D1(GND_net), .CIN(n10826), 
          .COUT(n10827), .S0(d4_71__N_633[8]), .S1(d4_71__N_633[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_997_10.INIT0 = 16'h5666;
    defparam add_997_10.INIT1 = 16'h5666;
    defparam add_997_10.INJECT1_0 = "NO";
    defparam add_997_10.INJECT1_1 = "NO";
    CCU2D add_997_8 (.A0(d3[6]), .B0(d4[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[7]), .B1(d4[7]), .C1(GND_net), .D1(GND_net), .CIN(n10825), 
          .COUT(n10826), .S0(d4_71__N_633[6]), .S1(d4_71__N_633[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_997_8.INIT0 = 16'h5666;
    defparam add_997_8.INIT1 = 16'h5666;
    defparam add_997_8.INJECT1_0 = "NO";
    defparam add_997_8.INJECT1_1 = "NO";
    CCU2D add_997_6 (.A0(d3[4]), .B0(d4[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[5]), .B1(d4[5]), .C1(GND_net), .D1(GND_net), .CIN(n10824), 
          .COUT(n10825), .S0(d4_71__N_633[4]), .S1(d4_71__N_633[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_997_6.INIT0 = 16'h5666;
    defparam add_997_6.INIT1 = 16'h5666;
    defparam add_997_6.INJECT1_0 = "NO";
    defparam add_997_6.INJECT1_1 = "NO";
    CCU2D add_997_4 (.A0(d3[2]), .B0(d4[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[3]), .B1(d4[3]), .C1(GND_net), .D1(GND_net), .CIN(n10823), 
          .COUT(n10824), .S0(d4_71__N_633[2]), .S1(d4_71__N_633[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_997_4.INIT0 = 16'h5666;
    defparam add_997_4.INIT1 = 16'h5666;
    defparam add_997_4.INJECT1_0 = "NO";
    defparam add_997_4.INJECT1_1 = "NO";
    CCU2D add_997_2 (.A0(d3[0]), .B0(d4[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[1]), .B1(d4[1]), .C1(GND_net), .D1(GND_net), .COUT(n10823), 
          .S1(d4_71__N_633[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_997_2.INIT0 = 16'h7000;
    defparam add_997_2.INIT1 = 16'h5666;
    defparam add_997_2.INJECT1_0 = "NO";
    defparam add_997_2.INJECT1_1 = "NO";
    CCU2D add_992_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10821), 
          .S0(n4342));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_992_cout.INIT0 = 16'h0000;
    defparam add_992_cout.INIT1 = 16'h0000;
    defparam add_992_cout.INJECT1_0 = "NO";
    defparam add_992_cout.INJECT1_1 = "NO";
    CCU2D add_992_36 (.A0(d2[34]), .B0(d3[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[35]), .B1(d3[35]), .C1(GND_net), .D1(GND_net), .CIN(n10820), 
          .COUT(n10821), .S0(d3_71__N_561[34]), .S1(d3_71__N_561[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_992_36.INIT0 = 16'h5666;
    defparam add_992_36.INIT1 = 16'h5666;
    defparam add_992_36.INJECT1_0 = "NO";
    defparam add_992_36.INJECT1_1 = "NO";
    CCU2D add_992_34 (.A0(d2[32]), .B0(d3[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[33]), .B1(d3[33]), .C1(GND_net), .D1(GND_net), .CIN(n10819), 
          .COUT(n10820), .S0(d3_71__N_561[32]), .S1(d3_71__N_561[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_992_34.INIT0 = 16'h5666;
    defparam add_992_34.INIT1 = 16'h5666;
    defparam add_992_34.INJECT1_0 = "NO";
    defparam add_992_34.INJECT1_1 = "NO";
    CCU2D add_992_32 (.A0(d2[30]), .B0(d3[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[31]), .B1(d3[31]), .C1(GND_net), .D1(GND_net), .CIN(n10818), 
          .COUT(n10819), .S0(d3_71__N_561[30]), .S1(d3_71__N_561[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_992_32.INIT0 = 16'h5666;
    defparam add_992_32.INIT1 = 16'h5666;
    defparam add_992_32.INJECT1_0 = "NO";
    defparam add_992_32.INJECT1_1 = "NO";
    CCU2D add_992_30 (.A0(d2[28]), .B0(d3[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[29]), .B1(d3[29]), .C1(GND_net), .D1(GND_net), .CIN(n10817), 
          .COUT(n10818), .S0(d3_71__N_561[28]), .S1(d3_71__N_561[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_992_30.INIT0 = 16'h5666;
    defparam add_992_30.INIT1 = 16'h5666;
    defparam add_992_30.INJECT1_0 = "NO";
    defparam add_992_30.INJECT1_1 = "NO";
    CCU2D add_992_28 (.A0(d2[26]), .B0(d3[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[27]), .B1(d3[27]), .C1(GND_net), .D1(GND_net), .CIN(n10816), 
          .COUT(n10817), .S0(d3_71__N_561[26]), .S1(d3_71__N_561[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_992_28.INIT0 = 16'h5666;
    defparam add_992_28.INIT1 = 16'h5666;
    defparam add_992_28.INJECT1_0 = "NO";
    defparam add_992_28.INJECT1_1 = "NO";
    CCU2D add_992_26 (.A0(d2[24]), .B0(d3[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[25]), .B1(d3[25]), .C1(GND_net), .D1(GND_net), .CIN(n10815), 
          .COUT(n10816), .S0(d3_71__N_561[24]), .S1(d3_71__N_561[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_992_26.INIT0 = 16'h5666;
    defparam add_992_26.INIT1 = 16'h5666;
    defparam add_992_26.INJECT1_0 = "NO";
    defparam add_992_26.INJECT1_1 = "NO";
    CCU2D add_992_24 (.A0(d2[22]), .B0(d3[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[23]), .B1(d3[23]), .C1(GND_net), .D1(GND_net), .CIN(n10814), 
          .COUT(n10815), .S0(d3_71__N_561[22]), .S1(d3_71__N_561[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_992_24.INIT0 = 16'h5666;
    defparam add_992_24.INIT1 = 16'h5666;
    defparam add_992_24.INJECT1_0 = "NO";
    defparam add_992_24.INJECT1_1 = "NO";
    CCU2D add_992_22 (.A0(d2[20]), .B0(d3[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[21]), .B1(d3[21]), .C1(GND_net), .D1(GND_net), .CIN(n10813), 
          .COUT(n10814), .S0(d3_71__N_561[20]), .S1(d3_71__N_561[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_992_22.INIT0 = 16'h5666;
    defparam add_992_22.INIT1 = 16'h5666;
    defparam add_992_22.INJECT1_0 = "NO";
    defparam add_992_22.INJECT1_1 = "NO";
    CCU2D add_992_20 (.A0(d2[18]), .B0(d3[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[19]), .B1(d3[19]), .C1(GND_net), .D1(GND_net), .CIN(n10812), 
          .COUT(n10813), .S0(d3_71__N_561[18]), .S1(d3_71__N_561[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_992_20.INIT0 = 16'h5666;
    defparam add_992_20.INIT1 = 16'h5666;
    defparam add_992_20.INJECT1_0 = "NO";
    defparam add_992_20.INJECT1_1 = "NO";
    CCU2D add_992_18 (.A0(d2[16]), .B0(d3[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[17]), .B1(d3[17]), .C1(GND_net), .D1(GND_net), .CIN(n10811), 
          .COUT(n10812), .S0(d3_71__N_561[16]), .S1(d3_71__N_561[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_992_18.INIT0 = 16'h5666;
    defparam add_992_18.INIT1 = 16'h5666;
    defparam add_992_18.INJECT1_0 = "NO";
    defparam add_992_18.INJECT1_1 = "NO";
    CCU2D add_992_16 (.A0(d2[14]), .B0(d3[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[15]), .B1(d3[15]), .C1(GND_net), .D1(GND_net), .CIN(n10810), 
          .COUT(n10811), .S0(d3_71__N_561[14]), .S1(d3_71__N_561[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_992_16.INIT0 = 16'h5666;
    defparam add_992_16.INIT1 = 16'h5666;
    defparam add_992_16.INJECT1_0 = "NO";
    defparam add_992_16.INJECT1_1 = "NO";
    CCU2D add_992_14 (.A0(d2[12]), .B0(d3[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[13]), .B1(d3[13]), .C1(GND_net), .D1(GND_net), .CIN(n10809), 
          .COUT(n10810), .S0(d3_71__N_561[12]), .S1(d3_71__N_561[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_992_14.INIT0 = 16'h5666;
    defparam add_992_14.INIT1 = 16'h5666;
    defparam add_992_14.INJECT1_0 = "NO";
    defparam add_992_14.INJECT1_1 = "NO";
    CCU2D add_992_12 (.A0(d2[10]), .B0(d3[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[11]), .B1(d3[11]), .C1(GND_net), .D1(GND_net), .CIN(n10808), 
          .COUT(n10809), .S0(d3_71__N_561[10]), .S1(d3_71__N_561[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_992_12.INIT0 = 16'h5666;
    defparam add_992_12.INIT1 = 16'h5666;
    defparam add_992_12.INJECT1_0 = "NO";
    defparam add_992_12.INJECT1_1 = "NO";
    CCU2D add_992_10 (.A0(d2[8]), .B0(d3[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[9]), .B1(d3[9]), .C1(GND_net), .D1(GND_net), .CIN(n10807), 
          .COUT(n10808), .S0(d3_71__N_561[8]), .S1(d3_71__N_561[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_992_10.INIT0 = 16'h5666;
    defparam add_992_10.INIT1 = 16'h5666;
    defparam add_992_10.INJECT1_0 = "NO";
    defparam add_992_10.INJECT1_1 = "NO";
    CCU2D add_992_8 (.A0(d2[6]), .B0(d3[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[7]), .B1(d3[7]), .C1(GND_net), .D1(GND_net), .CIN(n10806), 
          .COUT(n10807), .S0(d3_71__N_561[6]), .S1(d3_71__N_561[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_992_8.INIT0 = 16'h5666;
    defparam add_992_8.INIT1 = 16'h5666;
    defparam add_992_8.INJECT1_0 = "NO";
    defparam add_992_8.INJECT1_1 = "NO";
    CCU2D add_992_6 (.A0(d2[4]), .B0(d3[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[5]), .B1(d3[5]), .C1(GND_net), .D1(GND_net), .CIN(n10805), 
          .COUT(n10806), .S0(d3_71__N_561[4]), .S1(d3_71__N_561[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_992_6.INIT0 = 16'h5666;
    defparam add_992_6.INIT1 = 16'h5666;
    defparam add_992_6.INJECT1_0 = "NO";
    defparam add_992_6.INJECT1_1 = "NO";
    CCU2D add_992_4 (.A0(d2[2]), .B0(d3[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[3]), .B1(d3[3]), .C1(GND_net), .D1(GND_net), .CIN(n10804), 
          .COUT(n10805), .S0(d3_71__N_561[2]), .S1(d3_71__N_561[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_992_4.INIT0 = 16'h5666;
    defparam add_992_4.INIT1 = 16'h5666;
    defparam add_992_4.INJECT1_0 = "NO";
    defparam add_992_4.INJECT1_1 = "NO";
    CCU2D add_992_2 (.A0(d2[0]), .B0(d3[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[1]), .B1(d3[1]), .C1(GND_net), .D1(GND_net), .COUT(n10804), 
          .S1(d3_71__N_561[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_992_2.INIT0 = 16'h7000;
    defparam add_992_2.INIT1 = 16'h5666;
    defparam add_992_2.INJECT1_0 = "NO";
    defparam add_992_2.INJECT1_1 = "NO";
    CCU2D add_987_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10802), 
          .S0(n4190));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_987_cout.INIT0 = 16'h0000;
    defparam add_987_cout.INIT1 = 16'h0000;
    defparam add_987_cout.INJECT1_0 = "NO";
    defparam add_987_cout.INJECT1_1 = "NO";
    CCU2D add_987_36 (.A0(d1[34]), .B0(d2[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[35]), .B1(d2[35]), .C1(GND_net), .D1(GND_net), .CIN(n10801), 
          .COUT(n10802), .S0(d2_71__N_489[34]), .S1(d2_71__N_489[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_987_36.INIT0 = 16'h5666;
    defparam add_987_36.INIT1 = 16'h5666;
    defparam add_987_36.INJECT1_0 = "NO";
    defparam add_987_36.INJECT1_1 = "NO";
    CCU2D add_987_34 (.A0(d1[32]), .B0(d2[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[33]), .B1(d2[33]), .C1(GND_net), .D1(GND_net), .CIN(n10800), 
          .COUT(n10801), .S0(d2_71__N_489[32]), .S1(d2_71__N_489[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_987_34.INIT0 = 16'h5666;
    defparam add_987_34.INIT1 = 16'h5666;
    defparam add_987_34.INJECT1_0 = "NO";
    defparam add_987_34.INJECT1_1 = "NO";
    CCU2D add_987_32 (.A0(d1[30]), .B0(d2[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[31]), .B1(d2[31]), .C1(GND_net), .D1(GND_net), .CIN(n10799), 
          .COUT(n10800), .S0(d2_71__N_489[30]), .S1(d2_71__N_489[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_987_32.INIT0 = 16'h5666;
    defparam add_987_32.INIT1 = 16'h5666;
    defparam add_987_32.INJECT1_0 = "NO";
    defparam add_987_32.INJECT1_1 = "NO";
    CCU2D add_987_30 (.A0(d1[28]), .B0(d2[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[29]), .B1(d2[29]), .C1(GND_net), .D1(GND_net), .CIN(n10798), 
          .COUT(n10799), .S0(d2_71__N_489[28]), .S1(d2_71__N_489[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_987_30.INIT0 = 16'h5666;
    defparam add_987_30.INIT1 = 16'h5666;
    defparam add_987_30.INJECT1_0 = "NO";
    defparam add_987_30.INJECT1_1 = "NO";
    CCU2D add_987_28 (.A0(d1[26]), .B0(d2[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[27]), .B1(d2[27]), .C1(GND_net), .D1(GND_net), .CIN(n10797), 
          .COUT(n10798), .S0(d2_71__N_489[26]), .S1(d2_71__N_489[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_987_28.INIT0 = 16'h5666;
    defparam add_987_28.INIT1 = 16'h5666;
    defparam add_987_28.INJECT1_0 = "NO";
    defparam add_987_28.INJECT1_1 = "NO";
    CCU2D add_987_26 (.A0(d1[24]), .B0(d2[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[25]), .B1(d2[25]), .C1(GND_net), .D1(GND_net), .CIN(n10796), 
          .COUT(n10797), .S0(d2_71__N_489[24]), .S1(d2_71__N_489[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_987_26.INIT0 = 16'h5666;
    defparam add_987_26.INIT1 = 16'h5666;
    defparam add_987_26.INJECT1_0 = "NO";
    defparam add_987_26.INJECT1_1 = "NO";
    CCU2D add_987_24 (.A0(d1[22]), .B0(d2[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[23]), .B1(d2[23]), .C1(GND_net), .D1(GND_net), .CIN(n10795), 
          .COUT(n10796), .S0(d2_71__N_489[22]), .S1(d2_71__N_489[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_987_24.INIT0 = 16'h5666;
    defparam add_987_24.INIT1 = 16'h5666;
    defparam add_987_24.INJECT1_0 = "NO";
    defparam add_987_24.INJECT1_1 = "NO";
    CCU2D add_987_22 (.A0(d1[20]), .B0(d2[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[21]), .B1(d2[21]), .C1(GND_net), .D1(GND_net), .CIN(n10794), 
          .COUT(n10795), .S0(d2_71__N_489[20]), .S1(d2_71__N_489[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_987_22.INIT0 = 16'h5666;
    defparam add_987_22.INIT1 = 16'h5666;
    defparam add_987_22.INJECT1_0 = "NO";
    defparam add_987_22.INJECT1_1 = "NO";
    CCU2D add_987_20 (.A0(d1[18]), .B0(d2[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[19]), .B1(d2[19]), .C1(GND_net), .D1(GND_net), .CIN(n10793), 
          .COUT(n10794), .S0(d2_71__N_489[18]), .S1(d2_71__N_489[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_987_20.INIT0 = 16'h5666;
    defparam add_987_20.INIT1 = 16'h5666;
    defparam add_987_20.INJECT1_0 = "NO";
    defparam add_987_20.INJECT1_1 = "NO";
    CCU2D add_987_18 (.A0(d1[16]), .B0(d2[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[17]), .B1(d2[17]), .C1(GND_net), .D1(GND_net), .CIN(n10792), 
          .COUT(n10793), .S0(d2_71__N_489[16]), .S1(d2_71__N_489[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_987_18.INIT0 = 16'h5666;
    defparam add_987_18.INIT1 = 16'h5666;
    defparam add_987_18.INJECT1_0 = "NO";
    defparam add_987_18.INJECT1_1 = "NO";
    CCU2D add_987_16 (.A0(d1[14]), .B0(d2[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[15]), .B1(d2[15]), .C1(GND_net), .D1(GND_net), .CIN(n10791), 
          .COUT(n10792), .S0(d2_71__N_489[14]), .S1(d2_71__N_489[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_987_16.INIT0 = 16'h5666;
    defparam add_987_16.INIT1 = 16'h5666;
    defparam add_987_16.INJECT1_0 = "NO";
    defparam add_987_16.INJECT1_1 = "NO";
    CCU2D add_987_14 (.A0(d1[12]), .B0(d2[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[13]), .B1(d2[13]), .C1(GND_net), .D1(GND_net), .CIN(n10790), 
          .COUT(n10791), .S0(d2_71__N_489[12]), .S1(d2_71__N_489[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_987_14.INIT0 = 16'h5666;
    defparam add_987_14.INIT1 = 16'h5666;
    defparam add_987_14.INJECT1_0 = "NO";
    defparam add_987_14.INJECT1_1 = "NO";
    CCU2D add_987_12 (.A0(d1[10]), .B0(d2[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[11]), .B1(d2[11]), .C1(GND_net), .D1(GND_net), .CIN(n10789), 
          .COUT(n10790), .S0(d2_71__N_489[10]), .S1(d2_71__N_489[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_987_12.INIT0 = 16'h5666;
    defparam add_987_12.INIT1 = 16'h5666;
    defparam add_987_12.INJECT1_0 = "NO";
    defparam add_987_12.INJECT1_1 = "NO";
    CCU2D add_987_10 (.A0(d1[8]), .B0(d2[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[9]), .B1(d2[9]), .C1(GND_net), .D1(GND_net), .CIN(n10788), 
          .COUT(n10789), .S0(d2_71__N_489[8]), .S1(d2_71__N_489[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_987_10.INIT0 = 16'h5666;
    defparam add_987_10.INIT1 = 16'h5666;
    defparam add_987_10.INJECT1_0 = "NO";
    defparam add_987_10.INJECT1_1 = "NO";
    CCU2D add_987_8 (.A0(d1[6]), .B0(d2[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[7]), .B1(d2[7]), .C1(GND_net), .D1(GND_net), .CIN(n10787), 
          .COUT(n10788), .S0(d2_71__N_489[6]), .S1(d2_71__N_489[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_987_8.INIT0 = 16'h5666;
    defparam add_987_8.INIT1 = 16'h5666;
    defparam add_987_8.INJECT1_0 = "NO";
    defparam add_987_8.INJECT1_1 = "NO";
    CCU2D add_987_6 (.A0(d1[4]), .B0(d2[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[5]), .B1(d2[5]), .C1(GND_net), .D1(GND_net), .CIN(n10786), 
          .COUT(n10787), .S0(d2_71__N_489[4]), .S1(d2_71__N_489[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_987_6.INIT0 = 16'h5666;
    defparam add_987_6.INIT1 = 16'h5666;
    defparam add_987_6.INJECT1_0 = "NO";
    defparam add_987_6.INJECT1_1 = "NO";
    CCU2D add_987_4 (.A0(d1[2]), .B0(d2[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[3]), .B1(d2[3]), .C1(GND_net), .D1(GND_net), .CIN(n10785), 
          .COUT(n10786), .S0(d2_71__N_489[2]), .S1(d2_71__N_489[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_987_4.INIT0 = 16'h5666;
    defparam add_987_4.INIT1 = 16'h5666;
    defparam add_987_4.INJECT1_0 = "NO";
    defparam add_987_4.INJECT1_1 = "NO";
    CCU2D add_987_2 (.A0(d1[0]), .B0(d2[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[1]), .B1(d2[1]), .C1(GND_net), .D1(GND_net), .COUT(n10785), 
          .S1(d2_71__N_489[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_987_2.INIT0 = 16'h7000;
    defparam add_987_2.INIT1 = 16'h5666;
    defparam add_987_2.INJECT1_0 = "NO";
    defparam add_987_2.INJECT1_1 = "NO";
    LUT4 shift_right_31_i210_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n70_c), .D(n138), .Z(d_out_11__N_1818[9])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i210_3_lut_4_lut.init = 16'hfe10;
    LUT4 i2666_2_lut (.A(n375[0]), .B(n31), .Z(count_15__N_1441[0])) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(86[13] 89[16])
    defparam i2666_2_lut.init = 16'hbbbb;
    LUT4 i5789_2_lut (.A(count[10]), .B(count[5]), .Z(n13238)) /* synthesis lut_function=(A (B)) */ ;
    defparam i5789_2_lut.init = 16'h8888;
    LUT4 i5857_2_lut (.A(n31), .B(n14123), .Z(n8367)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam i5857_2_lut.init = 16'hdddd;
    LUT4 i2722_2_lut (.A(n375[11]), .B(n31), .Z(count_15__N_1441[11])) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(86[13] 89[16])
    defparam i2722_2_lut.init = 16'hbbbb;
    LUT4 shift_right_31_i212_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(d10[71]), .D(n140), .Z(d_out_11__N_1818[11])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i212_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i203_3_lut_4_lut_adj_37 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63), .D(n131_adj_2576), .Z(\d_out_11__N_1818[2] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i203_3_lut_4_lut_adj_37.init = 16'hfe10;
    LUT4 i6014_then_3_lut (.A(\CICGain[1] ), .B(d10[60]), .C(d10[58]), 
         .Z(n13820)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i6014_then_3_lut.init = 16'he4e4;
    LUT4 i6014_else_3_lut (.A(n62_c), .B(\CICGain[1] ), .C(d10[59]), .Z(n13819)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i6014_else_3_lut.init = 16'he2e2;
    LUT4 shift_right_31_i204_3_lut_4_lut_adj_38 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64), .D(n132_adj_2579), .Z(\d_out_11__N_1818[3] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i204_3_lut_4_lut_adj_38.init = 16'hfe10;
    LUT4 i4_4_lut (.A(n7), .B(count[15]), .C(count[11]), .D(count[14]), 
         .Z(n12864)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i4_4_lut.init = 16'hffef;
    FD1S3AX v_comb_66_rep_190 (.D(osc_clk_enable_62), .CK(osc_clk), .Q(osc_clk_enable_496)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_190.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_189 (.D(osc_clk_enable_62), .CK(osc_clk), .Q(osc_clk_enable_446)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_189.GSR = "ENABLED";
    LUT4 i5855_4_lut (.A(n13252), .B(n13), .C(n13254), .D(n13238), .Z(d_clk_tmp_N_1830)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i5855_4_lut.init = 16'h2000;
    CCU2D add_999_17 (.A0(d4[50]), .B0(n4494), .C0(n4495[14]), .D0(d3[50]), 
          .A1(d4[51]), .B1(n4494), .C1(n4495[15]), .D1(d3[51]), .CIN(n12003), 
          .COUT(n12004), .S0(d4_71__N_633[50]), .S1(d4_71__N_633[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_999_17.INIT0 = 16'h74b8;
    defparam add_999_17.INIT1 = 16'h74b8;
    defparam add_999_17.INJECT1_0 = "NO";
    defparam add_999_17.INJECT1_1 = "NO";
    LUT4 shift_right_31_i137_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n67_c), .D(d10[65]), .Z(n137)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i137_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i133_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63_c), .D(d10[61]), .Z(n133)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i133_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i136_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66_c), .D(d10[64]), .Z(n136)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i136_3_lut_4_lut.init = 16'hf960;
    PFUMX i6054 (.BLUT(n13819), .ALUT(n13820), .C0(\CICGain[0] ), .Z(d_out_11__N_1818[1]));
    LUT4 shift_right_31_i132_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n62_c), .D(d10[60]), .Z(n132)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i132_3_lut_4_lut.init = 16'hf960;
    LUT4 i5803_4_lut (.A(count[8]), .B(count[0]), .C(count[4]), .D(count[6]), 
         .Z(n13252)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5803_4_lut.init = 16'h8000;
    LUT4 shift_right_31_i140_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n70), .D(\d10[68] ), .Z(n140_adj_2582)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i140_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i137_3_lut_4_lut_adj_39 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n67), .D(\d10[65] ), .Z(n137_adj_2585)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i137_3_lut_4_lut_adj_39.init = 16'hf960;
    LUT4 shift_right_31_i138_3_lut_4_lut_adj_40 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n68), .D(\d10[66] ), .Z(n138_adj_2588)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i138_3_lut_4_lut_adj_40.init = 16'hf960;
    LUT4 shift_right_31_i135_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65), .D(\d10[63] ), .Z(n135_adj_2591)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i135_3_lut_4_lut.init = 16'hf960;
    FD1S3AX v_comb_66_rep_188 (.D(osc_clk_enable_62), .CK(osc_clk), .Q(osc_clk_enable_396)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_188.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_187 (.D(osc_clk_enable_62), .CK(osc_clk), .Q(osc_clk_enable_346)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_187.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_186 (.D(osc_clk_enable_62), .CK(osc_clk), .Q(osc_clk_enable_296)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_186.GSR = "ENABLED";
    LUT4 shift_right_31_i136_3_lut_4_lut_adj_41 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66), .D(\d10[64] ), .Z(n136_adj_2594)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i136_3_lut_4_lut_adj_41.init = 16'hf960;
    FD1S3AX v_comb_66_rep_192 (.D(osc_clk_enable_62), .CK(osc_clk), .Q(osc_clk_enable_596)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_192.GSR = "ENABLED";
    LUT4 shift_right_31_i133_3_lut_4_lut_adj_42 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63), .D(\d10[61] ), .Z(n133_adj_2596)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i133_3_lut_4_lut_adj_42.init = 16'hf960;
    LUT4 shift_right_31_i134_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64), .D(\d10[62] ), .Z(n134_adj_2598)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i134_3_lut_4_lut.init = 16'hf960;
    PFUMX i6046 (.BLUT(n13807), .ALUT(n13808), .C0(\CICGain[1] ), .Z(\d_out_11__N_1818[10] ));
    LUT4 shift_right_31_i131_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n61), .D(\d10[59] ), .Z(n131_adj_2576)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i131_3_lut_4_lut.init = 16'hf960;
    LUT4 i1_2_lut (.A(n12864), .B(count[3]), .Z(n13)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 i4750_2_lut (.A(d2[0]), .B(d3[0]), .Z(d3_71__N_561[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4750_2_lut.init = 16'h6666;
    LUT4 shift_right_31_i132_3_lut_4_lut_adj_43 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n62), .D(\d10[60] ), .Z(n132_adj_2579)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i132_3_lut_4_lut_adj_43.init = 16'hf960;
    LUT4 i4751_2_lut (.A(d3[0]), .B(d4[0]), .Z(d4_71__N_633[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4751_2_lut.init = 16'h6666;
    PFUMX i6040 (.BLUT(n13798), .ALUT(n13799), .C0(\CICGain[0] ), .Z(d_out_11__N_1818[0]));
    LUT4 shift_right_31_i140_3_lut_4_lut_adj_44 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n70_c), .D(d10[68]), .Z(n140)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i140_3_lut_4_lut_adj_44.init = 16'hf960;
    LUT4 i4752_2_lut (.A(d4[0]), .B(d5[0]), .Z(d5_71__N_705[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4752_2_lut.init = 16'h6666;
    LUT4 shift_right_31_i135_3_lut_4_lut_adj_45 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65_c), .D(d10[63]), .Z(n135)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i135_3_lut_4_lut_adj_45.init = 16'hf960;
    FD1S3AX v_comb_66_rep_191 (.D(osc_clk_enable_62), .CK(osc_clk), .Q(osc_clk_enable_546)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_191.GSR = "ENABLED";
    LUT4 shift_right_31_i134_3_lut_4_lut_adj_46 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64_c), .D(d10[62]), .Z(n134)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i134_3_lut_4_lut_adj_46.init = 16'hf960;
    LUT4 shift_right_31_i131_3_lut_4_lut_adj_47 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n61_c), .D(d10[59]), .Z(n131)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i131_3_lut_4_lut_adj_47.init = 16'hf960;
    FD1S3AX v_comb_66_rep_185 (.D(osc_clk_enable_62), .CK(osc_clk), .Q(osc_clk_enable_246)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_185.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_184 (.D(osc_clk_enable_62), .CK(osc_clk), .Q(osc_clk_enable_196)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_184.GSR = "ENABLED";
    LUT4 shift_right_31_i206_3_lut_4_lut_adj_48 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66), .D(n134_adj_2598), .Z(\d_out_11__N_1818[5] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i206_3_lut_4_lut_adj_48.init = 16'hfe10;
    FD1S3AX v_comb_66_rep_183 (.D(osc_clk_enable_62), .CK(osc_clk), .Q(osc_clk_enable_146)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_183.GSR = "ENABLED";
    LUT4 shift_right_31_i205_3_lut_4_lut_adj_49 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65), .D(n133_adj_2596), .Z(\d_out_11__N_1818[4] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i205_3_lut_4_lut_adj_49.init = 16'hfe10;
    LUT4 shift_right_31_i207_3_lut_4_lut_adj_50 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n67), .D(n135_adj_2591), .Z(\d_out_11__N_1818[6] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i207_3_lut_4_lut_adj_50.init = 16'hfe10;
    FD1S3AX v_comb_66_rep_182 (.D(osc_clk_enable_62), .CK(osc_clk), .Q(osc_clk_enable_1395)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_182.GSR = "ENABLED";
    CCU2D add_999_15 (.A0(d4[48]), .B0(n4494), .C0(n4495[12]), .D0(d3[48]), 
          .A1(d4[49]), .B1(n4494), .C1(n4495[13]), .D1(d3[49]), .CIN(n12002), 
          .COUT(n12003), .S0(d4_71__N_633[48]), .S1(d4_71__N_633[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_999_15.INIT0 = 16'h74b8;
    defparam add_999_15.INIT1 = 16'h74b8;
    defparam add_999_15.INJECT1_0 = "NO";
    defparam add_999_15.INJECT1_1 = "NO";
    CCU2D add_999_13 (.A0(d4[46]), .B0(n4494), .C0(n4495[10]), .D0(d3[46]), 
          .A1(d4[47]), .B1(n4494), .C1(n4495[11]), .D1(d3[47]), .CIN(n12001), 
          .COUT(n12002), .S0(d4_71__N_633[46]), .S1(d4_71__N_633[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_999_13.INIT0 = 16'h74b8;
    defparam add_999_13.INIT1 = 16'h74b8;
    defparam add_999_13.INJECT1_0 = "NO";
    defparam add_999_13.INJECT1_1 = "NO";
    CCU2D add_999_11 (.A0(d4[44]), .B0(n4494), .C0(n4495[8]), .D0(d3[44]), 
          .A1(d4[45]), .B1(n4494), .C1(n4495[9]), .D1(d3[45]), .CIN(n12000), 
          .COUT(n12001), .S0(d4_71__N_633[44]), .S1(d4_71__N_633[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_999_11.INIT0 = 16'h74b8;
    defparam add_999_11.INIT1 = 16'h74b8;
    defparam add_999_11.INJECT1_0 = "NO";
    defparam add_999_11.INJECT1_1 = "NO";
    CCU2D add_999_9 (.A0(d4[42]), .B0(n4494), .C0(n4495[6]), .D0(d3[42]), 
          .A1(d4[43]), .B1(n4494), .C1(n4495[7]), .D1(d3[43]), .CIN(n11999), 
          .COUT(n12000), .S0(d4_71__N_633[42]), .S1(d4_71__N_633[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_999_9.INIT0 = 16'h74b8;
    defparam add_999_9.INIT1 = 16'h74b8;
    defparam add_999_9.INJECT1_0 = "NO";
    defparam add_999_9.INJECT1_1 = "NO";
    LUT4 shift_right_31_i208_3_lut_4_lut_adj_51 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n68), .D(n136_adj_2594), .Z(\d_out_11__N_1818[7] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i208_3_lut_4_lut_adj_51.init = 16'hfe10;
    CCU2D add_999_7 (.A0(d4[40]), .B0(n4494), .C0(n4495[4]), .D0(d3[40]), 
          .A1(d4[41]), .B1(n4494), .C1(n4495[5]), .D1(d3[41]), .CIN(n11998), 
          .COUT(n11999), .S0(d4_71__N_633[40]), .S1(d4_71__N_633[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_999_7.INIT0 = 16'h74b8;
    defparam add_999_7.INIT1 = 16'h74b8;
    defparam add_999_7.INJECT1_0 = "NO";
    defparam add_999_7.INJECT1_1 = "NO";
    CCU2D add_999_5 (.A0(d4[38]), .B0(n4494), .C0(n4495[2]), .D0(d3[38]), 
          .A1(d4[39]), .B1(n4494), .C1(n4495[3]), .D1(d3[39]), .CIN(n11997), 
          .COUT(n11998), .S0(d4_71__N_633[38]), .S1(d4_71__N_633[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_999_5.INIT0 = 16'h74b8;
    defparam add_999_5.INIT1 = 16'h74b8;
    defparam add_999_5.INJECT1_0 = "NO";
    defparam add_999_5.INJECT1_1 = "NO";
    CCU2D add_999_3 (.A0(d4[36]), .B0(n4494), .C0(n4495[0]), .D0(d3[36]), 
          .A1(d4[37]), .B1(n4494), .C1(n4495[1]), .D1(d3[37]), .CIN(n11996), 
          .COUT(n11997), .S0(d4_71__N_633[36]), .S1(d4_71__N_633[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_999_3.INIT0 = 16'h74b8;
    defparam add_999_3.INIT1 = 16'h74b8;
    defparam add_999_3.INJECT1_0 = "NO";
    defparam add_999_3.INJECT1_1 = "NO";
    LUT4 shift_right_31_i141_3_lut_4_lut_adj_52 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n137_adj_2585), .D(\d10[68] ), .Z(\d_out_11__N_1818[8] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i141_3_lut_4_lut_adj_52.init = 16'hf1e0;
    CCU2D add_999_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n4494), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11996));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_999_1.INIT0 = 16'hF000;
    defparam add_999_1.INIT1 = 16'h0555;
    defparam add_999_1.INJECT1_0 = "NO";
    defparam add_999_1.INJECT1_1 = "NO";
    CCU2D add_1003_36 (.A0(d4[70]), .B0(d5[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[71]), .B1(d5[71]), .C1(GND_net), .D1(GND_net), .CIN(n11991), 
          .S0(n4647[34]), .S1(n4647[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1003_36.INIT0 = 16'h5666;
    defparam add_1003_36.INIT1 = 16'h5666;
    defparam add_1003_36.INJECT1_0 = "NO";
    defparam add_1003_36.INJECT1_1 = "NO";
    CCU2D add_1003_34 (.A0(d4[68]), .B0(d5[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[69]), .B1(d5[69]), .C1(GND_net), .D1(GND_net), .CIN(n11990), 
          .COUT(n11991), .S0(n4647[32]), .S1(n4647[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1003_34.INIT0 = 16'h5666;
    defparam add_1003_34.INIT1 = 16'h5666;
    defparam add_1003_34.INJECT1_0 = "NO";
    defparam add_1003_34.INJECT1_1 = "NO";
    CCU2D add_1003_32 (.A0(d4[66]), .B0(d5[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[67]), .B1(d5[67]), .C1(GND_net), .D1(GND_net), .CIN(n11989), 
          .COUT(n11990), .S0(n4647[30]), .S1(n4647[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1003_32.INIT0 = 16'h5666;
    defparam add_1003_32.INIT1 = 16'h5666;
    defparam add_1003_32.INJECT1_0 = "NO";
    defparam add_1003_32.INJECT1_1 = "NO";
    CCU2D add_1003_30 (.A0(d4[64]), .B0(d5[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[65]), .B1(d5[65]), .C1(GND_net), .D1(GND_net), .CIN(n11988), 
          .COUT(n11989), .S0(n4647[28]), .S1(n4647[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1003_30.INIT0 = 16'h5666;
    defparam add_1003_30.INIT1 = 16'h5666;
    defparam add_1003_30.INJECT1_0 = "NO";
    defparam add_1003_30.INJECT1_1 = "NO";
    CCU2D add_1003_28 (.A0(d4[62]), .B0(d5[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[63]), .B1(d5[63]), .C1(GND_net), .D1(GND_net), .CIN(n11987), 
          .COUT(n11988), .S0(n4647[26]), .S1(n4647[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1003_28.INIT0 = 16'h5666;
    defparam add_1003_28.INIT1 = 16'h5666;
    defparam add_1003_28.INJECT1_0 = "NO";
    defparam add_1003_28.INJECT1_1 = "NO";
    CCU2D add_1003_26 (.A0(d4[60]), .B0(d5[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[61]), .B1(d5[61]), .C1(GND_net), .D1(GND_net), .CIN(n11986), 
          .COUT(n11987), .S0(n4647[24]), .S1(n4647[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1003_26.INIT0 = 16'h5666;
    defparam add_1003_26.INIT1 = 16'h5666;
    defparam add_1003_26.INJECT1_0 = "NO";
    defparam add_1003_26.INJECT1_1 = "NO";
    CCU2D add_1003_24 (.A0(d4[58]), .B0(d5[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[59]), .B1(d5[59]), .C1(GND_net), .D1(GND_net), .CIN(n11985), 
          .COUT(n11986), .S0(n4647[22]), .S1(n4647[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1003_24.INIT0 = 16'h5666;
    defparam add_1003_24.INIT1 = 16'h5666;
    defparam add_1003_24.INJECT1_0 = "NO";
    defparam add_1003_24.INJECT1_1 = "NO";
    CCU2D add_1003_22 (.A0(d4[56]), .B0(d5[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[57]), .B1(d5[57]), .C1(GND_net), .D1(GND_net), .CIN(n11984), 
          .COUT(n11985), .S0(n4647[20]), .S1(n4647[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1003_22.INIT0 = 16'h5666;
    defparam add_1003_22.INIT1 = 16'h5666;
    defparam add_1003_22.INJECT1_0 = "NO";
    defparam add_1003_22.INJECT1_1 = "NO";
    CCU2D add_1003_20 (.A0(d4[54]), .B0(d5[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[55]), .B1(d5[55]), .C1(GND_net), .D1(GND_net), .CIN(n11983), 
          .COUT(n11984), .S0(n4647[18]), .S1(n4647[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1003_20.INIT0 = 16'h5666;
    defparam add_1003_20.INIT1 = 16'h5666;
    defparam add_1003_20.INJECT1_0 = "NO";
    defparam add_1003_20.INJECT1_1 = "NO";
    CCU2D add_1003_18 (.A0(d4[52]), .B0(d5[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[53]), .B1(d5[53]), .C1(GND_net), .D1(GND_net), .CIN(n11982), 
          .COUT(n11983), .S0(n4647[16]), .S1(n4647[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1003_18.INIT0 = 16'h5666;
    defparam add_1003_18.INIT1 = 16'h5666;
    defparam add_1003_18.INJECT1_0 = "NO";
    defparam add_1003_18.INJECT1_1 = "NO";
    CCU2D add_1003_16 (.A0(d4[50]), .B0(d5[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[51]), .B1(d5[51]), .C1(GND_net), .D1(GND_net), .CIN(n11981), 
          .COUT(n11982), .S0(n4647[14]), .S1(n4647[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1003_16.INIT0 = 16'h5666;
    defparam add_1003_16.INIT1 = 16'h5666;
    defparam add_1003_16.INJECT1_0 = "NO";
    defparam add_1003_16.INJECT1_1 = "NO";
    CCU2D add_984_36 (.A0(MixerOutSin[11]), .B0(d1[70]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[71]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12134), .S0(n4077[34]), .S1(n4077[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_984_36.INIT0 = 16'h5666;
    defparam add_984_36.INIT1 = 16'h5666;
    defparam add_984_36.INJECT1_0 = "NO";
    defparam add_984_36.INJECT1_1 = "NO";
    CCU2D add_984_34 (.A0(MixerOutSin[11]), .B0(d1[68]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[69]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12133), .COUT(n12134), .S0(n4077[32]), 
          .S1(n4077[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_984_34.INIT0 = 16'h5666;
    defparam add_984_34.INIT1 = 16'h5666;
    defparam add_984_34.INJECT1_0 = "NO";
    defparam add_984_34.INJECT1_1 = "NO";
    CCU2D add_984_32 (.A0(MixerOutSin[11]), .B0(d1[66]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[67]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12132), .COUT(n12133), .S0(n4077[30]), 
          .S1(n4077[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_984_32.INIT0 = 16'h5666;
    defparam add_984_32.INIT1 = 16'h5666;
    defparam add_984_32.INJECT1_0 = "NO";
    defparam add_984_32.INJECT1_1 = "NO";
    CCU2D add_984_30 (.A0(MixerOutSin[11]), .B0(d1[64]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[65]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12131), .COUT(n12132), .S0(n4077[28]), 
          .S1(n4077[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_984_30.INIT0 = 16'h5666;
    defparam add_984_30.INIT1 = 16'h5666;
    defparam add_984_30.INJECT1_0 = "NO";
    defparam add_984_30.INJECT1_1 = "NO";
    CCU2D add_984_28 (.A0(MixerOutSin[11]), .B0(d1[62]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[63]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12130), .COUT(n12131), .S0(n4077[26]), 
          .S1(n4077[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_984_28.INIT0 = 16'h5666;
    defparam add_984_28.INIT1 = 16'h5666;
    defparam add_984_28.INJECT1_0 = "NO";
    defparam add_984_28.INJECT1_1 = "NO";
    CCU2D add_984_26 (.A0(MixerOutSin[11]), .B0(d1[60]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[61]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12129), .COUT(n12130), .S0(n4077[24]), 
          .S1(n4077[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_984_26.INIT0 = 16'h5666;
    defparam add_984_26.INIT1 = 16'h5666;
    defparam add_984_26.INJECT1_0 = "NO";
    defparam add_984_26.INJECT1_1 = "NO";
    CCU2D add_984_24 (.A0(MixerOutSin[11]), .B0(d1[58]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[59]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12128), .COUT(n12129), .S0(n4077[22]), 
          .S1(n4077[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_984_24.INIT0 = 16'h5666;
    defparam add_984_24.INIT1 = 16'h5666;
    defparam add_984_24.INJECT1_0 = "NO";
    defparam add_984_24.INJECT1_1 = "NO";
    CCU2D add_984_22 (.A0(MixerOutSin[11]), .B0(d1[56]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[57]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12127), .COUT(n12128), .S0(n4077[20]), 
          .S1(n4077[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_984_22.INIT0 = 16'h5666;
    defparam add_984_22.INIT1 = 16'h5666;
    defparam add_984_22.INJECT1_0 = "NO";
    defparam add_984_22.INJECT1_1 = "NO";
    CCU2D add_984_20 (.A0(MixerOutSin[11]), .B0(d1[54]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[55]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12126), .COUT(n12127), .S0(n4077[18]), 
          .S1(n4077[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_984_20.INIT0 = 16'h5666;
    defparam add_984_20.INIT1 = 16'h5666;
    defparam add_984_20.INJECT1_0 = "NO";
    defparam add_984_20.INJECT1_1 = "NO";
    CCU2D add_984_18 (.A0(MixerOutSin[11]), .B0(d1[52]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[53]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12125), .COUT(n12126), .S0(n4077[16]), 
          .S1(n4077[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_984_18.INIT0 = 16'h5666;
    defparam add_984_18.INIT1 = 16'h5666;
    defparam add_984_18.INJECT1_0 = "NO";
    defparam add_984_18.INJECT1_1 = "NO";
    LUT4 shift_right_31_i210_3_lut_4_lut_adj_53 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n70), .D(n138_adj_2588), .Z(\d_out_11__N_1818[9] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i210_3_lut_4_lut_adj_53.init = 16'hfe10;
    CCU2D add_984_16 (.A0(MixerOutSin[11]), .B0(d1[50]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[51]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12124), .COUT(n12125), .S0(n4077[14]), 
          .S1(n4077[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_984_16.INIT0 = 16'h5666;
    defparam add_984_16.INIT1 = 16'h5666;
    defparam add_984_16.INJECT1_0 = "NO";
    defparam add_984_16.INJECT1_1 = "NO";
    CCU2D add_984_14 (.A0(MixerOutSin[11]), .B0(d1[48]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[49]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12123), .COUT(n12124), .S0(n4077[12]), 
          .S1(n4077[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_984_14.INIT0 = 16'h5666;
    defparam add_984_14.INIT1 = 16'h5666;
    defparam add_984_14.INJECT1_0 = "NO";
    defparam add_984_14.INJECT1_1 = "NO";
    CCU2D add_984_12 (.A0(MixerOutSin[11]), .B0(d1[46]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[47]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12122), .COUT(n12123), .S0(n4077[10]), 
          .S1(n4077[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_984_12.INIT0 = 16'h5666;
    defparam add_984_12.INIT1 = 16'h5666;
    defparam add_984_12.INJECT1_0 = "NO";
    defparam add_984_12.INJECT1_1 = "NO";
    CCU2D add_1003_14 (.A0(d4[48]), .B0(d5[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[49]), .B1(d5[49]), .C1(GND_net), .D1(GND_net), .CIN(n11980), 
          .COUT(n11981), .S0(n4647[12]), .S1(n4647[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1003_14.INIT0 = 16'h5666;
    defparam add_1003_14.INIT1 = 16'h5666;
    defparam add_1003_14.INJECT1_0 = "NO";
    defparam add_1003_14.INJECT1_1 = "NO";
    CCU2D add_984_10 (.A0(MixerOutSin[11]), .B0(d1[44]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[45]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12121), .COUT(n12122), .S0(n4077[8]), 
          .S1(n4077[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_984_10.INIT0 = 16'h5666;
    defparam add_984_10.INIT1 = 16'h5666;
    defparam add_984_10.INJECT1_0 = "NO";
    defparam add_984_10.INJECT1_1 = "NO";
    CCU2D add_984_8 (.A0(MixerOutSin[11]), .B0(d1[42]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[43]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12120), .COUT(n12121), .S0(n4077[6]), 
          .S1(n4077[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_984_8.INIT0 = 16'h5666;
    defparam add_984_8.INIT1 = 16'h5666;
    defparam add_984_8.INJECT1_0 = "NO";
    defparam add_984_8.INJECT1_1 = "NO";
    CCU2D add_984_6 (.A0(MixerOutSin[11]), .B0(d1[40]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[41]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12119), .COUT(n12120), .S0(n4077[4]), 
          .S1(n4077[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_984_6.INIT0 = 16'h5666;
    defparam add_984_6.INIT1 = 16'h5666;
    defparam add_984_6.INJECT1_0 = "NO";
    defparam add_984_6.INJECT1_1 = "NO";
    CCU2D add_1003_12 (.A0(d4[46]), .B0(d5[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[47]), .B1(d5[47]), .C1(GND_net), .D1(GND_net), .CIN(n11979), 
          .COUT(n11980), .S0(n4647[10]), .S1(n4647[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1003_12.INIT0 = 16'h5666;
    defparam add_1003_12.INIT1 = 16'h5666;
    defparam add_1003_12.INJECT1_0 = "NO";
    defparam add_1003_12.INJECT1_1 = "NO";
    CCU2D add_984_4 (.A0(MixerOutSin[11]), .B0(d1[38]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[39]), .C1(GND_net), 
          .D1(GND_net), .CIN(n12118), .COUT(n12119), .S0(n4077[2]), 
          .S1(n4077[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_984_4.INIT0 = 16'h5666;
    defparam add_984_4.INIT1 = 16'h5666;
    defparam add_984_4.INJECT1_0 = "NO";
    defparam add_984_4.INJECT1_1 = "NO";
    CCU2D add_984_2 (.A0(MixerOutSin[11]), .B0(d1[36]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutSin[11]), .B1(d1[37]), .C1(GND_net), 
          .D1(GND_net), .COUT(n12118), .S1(n4077[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_984_2.INIT0 = 16'h1000;
    defparam add_984_2.INIT1 = 16'h5666;
    defparam add_984_2.INJECT1_0 = "NO";
    defparam add_984_2.INJECT1_1 = "NO";
    CCU2D add_1003_10 (.A0(d4[44]), .B0(d5[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[45]), .B1(d5[45]), .C1(GND_net), .D1(GND_net), .CIN(n11978), 
          .COUT(n11979), .S0(n4647[8]), .S1(n4647[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1003_10.INIT0 = 16'h5666;
    defparam add_1003_10.INIT1 = 16'h5666;
    defparam add_1003_10.INJECT1_0 = "NO";
    defparam add_1003_10.INJECT1_1 = "NO";
    CCU2D add_988_36 (.A0(d1[70]), .B0(d2[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[71]), .B1(d2[71]), .C1(GND_net), .D1(GND_net), .CIN(n12114), 
          .S0(n4191[34]), .S1(n4191[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_988_36.INIT0 = 16'h5666;
    defparam add_988_36.INIT1 = 16'h5666;
    defparam add_988_36.INJECT1_0 = "NO";
    defparam add_988_36.INJECT1_1 = "NO";
    CCU2D add_988_34 (.A0(d1[68]), .B0(d2[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[69]), .B1(d2[69]), .C1(GND_net), .D1(GND_net), .CIN(n12113), 
          .COUT(n12114), .S0(n4191[32]), .S1(n4191[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_988_34.INIT0 = 16'h5666;
    defparam add_988_34.INIT1 = 16'h5666;
    defparam add_988_34.INJECT1_0 = "NO";
    defparam add_988_34.INJECT1_1 = "NO";
    CCU2D add_1003_8 (.A0(d4[42]), .B0(d5[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[43]), .B1(d5[43]), .C1(GND_net), .D1(GND_net), .CIN(n11977), 
          .COUT(n11978), .S0(n4647[6]), .S1(n4647[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1003_8.INIT0 = 16'h5666;
    defparam add_1003_8.INIT1 = 16'h5666;
    defparam add_1003_8.INJECT1_0 = "NO";
    defparam add_1003_8.INJECT1_1 = "NO";
    CCU2D add_988_32 (.A0(d1[66]), .B0(d2[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[67]), .B1(d2[67]), .C1(GND_net), .D1(GND_net), .CIN(n12112), 
          .COUT(n12113), .S0(n4191[30]), .S1(n4191[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_988_32.INIT0 = 16'h5666;
    defparam add_988_32.INIT1 = 16'h5666;
    defparam add_988_32.INJECT1_0 = "NO";
    defparam add_988_32.INJECT1_1 = "NO";
    CCU2D add_988_30 (.A0(d1[64]), .B0(d2[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[65]), .B1(d2[65]), .C1(GND_net), .D1(GND_net), .CIN(n12111), 
          .COUT(n12112), .S0(n4191[28]), .S1(n4191[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_988_30.INIT0 = 16'h5666;
    defparam add_988_30.INIT1 = 16'h5666;
    defparam add_988_30.INJECT1_0 = "NO";
    defparam add_988_30.INJECT1_1 = "NO";
    CCU2D add_988_28 (.A0(d1[62]), .B0(d2[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[63]), .B1(d2[63]), .C1(GND_net), .D1(GND_net), .CIN(n12110), 
          .COUT(n12111), .S0(n4191[26]), .S1(n4191[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_988_28.INIT0 = 16'h5666;
    defparam add_988_28.INIT1 = 16'h5666;
    defparam add_988_28.INJECT1_0 = "NO";
    defparam add_988_28.INJECT1_1 = "NO";
    CCU2D add_988_26 (.A0(d1[60]), .B0(d2[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[61]), .B1(d2[61]), .C1(GND_net), .D1(GND_net), .CIN(n12109), 
          .COUT(n12110), .S0(n4191[24]), .S1(n4191[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_988_26.INIT0 = 16'h5666;
    defparam add_988_26.INIT1 = 16'h5666;
    defparam add_988_26.INJECT1_0 = "NO";
    defparam add_988_26.INJECT1_1 = "NO";
    CCU2D add_988_24 (.A0(d1[58]), .B0(d2[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[59]), .B1(d2[59]), .C1(GND_net), .D1(GND_net), .CIN(n12108), 
          .COUT(n12109), .S0(n4191[22]), .S1(n4191[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_988_24.INIT0 = 16'h5666;
    defparam add_988_24.INIT1 = 16'h5666;
    defparam add_988_24.INJECT1_0 = "NO";
    defparam add_988_24.INJECT1_1 = "NO";
    CCU2D add_988_22 (.A0(d1[56]), .B0(d2[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[57]), .B1(d2[57]), .C1(GND_net), .D1(GND_net), .CIN(n12107), 
          .COUT(n12108), .S0(n4191[20]), .S1(n4191[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_988_22.INIT0 = 16'h5666;
    defparam add_988_22.INIT1 = 16'h5666;
    defparam add_988_22.INJECT1_0 = "NO";
    defparam add_988_22.INJECT1_1 = "NO";
    CCU2D add_988_20 (.A0(d1[54]), .B0(d2[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[55]), .B1(d2[55]), .C1(GND_net), .D1(GND_net), .CIN(n12106), 
          .COUT(n12107), .S0(n4191[18]), .S1(n4191[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_988_20.INIT0 = 16'h5666;
    defparam add_988_20.INIT1 = 16'h5666;
    defparam add_988_20.INJECT1_0 = "NO";
    defparam add_988_20.INJECT1_1 = "NO";
    CCU2D add_988_18 (.A0(d1[52]), .B0(d2[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[53]), .B1(d2[53]), .C1(GND_net), .D1(GND_net), .CIN(n12105), 
          .COUT(n12106), .S0(n4191[16]), .S1(n4191[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_988_18.INIT0 = 16'h5666;
    defparam add_988_18.INIT1 = 16'h5666;
    defparam add_988_18.INJECT1_0 = "NO";
    defparam add_988_18.INJECT1_1 = "NO";
    CCU2D add_988_16 (.A0(d1[50]), .B0(d2[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[51]), .B1(d2[51]), .C1(GND_net), .D1(GND_net), .CIN(n12104), 
          .COUT(n12105), .S0(n4191[14]), .S1(n4191[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_988_16.INIT0 = 16'h5666;
    defparam add_988_16.INIT1 = 16'h5666;
    defparam add_988_16.INJECT1_0 = "NO";
    defparam add_988_16.INJECT1_1 = "NO";
    CCU2D add_988_14 (.A0(d1[48]), .B0(d2[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[49]), .B1(d2[49]), .C1(GND_net), .D1(GND_net), .CIN(n12103), 
          .COUT(n12104), .S0(n4191[12]), .S1(n4191[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_988_14.INIT0 = 16'h5666;
    defparam add_988_14.INIT1 = 16'h5666;
    defparam add_988_14.INJECT1_0 = "NO";
    defparam add_988_14.INJECT1_1 = "NO";
    CCU2D add_988_12 (.A0(d1[46]), .B0(d2[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[47]), .B1(d2[47]), .C1(GND_net), .D1(GND_net), .CIN(n12102), 
          .COUT(n12103), .S0(n4191[10]), .S1(n4191[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_988_12.INIT0 = 16'h5666;
    defparam add_988_12.INIT1 = 16'h5666;
    defparam add_988_12.INJECT1_0 = "NO";
    defparam add_988_12.INJECT1_1 = "NO";
    CCU2D add_988_10 (.A0(d1[44]), .B0(d2[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[45]), .B1(d2[45]), .C1(GND_net), .D1(GND_net), .CIN(n12101), 
          .COUT(n12102), .S0(n4191[8]), .S1(n4191[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_988_10.INIT0 = 16'h5666;
    defparam add_988_10.INIT1 = 16'h5666;
    defparam add_988_10.INJECT1_0 = "NO";
    defparam add_988_10.INJECT1_1 = "NO";
    CCU2D add_988_8 (.A0(d1[42]), .B0(d2[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[43]), .B1(d2[43]), .C1(GND_net), .D1(GND_net), .CIN(n12100), 
          .COUT(n12101), .S0(n4191[6]), .S1(n4191[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_988_8.INIT0 = 16'h5666;
    defparam add_988_8.INIT1 = 16'h5666;
    defparam add_988_8.INJECT1_0 = "NO";
    defparam add_988_8.INJECT1_1 = "NO";
    CCU2D add_988_6 (.A0(d1[40]), .B0(d2[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[41]), .B1(d2[41]), .C1(GND_net), .D1(GND_net), .CIN(n12099), 
          .COUT(n12100), .S0(n4191[4]), .S1(n4191[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_988_6.INIT0 = 16'h5666;
    defparam add_988_6.INIT1 = 16'h5666;
    defparam add_988_6.INJECT1_0 = "NO";
    defparam add_988_6.INJECT1_1 = "NO";
    CCU2D add_1003_6 (.A0(d4[40]), .B0(d5[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[41]), .B1(d5[41]), .C1(GND_net), .D1(GND_net), .CIN(n11976), 
          .COUT(n11977), .S0(n4647[4]), .S1(n4647[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1003_6.INIT0 = 16'h5666;
    defparam add_1003_6.INIT1 = 16'h5666;
    defparam add_1003_6.INJECT1_0 = "NO";
    defparam add_1003_6.INJECT1_1 = "NO";
    CCU2D add_988_4 (.A0(d1[38]), .B0(d2[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[39]), .B1(d2[39]), .C1(GND_net), .D1(GND_net), .CIN(n12098), 
          .COUT(n12099), .S0(n4191[2]), .S1(n4191[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_988_4.INIT0 = 16'h5666;
    defparam add_988_4.INIT1 = 16'h5666;
    defparam add_988_4.INJECT1_0 = "NO";
    defparam add_988_4.INJECT1_1 = "NO";
    CCU2D add_988_2 (.A0(d1[36]), .B0(d2[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[37]), .B1(d2[37]), .C1(GND_net), .D1(GND_net), .COUT(n12098), 
          .S1(n4191[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_988_2.INIT0 = 16'h7000;
    defparam add_988_2.INIT1 = 16'h5666;
    defparam add_988_2.INJECT1_0 = "NO";
    defparam add_988_2.INJECT1_1 = "NO";
    CCU2D add_989_37 (.A0(d2[70]), .B0(n4190), .C0(n4191[34]), .D0(d1[70]), 
          .A1(d2[71]), .B1(n4190), .C1(n4191[35]), .D1(d1[71]), .CIN(n12095), 
          .S0(d2_71__N_489[70]), .S1(d2_71__N_489[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_989_37.INIT0 = 16'h74b8;
    defparam add_989_37.INIT1 = 16'h74b8;
    defparam add_989_37.INJECT1_0 = "NO";
    defparam add_989_37.INJECT1_1 = "NO";
    CCU2D add_1034_31 (.A0(d_d6[64]), .B0(n5558), .C0(n5559[28]), .D0(d6[64]), 
          .A1(d_d6[65]), .B1(n5558), .C1(n5559[29]), .D1(d6[65]), .CIN(n11724), 
          .COUT(n11725), .S0(d7_71__N_1530[64]), .S1(d7_71__N_1530[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1034_31.INIT0 = 16'hb874;
    defparam add_1034_31.INIT1 = 16'hb874;
    defparam add_1034_31.INJECT1_0 = "NO";
    defparam add_1034_31.INJECT1_1 = "NO";
    CCU2D add_989_35 (.A0(d2[68]), .B0(n4190), .C0(n4191[32]), .D0(d1[68]), 
          .A1(d2[69]), .B1(n4190), .C1(n4191[33]), .D1(d1[69]), .CIN(n12094), 
          .COUT(n12095), .S0(d2_71__N_489[68]), .S1(d2_71__N_489[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_989_35.INIT0 = 16'h74b8;
    defparam add_989_35.INIT1 = 16'h74b8;
    defparam add_989_35.INJECT1_0 = "NO";
    defparam add_989_35.INJECT1_1 = "NO";
    LUT4 shift_right_31_i212_3_lut_4_lut_adj_54 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(\d10[71] ), .D(n140_adj_2582), .Z(\d_out_11__N_1818[11] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i212_3_lut_4_lut_adj_54.init = 16'hfe10;
    CCU2D add_1003_4 (.A0(d4[38]), .B0(d5[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[39]), .B1(d5[39]), .C1(GND_net), .D1(GND_net), .CIN(n11975), 
          .COUT(n11976), .S0(n4647[2]), .S1(n4647[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1003_4.INIT0 = 16'h5666;
    defparam add_1003_4.INIT1 = 16'h5666;
    defparam add_1003_4.INJECT1_0 = "NO";
    defparam add_1003_4.INJECT1_1 = "NO";
    CCU2D add_989_33 (.A0(d2[66]), .B0(n4190), .C0(n4191[30]), .D0(d1[66]), 
          .A1(d2[67]), .B1(n4190), .C1(n4191[31]), .D1(d1[67]), .CIN(n12093), 
          .COUT(n12094), .S0(d2_71__N_489[66]), .S1(d2_71__N_489[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_989_33.INIT0 = 16'h74b8;
    defparam add_989_33.INIT1 = 16'h74b8;
    defparam add_989_33.INJECT1_0 = "NO";
    defparam add_989_33.INJECT1_1 = "NO";
    CCU2D add_1003_2 (.A0(d4[36]), .B0(d5[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[37]), .B1(d5[37]), .C1(GND_net), .D1(GND_net), .COUT(n11975), 
          .S1(n4647[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1003_2.INIT0 = 16'h7000;
    defparam add_1003_2.INIT1 = 16'h5666;
    defparam add_1003_2.INJECT1_0 = "NO";
    defparam add_1003_2.INJECT1_1 = "NO";
    CCU2D add_1004_37 (.A0(d5[70]), .B0(n4646), .C0(n4647[34]), .D0(d4[70]), 
          .A1(d5[71]), .B1(n4646), .C1(n4647[35]), .D1(d4[71]), .CIN(n11972), 
          .S0(d5_71__N_705[70]), .S1(d5_71__N_705[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1004_37.INIT0 = 16'h74b8;
    defparam add_1004_37.INIT1 = 16'h74b8;
    defparam add_1004_37.INJECT1_0 = "NO";
    defparam add_1004_37.INJECT1_1 = "NO";
    FD1S3IX count__i1 (.D(n375[1]), .CK(osc_clk), .CD(n8367), .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=128, LSE_RLINE=134 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i1.GSR = "ENABLED";
    PFUMX i6026 (.BLUT(n13777), .ALUT(n13778), .C0(\CICGain[1] ), .Z(d_out_11__N_1818[10]));
    CCU2D add_1004_35 (.A0(d5[68]), .B0(n4646), .C0(n4647[32]), .D0(d4[68]), 
          .A1(d5[69]), .B1(n4646), .C1(n4647[33]), .D1(d4[69]), .CIN(n11971), 
          .COUT(n11972), .S0(d5_71__N_705[68]), .S1(d5_71__N_705[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1004_35.INIT0 = 16'h74b8;
    defparam add_1004_35.INIT1 = 16'h74b8;
    defparam add_1004_35.INJECT1_0 = "NO";
    defparam add_1004_35.INJECT1_1 = "NO";
    CCU2D add_1004_33 (.A0(d5[66]), .B0(n4646), .C0(n4647[30]), .D0(d4[66]), 
          .A1(d5[67]), .B1(n4646), .C1(n4647[31]), .D1(d4[67]), .CIN(n11970), 
          .COUT(n11971), .S0(d5_71__N_705[66]), .S1(d5_71__N_705[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1004_33.INIT0 = 16'h74b8;
    defparam add_1004_33.INIT1 = 16'h74b8;
    defparam add_1004_33.INJECT1_0 = "NO";
    defparam add_1004_33.INJECT1_1 = "NO";
    CCU2D add_1004_31 (.A0(d5[64]), .B0(n4646), .C0(n4647[28]), .D0(d4[64]), 
          .A1(d5[65]), .B1(n4646), .C1(n4647[29]), .D1(d4[65]), .CIN(n11969), 
          .COUT(n11970), .S0(d5_71__N_705[64]), .S1(d5_71__N_705[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1004_31.INIT0 = 16'h74b8;
    defparam add_1004_31.INIT1 = 16'h74b8;
    defparam add_1004_31.INJECT1_0 = "NO";
    defparam add_1004_31.INJECT1_1 = "NO";
    CCU2D add_1004_29 (.A0(d5[62]), .B0(n4646), .C0(n4647[26]), .D0(d4[62]), 
          .A1(d5[63]), .B1(n4646), .C1(n4647[27]), .D1(d4[63]), .CIN(n11968), 
          .COUT(n11969), .S0(d5_71__N_705[62]), .S1(d5_71__N_705[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1004_29.INIT0 = 16'h74b8;
    defparam add_1004_29.INIT1 = 16'h74b8;
    defparam add_1004_29.INJECT1_0 = "NO";
    defparam add_1004_29.INJECT1_1 = "NO";
    CCU2D add_1004_27 (.A0(d5[60]), .B0(n4646), .C0(n4647[24]), .D0(d4[60]), 
          .A1(d5[61]), .B1(n4646), .C1(n4647[25]), .D1(d4[61]), .CIN(n11967), 
          .COUT(n11968), .S0(d5_71__N_705[60]), .S1(d5_71__N_705[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1004_27.INIT0 = 16'h74b8;
    defparam add_1004_27.INIT1 = 16'h74b8;
    defparam add_1004_27.INJECT1_0 = "NO";
    defparam add_1004_27.INJECT1_1 = "NO";
    CCU2D add_1004_25 (.A0(d5[58]), .B0(n4646), .C0(n4647[22]), .D0(d4[58]), 
          .A1(d5[59]), .B1(n4646), .C1(n4647[23]), .D1(d4[59]), .CIN(n11966), 
          .COUT(n11967), .S0(d5_71__N_705[58]), .S1(d5_71__N_705[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1004_25.INIT0 = 16'h74b8;
    defparam add_1004_25.INIT1 = 16'h74b8;
    defparam add_1004_25.INJECT1_0 = "NO";
    defparam add_1004_25.INJECT1_1 = "NO";
    CCU2D add_1004_23 (.A0(d5[56]), .B0(n4646), .C0(n4647[20]), .D0(d4[56]), 
          .A1(d5[57]), .B1(n4646), .C1(n4647[21]), .D1(d4[57]), .CIN(n11965), 
          .COUT(n11966), .S0(d5_71__N_705[56]), .S1(d5_71__N_705[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1004_23.INIT0 = 16'h74b8;
    defparam add_1004_23.INIT1 = 16'h74b8;
    defparam add_1004_23.INJECT1_0 = "NO";
    defparam add_1004_23.INJECT1_1 = "NO";
    CCU2D add_1004_21 (.A0(d5[54]), .B0(n4646), .C0(n4647[18]), .D0(d4[54]), 
          .A1(d5[55]), .B1(n4646), .C1(n4647[19]), .D1(d4[55]), .CIN(n11964), 
          .COUT(n11965), .S0(d5_71__N_705[54]), .S1(d5_71__N_705[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1004_21.INIT0 = 16'h74b8;
    defparam add_1004_21.INIT1 = 16'h74b8;
    defparam add_1004_21.INJECT1_0 = "NO";
    defparam add_1004_21.INJECT1_1 = "NO";
    CCU2D add_989_31 (.A0(d2[64]), .B0(n4190), .C0(n4191[28]), .D0(d1[64]), 
          .A1(d2[65]), .B1(n4190), .C1(n4191[29]), .D1(d1[65]), .CIN(n12092), 
          .COUT(n12093), .S0(d2_71__N_489[64]), .S1(d2_71__N_489[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_989_31.INIT0 = 16'h74b8;
    defparam add_989_31.INIT1 = 16'h74b8;
    defparam add_989_31.INJECT1_0 = "NO";
    defparam add_989_31.INJECT1_1 = "NO";
    CCU2D add_1004_19 (.A0(d5[52]), .B0(n4646), .C0(n4647[16]), .D0(d4[52]), 
          .A1(d5[53]), .B1(n4646), .C1(n4647[17]), .D1(d4[53]), .CIN(n11963), 
          .COUT(n11964), .S0(d5_71__N_705[52]), .S1(d5_71__N_705[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1004_19.INIT0 = 16'h74b8;
    defparam add_1004_19.INIT1 = 16'h74b8;
    defparam add_1004_19.INJECT1_0 = "NO";
    defparam add_1004_19.INJECT1_1 = "NO";
    CCU2D add_1004_17 (.A0(d5[50]), .B0(n4646), .C0(n4647[14]), .D0(d4[50]), 
          .A1(d5[51]), .B1(n4646), .C1(n4647[15]), .D1(d4[51]), .CIN(n11962), 
          .COUT(n11963), .S0(d5_71__N_705[50]), .S1(d5_71__N_705[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1004_17.INIT0 = 16'h74b8;
    defparam add_1004_17.INIT1 = 16'h74b8;
    defparam add_1004_17.INJECT1_0 = "NO";
    defparam add_1004_17.INJECT1_1 = "NO";
    CCU2D add_1004_15 (.A0(d5[48]), .B0(n4646), .C0(n4647[12]), .D0(d4[48]), 
          .A1(d5[49]), .B1(n4646), .C1(n4647[13]), .D1(d4[49]), .CIN(n11961), 
          .COUT(n11962), .S0(d5_71__N_705[48]), .S1(d5_71__N_705[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1004_15.INIT0 = 16'h74b8;
    defparam add_1004_15.INIT1 = 16'h74b8;
    defparam add_1004_15.INJECT1_0 = "NO";
    defparam add_1004_15.INJECT1_1 = "NO";
    CCU2D add_1004_13 (.A0(d5[46]), .B0(n4646), .C0(n4647[10]), .D0(d4[46]), 
          .A1(d5[47]), .B1(n4646), .C1(n4647[11]), .D1(d4[47]), .CIN(n11960), 
          .COUT(n11961), .S0(d5_71__N_705[46]), .S1(d5_71__N_705[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1004_13.INIT0 = 16'h74b8;
    defparam add_1004_13.INIT1 = 16'h74b8;
    defparam add_1004_13.INJECT1_0 = "NO";
    defparam add_1004_13.INJECT1_1 = "NO";
    CCU2D add_1004_11 (.A0(d5[44]), .B0(n4646), .C0(n4647[8]), .D0(d4[44]), 
          .A1(d5[45]), .B1(n4646), .C1(n4647[9]), .D1(d4[45]), .CIN(n11959), 
          .COUT(n11960), .S0(d5_71__N_705[44]), .S1(d5_71__N_705[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1004_11.INIT0 = 16'h74b8;
    defparam add_1004_11.INIT1 = 16'h74b8;
    defparam add_1004_11.INJECT1_0 = "NO";
    defparam add_1004_11.INJECT1_1 = "NO";
    CCU2D add_1004_9 (.A0(d5[42]), .B0(n4646), .C0(n4647[6]), .D0(d4[42]), 
          .A1(d5[43]), .B1(n4646), .C1(n4647[7]), .D1(d4[43]), .CIN(n11958), 
          .COUT(n11959), .S0(d5_71__N_705[42]), .S1(d5_71__N_705[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1004_9.INIT0 = 16'h74b8;
    defparam add_1004_9.INIT1 = 16'h74b8;
    defparam add_1004_9.INJECT1_0 = "NO";
    defparam add_1004_9.INJECT1_1 = "NO";
    CCU2D add_1004_7 (.A0(d5[40]), .B0(n4646), .C0(n4647[4]), .D0(d4[40]), 
          .A1(d5[41]), .B1(n4646), .C1(n4647[5]), .D1(d4[41]), .CIN(n11957), 
          .COUT(n11958), .S0(d5_71__N_705[40]), .S1(d5_71__N_705[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1004_7.INIT0 = 16'h74b8;
    defparam add_1004_7.INIT1 = 16'h74b8;
    defparam add_1004_7.INJECT1_0 = "NO";
    defparam add_1004_7.INJECT1_1 = "NO";
    CCU2D add_1004_5 (.A0(d5[38]), .B0(n4646), .C0(n4647[2]), .D0(d4[38]), 
          .A1(d5[39]), .B1(n4646), .C1(n4647[3]), .D1(d4[39]), .CIN(n11956), 
          .COUT(n11957), .S0(d5_71__N_705[38]), .S1(d5_71__N_705[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1004_5.INIT0 = 16'h74b8;
    defparam add_1004_5.INIT1 = 16'h74b8;
    defparam add_1004_5.INJECT1_0 = "NO";
    defparam add_1004_5.INJECT1_1 = "NO";
    CCU2D add_1004_3 (.A0(d5[36]), .B0(n4646), .C0(n4647[0]), .D0(d4[36]), 
          .A1(d5[37]), .B1(n4646), .C1(n4647[1]), .D1(d4[37]), .CIN(n11955), 
          .COUT(n11956), .S0(d5_71__N_705[36]), .S1(d5_71__N_705[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1004_3.INIT0 = 16'h74b8;
    defparam add_1004_3.INIT1 = 16'h74b8;
    defparam add_1004_3.INJECT1_0 = "NO";
    defparam add_1004_3.INJECT1_1 = "NO";
    CCU2D add_1004_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n4646), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11955));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1004_1.INIT0 = 16'hF000;
    defparam add_1004_1.INIT1 = 16'h0555;
    defparam add_1004_1.INJECT1_0 = "NO";
    defparam add_1004_1.INJECT1_1 = "NO";
    LUT4 i2328_2_lut (.A(n31), .B(d_clk_tmp), .Z(n8331)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam i2328_2_lut.init = 16'h8888;
    CCU2D add_989_29 (.A0(d2[62]), .B0(n4190), .C0(n4191[26]), .D0(d1[62]), 
          .A1(d2[63]), .B1(n4190), .C1(n4191[27]), .D1(d1[63]), .CIN(n12091), 
          .COUT(n12092), .S0(d2_71__N_489[62]), .S1(d2_71__N_489[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_989_29.INIT0 = 16'h74b8;
    defparam add_989_29.INIT1 = 16'h74b8;
    defparam add_989_29.INJECT1_0 = "NO";
    defparam add_989_29.INJECT1_1 = "NO";
    CCU2D add_989_27 (.A0(d2[60]), .B0(n4190), .C0(n4191[24]), .D0(d1[60]), 
          .A1(d2[61]), .B1(n4190), .C1(n4191[25]), .D1(d1[61]), .CIN(n12090), 
          .COUT(n12091), .S0(d2_71__N_489[60]), .S1(d2_71__N_489[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_989_27.INIT0 = 16'h74b8;
    defparam add_989_27.INIT1 = 16'h74b8;
    defparam add_989_27.INJECT1_0 = "NO";
    defparam add_989_27.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PLL
//

module PLL (XIn_c, osc_clk, GND_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input XIn_c;
    output osc_clk;
    input GND_net;
    
    wire XIn_c /* synthesis is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(46[8:11])
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(55[8:15])
    
    EHXPLLJ PLLInst_0 (.CLKI(XIn_c), .CLKFB(osc_clk), .PHASESEL0(GND_net), 
            .PHASESEL1(GND_net), .PHASEDIR(GND_net), .PHASESTEP(GND_net), 
            .LOADREG(GND_net), .STDBY(GND_net), .PLLWAKESYNC(GND_net), 
            .RST(GND_net), .RESETC(GND_net), .RESETD(GND_net), .RESETM(GND_net), 
            .ENCLKOP(GND_net), .ENCLKOS(GND_net), .ENCLKOS2(GND_net), 
            .ENCLKOS3(GND_net), .PLLCLK(GND_net), .PLLRST(GND_net), .PLLSTB(GND_net), 
            .PLLWE(GND_net), .PLLDATI0(GND_net), .PLLDATI1(GND_net), .PLLDATI2(GND_net), 
            .PLLDATI3(GND_net), .PLLDATI4(GND_net), .PLLDATI5(GND_net), 
            .PLLDATI6(GND_net), .PLLDATI7(GND_net), .PLLADDR0(GND_net), 
            .PLLADDR1(GND_net), .PLLADDR2(GND_net), .PLLADDR3(GND_net), 
            .PLLADDR4(GND_net), .CLKOP(osc_clk)) /* synthesis FREQUENCY_PIN_CLKOP="80.000000", FREQUENCY_PIN_CLKI="8.000000", ICP_CURRENT="7", LPF_RESISTOR="8", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=154, LSE_RLINE=156 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(154[5] 156[2])
    defparam PLLInst_0.CLKI_DIV = 1;
    defparam PLLInst_0.CLKFB_DIV = 10;
    defparam PLLInst_0.CLKOP_DIV = 6;
    defparam PLLInst_0.CLKOS_DIV = 1;
    defparam PLLInst_0.CLKOS2_DIV = 1;
    defparam PLLInst_0.CLKOS3_DIV = 1;
    defparam PLLInst_0.CLKOP_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS2_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS3_ENABLE = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_A0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_B0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_C0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_D0 = "DISABLED";
    defparam PLLInst_0.CLKOP_CPHASE = 5;
    defparam PLLInst_0.CLKOS_CPHASE = 0;
    defparam PLLInst_0.CLKOS2_CPHASE = 0;
    defparam PLLInst_0.CLKOS3_CPHASE = 0;
    defparam PLLInst_0.CLKOP_FPHASE = 0;
    defparam PLLInst_0.CLKOS_FPHASE = 0;
    defparam PLLInst_0.CLKOS2_FPHASE = 0;
    defparam PLLInst_0.CLKOS3_FPHASE = 0;
    defparam PLLInst_0.FEEDBK_PATH = "CLKOP";
    defparam PLLInst_0.FRACN_ENABLE = "DISABLED";
    defparam PLLInst_0.FRACN_DIV = 0;
    defparam PLLInst_0.CLKOP_TRIM_POL = "RISING";
    defparam PLLInst_0.CLKOP_TRIM_DELAY = 0;
    defparam PLLInst_0.CLKOS_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOS_TRIM_DELAY = 0;
    defparam PLLInst_0.PLL_USE_WB = "DISABLED";
    defparam PLLInst_0.PREDIVIDER_MUXA1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXB1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXC1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXD1 = 0;
    defparam PLLInst_0.OUTDIVIDER_MUXA2 = "DIVA";
    defparam PLLInst_0.OUTDIVIDER_MUXB2 = "DIVB";
    defparam PLLInst_0.OUTDIVIDER_MUXC2 = "DIVC";
    defparam PLLInst_0.OUTDIVIDER_MUXD2 = "DIVD";
    defparam PLLInst_0.PLL_LOCK_MODE = 0;
    defparam PLLInst_0.STDBY_ENABLE = "DISABLED";
    defparam PLLInst_0.DPHASE_SOURCE = "DISABLED";
    defparam PLLInst_0.PLLRST_ENA = "DISABLED";
    defparam PLLInst_0.MRST_ENA = "DISABLED";
    defparam PLLInst_0.DCRST_ENA = "DISABLED";
    defparam PLLInst_0.DDRST_ENA = "DISABLED";
    defparam PLLInst_0.INTFB_WAKE = "DISABLED";
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module nco_sig
//

module nco_sig (osc_clk, \phase_accum[63] , \phase_accum[62] , \phase_accum[61] , 
            \phase_accum[60] , \phase_accum[59] , \phase_accum[58] , \phase_accum[57] , 
            \phase_accum[56] , sinGen_c, phase_inc_carrGen1, GND_net) /* synthesis syn_module_defined=1 */ ;
    input osc_clk;
    output \phase_accum[63] ;
    output \phase_accum[62] ;
    output \phase_accum[61] ;
    output \phase_accum[60] ;
    output \phase_accum[59] ;
    output \phase_accum[58] ;
    output \phase_accum[57] ;
    output \phase_accum[56] ;
    output sinGen_c;
    input [63:0]phase_inc_carrGen1;
    input GND_net;
    
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(55[8:15])
    wire [63:0]phase_accum;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(29[19:30])
    wire [63:0]phase_accum_63__N_145;
    
    wire n10782, n10781, n10780, n10779, n10778, n10777, n10776, 
        n10775, n10774, n10773, n10772, n10771, n10770, n10769, 
        n10768, n10767, n10766, n10765, n10764, n10763, n10762, 
        n10761, n10760, n10759, n10758, n10757, n10756, n10755, 
        n10754, n10753, n10752;
    
    FD1S3AX phase_accum_i0 (.D(phase_accum_63__N_145[0]), .CK(osc_clk), 
            .Q(phase_accum[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i0.GSR = "ENABLED";
    FD1S3AX phase_accum_i63 (.D(phase_accum_63__N_145[63]), .CK(osc_clk), 
            .Q(\phase_accum[63] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i63.GSR = "ENABLED";
    FD1S3AX phase_accum_i62 (.D(phase_accum_63__N_145[62]), .CK(osc_clk), 
            .Q(\phase_accum[62] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i62.GSR = "ENABLED";
    FD1S3AX phase_accum_i61 (.D(phase_accum_63__N_145[61]), .CK(osc_clk), 
            .Q(\phase_accum[61] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i61.GSR = "ENABLED";
    FD1S3AX phase_accum_i60 (.D(phase_accum_63__N_145[60]), .CK(osc_clk), 
            .Q(\phase_accum[60] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i60.GSR = "ENABLED";
    FD1S3AX phase_accum_i59 (.D(phase_accum_63__N_145[59]), .CK(osc_clk), 
            .Q(\phase_accum[59] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i59.GSR = "ENABLED";
    FD1S3AX phase_accum_i58 (.D(phase_accum_63__N_145[58]), .CK(osc_clk), 
            .Q(\phase_accum[58] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i58.GSR = "ENABLED";
    FD1S3AX phase_accum_i57 (.D(phase_accum_63__N_145[57]), .CK(osc_clk), 
            .Q(\phase_accum[57] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i57.GSR = "ENABLED";
    FD1S3AX phase_accum_i56 (.D(phase_accum_63__N_145[56]), .CK(osc_clk), 
            .Q(\phase_accum[56] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i56.GSR = "ENABLED";
    FD1S3AX phase_accum_i55 (.D(phase_accum_63__N_145[55]), .CK(osc_clk), 
            .Q(phase_accum[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i55.GSR = "ENABLED";
    FD1S3AX phase_accum_i54 (.D(phase_accum_63__N_145[54]), .CK(osc_clk), 
            .Q(phase_accum[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i54.GSR = "ENABLED";
    FD1S3AX phase_accum_i53 (.D(phase_accum_63__N_145[53]), .CK(osc_clk), 
            .Q(phase_accum[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i53.GSR = "ENABLED";
    FD1S3AX phase_accum_i52 (.D(phase_accum_63__N_145[52]), .CK(osc_clk), 
            .Q(phase_accum[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i52.GSR = "ENABLED";
    FD1S3AX phase_accum_i51 (.D(phase_accum_63__N_145[51]), .CK(osc_clk), 
            .Q(phase_accum[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i51.GSR = "ENABLED";
    FD1S3AX phase_accum_i50 (.D(phase_accum_63__N_145[50]), .CK(osc_clk), 
            .Q(phase_accum[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i50.GSR = "ENABLED";
    FD1S3AX phase_accum_i49 (.D(phase_accum_63__N_145[49]), .CK(osc_clk), 
            .Q(phase_accum[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i49.GSR = "ENABLED";
    FD1S3AX phase_accum_i48 (.D(phase_accum_63__N_145[48]), .CK(osc_clk), 
            .Q(phase_accum[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i48.GSR = "ENABLED";
    FD1S3AX phase_accum_i47 (.D(phase_accum_63__N_145[47]), .CK(osc_clk), 
            .Q(phase_accum[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i47.GSR = "ENABLED";
    FD1S3AX phase_accum_i46 (.D(phase_accum_63__N_145[46]), .CK(osc_clk), 
            .Q(phase_accum[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i46.GSR = "ENABLED";
    FD1S3AX phase_accum_i45 (.D(phase_accum_63__N_145[45]), .CK(osc_clk), 
            .Q(phase_accum[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i45.GSR = "ENABLED";
    FD1S3AX phase_accum_i44 (.D(phase_accum_63__N_145[44]), .CK(osc_clk), 
            .Q(phase_accum[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i44.GSR = "ENABLED";
    FD1S3AX phase_accum_i43 (.D(phase_accum_63__N_145[43]), .CK(osc_clk), 
            .Q(phase_accum[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i43.GSR = "ENABLED";
    FD1S3AX phase_accum_i42 (.D(phase_accum_63__N_145[42]), .CK(osc_clk), 
            .Q(phase_accum[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i42.GSR = "ENABLED";
    FD1S3AX phase_accum_i41 (.D(phase_accum_63__N_145[41]), .CK(osc_clk), 
            .Q(phase_accum[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i41.GSR = "ENABLED";
    FD1S3AX phase_accum_i40 (.D(phase_accum_63__N_145[40]), .CK(osc_clk), 
            .Q(phase_accum[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i40.GSR = "ENABLED";
    FD1S3AX phase_accum_i39 (.D(phase_accum_63__N_145[39]), .CK(osc_clk), 
            .Q(phase_accum[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i39.GSR = "ENABLED";
    FD1S3AX phase_accum_i38 (.D(phase_accum_63__N_145[38]), .CK(osc_clk), 
            .Q(phase_accum[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i38.GSR = "ENABLED";
    FD1S3AX phase_accum_i37 (.D(phase_accum_63__N_145[37]), .CK(osc_clk), 
            .Q(phase_accum[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i37.GSR = "ENABLED";
    FD1S3AX phase_accum_i36 (.D(phase_accum_63__N_145[36]), .CK(osc_clk), 
            .Q(phase_accum[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i36.GSR = "ENABLED";
    FD1S3AX phase_accum_i35 (.D(phase_accum_63__N_145[35]), .CK(osc_clk), 
            .Q(phase_accum[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i35.GSR = "ENABLED";
    FD1S3AX phase_accum_i34 (.D(phase_accum_63__N_145[34]), .CK(osc_clk), 
            .Q(phase_accum[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i34.GSR = "ENABLED";
    FD1S3AX phase_accum_i33 (.D(phase_accum_63__N_145[33]), .CK(osc_clk), 
            .Q(phase_accum[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i33.GSR = "ENABLED";
    FD1S3AX phase_accum_i32 (.D(phase_accum_63__N_145[32]), .CK(osc_clk), 
            .Q(phase_accum[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i32.GSR = "ENABLED";
    FD1S3AX phase_accum_i31 (.D(phase_accum_63__N_145[31]), .CK(osc_clk), 
            .Q(phase_accum[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i31.GSR = "ENABLED";
    FD1S3AX phase_accum_i30 (.D(phase_accum_63__N_145[30]), .CK(osc_clk), 
            .Q(phase_accum[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i30.GSR = "ENABLED";
    FD1S3AX phase_accum_i29 (.D(phase_accum_63__N_145[29]), .CK(osc_clk), 
            .Q(phase_accum[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i29.GSR = "ENABLED";
    FD1S3AX phase_accum_i28 (.D(phase_accum_63__N_145[28]), .CK(osc_clk), 
            .Q(phase_accum[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i28.GSR = "ENABLED";
    FD1S3AX phase_accum_i27 (.D(phase_accum_63__N_145[27]), .CK(osc_clk), 
            .Q(phase_accum[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i27.GSR = "ENABLED";
    FD1S3AX phase_accum_i26 (.D(phase_accum_63__N_145[26]), .CK(osc_clk), 
            .Q(phase_accum[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i26.GSR = "ENABLED";
    FD1S3AX phase_accum_i25 (.D(phase_accum_63__N_145[25]), .CK(osc_clk), 
            .Q(phase_accum[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i25.GSR = "ENABLED";
    FD1S3AX phase_accum_i24 (.D(phase_accum_63__N_145[24]), .CK(osc_clk), 
            .Q(phase_accum[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i24.GSR = "ENABLED";
    FD1S3AX phase_accum_i23 (.D(phase_accum_63__N_145[23]), .CK(osc_clk), 
            .Q(phase_accum[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i23.GSR = "ENABLED";
    FD1S3AX phase_accum_i22 (.D(phase_accum_63__N_145[22]), .CK(osc_clk), 
            .Q(phase_accum[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i22.GSR = "ENABLED";
    FD1S3AX phase_accum_i21 (.D(phase_accum_63__N_145[21]), .CK(osc_clk), 
            .Q(phase_accum[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i21.GSR = "ENABLED";
    FD1S3AX phase_accum_i20 (.D(phase_accum_63__N_145[20]), .CK(osc_clk), 
            .Q(phase_accum[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i20.GSR = "ENABLED";
    FD1S3AX phase_accum_i19 (.D(phase_accum_63__N_145[19]), .CK(osc_clk), 
            .Q(phase_accum[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i19.GSR = "ENABLED";
    FD1S3AX phase_accum_i18 (.D(phase_accum_63__N_145[18]), .CK(osc_clk), 
            .Q(phase_accum[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i18.GSR = "ENABLED";
    FD1S3AX phase_accum_i17 (.D(phase_accum_63__N_145[17]), .CK(osc_clk), 
            .Q(phase_accum[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i17.GSR = "ENABLED";
    FD1S3AX phase_accum_i16 (.D(phase_accum_63__N_145[16]), .CK(osc_clk), 
            .Q(phase_accum[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i16.GSR = "ENABLED";
    FD1S3AX phase_accum_i15 (.D(phase_accum_63__N_145[15]), .CK(osc_clk), 
            .Q(phase_accum[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i15.GSR = "ENABLED";
    FD1S3AX phase_accum_i14 (.D(phase_accum_63__N_145[14]), .CK(osc_clk), 
            .Q(phase_accum[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i14.GSR = "ENABLED";
    FD1S3AX phase_accum_i13 (.D(phase_accum_63__N_145[13]), .CK(osc_clk), 
            .Q(phase_accum[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i13.GSR = "ENABLED";
    LUT4 phase_accum_63__I_0_13_1_lut (.A(\phase_accum[63] ), .Z(sinGen_c)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(32[18:56])
    defparam phase_accum_63__I_0_13_1_lut.init = 16'h5555;
    FD1S3AX phase_accum_i12 (.D(phase_accum_63__N_145[12]), .CK(osc_clk), 
            .Q(phase_accum[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i12.GSR = "ENABLED";
    FD1S3AX phase_accum_i11 (.D(phase_accum_63__N_145[11]), .CK(osc_clk), 
            .Q(phase_accum[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i11.GSR = "ENABLED";
    FD1S3AX phase_accum_i10 (.D(phase_accum_63__N_145[10]), .CK(osc_clk), 
            .Q(phase_accum[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i10.GSR = "ENABLED";
    FD1S3AX phase_accum_i9 (.D(phase_accum_63__N_145[9]), .CK(osc_clk), 
            .Q(phase_accum[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i9.GSR = "ENABLED";
    FD1S3AX phase_accum_i8 (.D(phase_accum_63__N_145[8]), .CK(osc_clk), 
            .Q(phase_accum[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i8.GSR = "ENABLED";
    FD1S3AX phase_accum_i7 (.D(phase_accum_63__N_145[7]), .CK(osc_clk), 
            .Q(phase_accum[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i7.GSR = "ENABLED";
    FD1S3AX phase_accum_i6 (.D(phase_accum_63__N_145[6]), .CK(osc_clk), 
            .Q(phase_accum[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i6.GSR = "ENABLED";
    FD1S3AX phase_accum_i5 (.D(phase_accum_63__N_145[5]), .CK(osc_clk), 
            .Q(phase_accum[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i5.GSR = "ENABLED";
    FD1S3AX phase_accum_i4 (.D(phase_accum_63__N_145[4]), .CK(osc_clk), 
            .Q(phase_accum[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i4.GSR = "ENABLED";
    FD1S3AX phase_accum_i3 (.D(phase_accum_63__N_145[3]), .CK(osc_clk), 
            .Q(phase_accum[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i3.GSR = "ENABLED";
    FD1S3AX phase_accum_i2 (.D(phase_accum_63__N_145[2]), .CK(osc_clk), 
            .Q(phase_accum[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i2.GSR = "ENABLED";
    FD1S3AX phase_accum_i1 (.D(phase_accum_63__N_145[1]), .CK(osc_clk), 
            .Q(phase_accum[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(36[7] 38[4])
    defparam phase_accum_i1.GSR = "ENABLED";
    LUT4 i4748_2_lut (.A(phase_accum[0]), .B(phase_inc_carrGen1[0]), .Z(phase_accum_63__N_145[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4748_2_lut.init = 16'h6666;
    CCU2D phase_accum_63__I_0_12_64 (.A0(\phase_accum[62] ), .B0(phase_inc_carrGen1[62]), 
          .C0(GND_net), .D0(GND_net), .A1(\phase_accum[63] ), .B1(phase_inc_carrGen1[63]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10782), .S0(phase_accum_63__N_145[62]), 
          .S1(phase_accum_63__N_145[63]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_64.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_64.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_64.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_64.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_62 (.A0(\phase_accum[60] ), .B0(phase_inc_carrGen1[60]), 
          .C0(GND_net), .D0(GND_net), .A1(\phase_accum[61] ), .B1(phase_inc_carrGen1[61]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10781), .COUT(n10782), .S0(phase_accum_63__N_145[60]), 
          .S1(phase_accum_63__N_145[61]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_62.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_62.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_62.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_62.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_60 (.A0(\phase_accum[58] ), .B0(phase_inc_carrGen1[58]), 
          .C0(GND_net), .D0(GND_net), .A1(\phase_accum[59] ), .B1(phase_inc_carrGen1[59]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10780), .COUT(n10781), .S0(phase_accum_63__N_145[58]), 
          .S1(phase_accum_63__N_145[59]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_60.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_60.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_60.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_60.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_58 (.A0(\phase_accum[56] ), .B0(phase_inc_carrGen1[56]), 
          .C0(GND_net), .D0(GND_net), .A1(\phase_accum[57] ), .B1(phase_inc_carrGen1[57]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10779), .COUT(n10780), .S0(phase_accum_63__N_145[56]), 
          .S1(phase_accum_63__N_145[57]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_58.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_58.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_58.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_58.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_56 (.A0(phase_accum[54]), .B0(phase_inc_carrGen1[54]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[55]), .B1(phase_inc_carrGen1[55]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10778), .COUT(n10779), .S0(phase_accum_63__N_145[54]), 
          .S1(phase_accum_63__N_145[55]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_56.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_56.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_56.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_56.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_54 (.A0(phase_accum[52]), .B0(phase_inc_carrGen1[52]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[53]), .B1(phase_inc_carrGen1[53]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10777), .COUT(n10778), .S0(phase_accum_63__N_145[52]), 
          .S1(phase_accum_63__N_145[53]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_54.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_54.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_54.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_54.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_52 (.A0(phase_accum[50]), .B0(phase_inc_carrGen1[50]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[51]), .B1(phase_inc_carrGen1[51]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10776), .COUT(n10777), .S0(phase_accum_63__N_145[50]), 
          .S1(phase_accum_63__N_145[51]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_52.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_52.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_52.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_52.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_50 (.A0(phase_accum[48]), .B0(phase_inc_carrGen1[48]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[49]), .B1(phase_inc_carrGen1[49]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10775), .COUT(n10776), .S0(phase_accum_63__N_145[48]), 
          .S1(phase_accum_63__N_145[49]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_50.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_50.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_50.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_50.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_48 (.A0(phase_accum[46]), .B0(phase_inc_carrGen1[46]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[47]), .B1(phase_inc_carrGen1[47]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10774), .COUT(n10775), .S0(phase_accum_63__N_145[46]), 
          .S1(phase_accum_63__N_145[47]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_48.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_48.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_48.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_48.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_46 (.A0(phase_accum[44]), .B0(phase_inc_carrGen1[44]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[45]), .B1(phase_inc_carrGen1[45]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10773), .COUT(n10774), .S0(phase_accum_63__N_145[44]), 
          .S1(phase_accum_63__N_145[45]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_46.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_46.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_46.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_46.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_44 (.A0(phase_accum[42]), .B0(phase_inc_carrGen1[42]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[43]), .B1(phase_inc_carrGen1[43]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10772), .COUT(n10773), .S0(phase_accum_63__N_145[42]), 
          .S1(phase_accum_63__N_145[43]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_44.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_44.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_44.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_44.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_42 (.A0(phase_accum[40]), .B0(phase_inc_carrGen1[40]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[41]), .B1(phase_inc_carrGen1[41]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10771), .COUT(n10772), .S0(phase_accum_63__N_145[40]), 
          .S1(phase_accum_63__N_145[41]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_42.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_42.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_42.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_42.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_40 (.A0(phase_accum[38]), .B0(phase_inc_carrGen1[38]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[39]), .B1(phase_inc_carrGen1[39]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10770), .COUT(n10771), .S0(phase_accum_63__N_145[38]), 
          .S1(phase_accum_63__N_145[39]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_40.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_40.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_40.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_40.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_38 (.A0(phase_accum[36]), .B0(phase_inc_carrGen1[36]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[37]), .B1(phase_inc_carrGen1[37]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10769), .COUT(n10770), .S0(phase_accum_63__N_145[36]), 
          .S1(phase_accum_63__N_145[37]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_38.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_38.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_38.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_38.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_36 (.A0(phase_accum[34]), .B0(phase_inc_carrGen1[34]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[35]), .B1(phase_inc_carrGen1[35]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10768), .COUT(n10769), .S0(phase_accum_63__N_145[34]), 
          .S1(phase_accum_63__N_145[35]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_36.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_36.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_36.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_36.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_34 (.A0(phase_accum[32]), .B0(phase_inc_carrGen1[32]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[33]), .B1(phase_inc_carrGen1[33]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10767), .COUT(n10768), .S0(phase_accum_63__N_145[32]), 
          .S1(phase_accum_63__N_145[33]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_34.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_34.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_34.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_34.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_32 (.A0(phase_accum[30]), .B0(phase_inc_carrGen1[30]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[31]), .B1(phase_inc_carrGen1[31]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10766), .COUT(n10767), .S0(phase_accum_63__N_145[30]), 
          .S1(phase_accum_63__N_145[31]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_32.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_32.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_32.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_32.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_30 (.A0(phase_accum[28]), .B0(phase_inc_carrGen1[28]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[29]), .B1(phase_inc_carrGen1[29]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10765), .COUT(n10766), .S0(phase_accum_63__N_145[28]), 
          .S1(phase_accum_63__N_145[29]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_30.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_30.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_30.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_30.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_28 (.A0(phase_accum[26]), .B0(phase_inc_carrGen1[26]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[27]), .B1(phase_inc_carrGen1[27]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10764), .COUT(n10765), .S0(phase_accum_63__N_145[26]), 
          .S1(phase_accum_63__N_145[27]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_28.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_28.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_28.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_28.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_26 (.A0(phase_accum[24]), .B0(phase_inc_carrGen1[24]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[25]), .B1(phase_inc_carrGen1[25]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10763), .COUT(n10764), .S0(phase_accum_63__N_145[24]), 
          .S1(phase_accum_63__N_145[25]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_26.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_26.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_26.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_26.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_24 (.A0(phase_accum[22]), .B0(phase_inc_carrGen1[22]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[23]), .B1(phase_inc_carrGen1[23]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10762), .COUT(n10763), .S0(phase_accum_63__N_145[22]), 
          .S1(phase_accum_63__N_145[23]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_24.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_24.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_24.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_24.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_22 (.A0(phase_accum[20]), .B0(phase_inc_carrGen1[20]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[21]), .B1(phase_inc_carrGen1[21]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10761), .COUT(n10762), .S0(phase_accum_63__N_145[20]), 
          .S1(phase_accum_63__N_145[21]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_22.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_22.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_22.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_22.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_20 (.A0(phase_accum[18]), .B0(phase_inc_carrGen1[18]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[19]), .B1(phase_inc_carrGen1[19]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10760), .COUT(n10761), .S0(phase_accum_63__N_145[18]), 
          .S1(phase_accum_63__N_145[19]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_20.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_20.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_20.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_20.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_18 (.A0(phase_accum[16]), .B0(phase_inc_carrGen1[16]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[17]), .B1(phase_inc_carrGen1[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10759), .COUT(n10760), .S0(phase_accum_63__N_145[16]), 
          .S1(phase_accum_63__N_145[17]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_18.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_18.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_18.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_18.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_16 (.A0(phase_accum[14]), .B0(phase_inc_carrGen1[14]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[15]), .B1(phase_inc_carrGen1[15]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10758), .COUT(n10759), .S0(phase_accum_63__N_145[14]), 
          .S1(phase_accum_63__N_145[15]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_16.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_16.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_16.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_16.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_14 (.A0(phase_accum[12]), .B0(phase_inc_carrGen1[12]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[13]), .B1(phase_inc_carrGen1[13]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10757), .COUT(n10758), .S0(phase_accum_63__N_145[12]), 
          .S1(phase_accum_63__N_145[13]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_14.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_14.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_14.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_14.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_12 (.A0(phase_accum[10]), .B0(phase_inc_carrGen1[10]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[11]), .B1(phase_inc_carrGen1[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10756), .COUT(n10757), .S0(phase_accum_63__N_145[10]), 
          .S1(phase_accum_63__N_145[11]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_12.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_12.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_12.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_12.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_10 (.A0(phase_accum[8]), .B0(phase_inc_carrGen1[8]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[9]), .B1(phase_inc_carrGen1[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10755), .COUT(n10756), .S0(phase_accum_63__N_145[8]), 
          .S1(phase_accum_63__N_145[9]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_10.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_10.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_10.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_10.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_8 (.A0(phase_accum[6]), .B0(phase_inc_carrGen1[6]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[7]), .B1(phase_inc_carrGen1[7]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10754), .COUT(n10755), .S0(phase_accum_63__N_145[6]), 
          .S1(phase_accum_63__N_145[7]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_8.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_8.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_8.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_8.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_6 (.A0(phase_accum[4]), .B0(phase_inc_carrGen1[4]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[5]), .B1(phase_inc_carrGen1[5]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10753), .COUT(n10754), .S0(phase_accum_63__N_145[4]), 
          .S1(phase_accum_63__N_145[5]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_6.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_6.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_6.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_6.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_4 (.A0(phase_accum[2]), .B0(phase_inc_carrGen1[2]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[3]), .B1(phase_inc_carrGen1[3]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10752), .COUT(n10753), .S0(phase_accum_63__N_145[2]), 
          .S1(phase_accum_63__N_145[3]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_4.INIT0 = 16'h5666;
    defparam phase_accum_63__I_0_12_4.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_4.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_4.INJECT1_1 = "NO";
    CCU2D phase_accum_63__I_0_12_2 (.A0(phase_accum[0]), .B0(phase_inc_carrGen1[0]), 
          .C0(GND_net), .D0(GND_net), .A1(phase_accum[1]), .B1(phase_inc_carrGen1[1]), 
          .C1(GND_net), .D1(GND_net), .COUT(n10752), .S1(phase_accum_63__N_145[1]));   // c:/users/user/lattice/1bitadcfpgasdr/nco.v(37[17:45])
    defparam phase_accum_63__I_0_12_2.INIT0 = 16'h7000;
    defparam phase_accum_63__I_0_12_2.INIT1 = 16'h5666;
    defparam phase_accum_63__I_0_12_2.INJECT1_0 = "NO";
    defparam phase_accum_63__I_0_12_2.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \CIC(width=72,decimation_ratio=4096)_U1 
//

module \CIC(width=72,decimation_ratio=4096)_U1  (GND_net, osc_clk, CIC1_outCos, 
            \d10[59] , \d10[60] , \d10[61] , \d10[62] , \d10[63] , 
            \d10[64] , \d10[65] , \d10[66] , \d10[67] , \d10[68] , 
            \d10[69] , \d10[70] , \d10[71] , \d_out_11__N_1818[2] , 
            \d_out_11__N_1818[3] , \d_out_11__N_1818[4] , \d_out_11__N_1818[5] , 
            \d_out_11__N_1818[6] , \d_out_11__N_1818[7] , \d_out_11__N_1818[8] , 
            \d_out_11__N_1818[9] , \d_out_11__N_1818[10] , \d_out_11__N_1818[11] , 
            \CICGain[0] , n61, MixerOutCos, n62, n63, n64, \CICGain[1] , 
            n65, n66, n67, n68, n70) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input osc_clk;
    output [11:0]CIC1_outCos;
    output \d10[59] ;
    output \d10[60] ;
    output \d10[61] ;
    output \d10[62] ;
    output \d10[63] ;
    output \d10[64] ;
    output \d10[65] ;
    output \d10[66] ;
    output \d10[67] ;
    output \d10[68] ;
    output \d10[69] ;
    output \d10[70] ;
    output \d10[71] ;
    input \d_out_11__N_1818[2] ;
    input \d_out_11__N_1818[3] ;
    input \d_out_11__N_1818[4] ;
    input \d_out_11__N_1818[5] ;
    input \d_out_11__N_1818[6] ;
    input \d_out_11__N_1818[7] ;
    input \d_out_11__N_1818[8] ;
    input \d_out_11__N_1818[9] ;
    input \d_out_11__N_1818[10] ;
    input \d_out_11__N_1818[11] ;
    input \CICGain[0] ;
    output n61;
    input [11:0]MixerOutCos;
    output n62;
    output n63;
    output n64;
    input \CICGain[1] ;
    output n65;
    output n66;
    output n67;
    output n68;
    output n70;
    
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(55[8:15])
    
    wire n11845;
    wire [71:0]d3;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(37[26:28])
    
    wire n5102;
    wire [35:0]n5103;
    wire [71:0]d2;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(36[26:28])
    wire [71:0]d3_71__N_561;
    
    wire n11846, n11842, n11843, n11839, n11840, n11841, n11844, 
        n11893;
    wire [71:0]d1;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(35[26:28])
    wire [35:0]n4951;
    
    wire n11894;
    wire [71:0]d_tmp;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(30[26:31])
    
    wire osc_clk_enable_743;
    wire [71:0]d5;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(39[26:28])
    wire [71:0]d_d_tmp;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(30[33:40])
    
    wire osc_clk_enable_783;
    wire [71:0]d2_71__N_489;
    wire [71:0]d4;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(38[26:28])
    wire [71:0]d4_71__N_633;
    wire [71:0]d5_71__N_705;
    wire [71:0]d6;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(43[26:28])
    wire [71:0]d6_71__N_1458;
    wire [71:0]d_d6;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(43[30:34])
    
    wire v_comb;
    wire [71:0]d7;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(44[26:28])
    wire [71:0]d7_71__N_1530;
    wire [71:0]d_d7;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(44[30:34])
    wire [71:0]d8;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(45[26:28])
    wire [71:0]d8_71__N_1602;
    wire [71:0]d_d8;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(45[30:34])
    wire [71:0]d9;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(46[26:28])
    wire [71:0]d9_71__N_1674;
    wire [71:0]d_d9;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(46[30:34])
    wire [71:0]d_out_11__N_1818;
    wire [71:0]d1_71__N_417;
    
    wire n11888, n4950, n11889, n11886, n11887, n11885, n11884, 
        n11883, n11882, n11881, n11880, n11837, n11838, n11890, 
        n11833, n11834, n11825;
    wire [35:0]n5255;
    
    wire n11826, n11795, n5254, n11796, n11824, n11832, n11435;
    wire [35:0]n6167;
    
    wire n11436, n11823, n11836, n11821, n11822, n11820, n11819, 
        n11818, n11815, n11816, n11812, n11813, n11794, n11814, 
        n11817, n11811, n11793, n11827, n11792, n11835, n11434, 
        n11433, n11432, n11431, n11791, n11786;
    wire [35:0]n5407;
    
    wire n11785, n11805, n11806, n11799, n11800, n11784, n11798, 
        n11804, n11797, n11803, n11808, n11802, n11801, n11807, 
        n11879, n11878, n11783, n11877, n11875, n11876, n11873, 
        n11874, n11429, n6166, n11428, n11427, n11426, n11425, 
        n11424, n11423, n11422, n11421, n11420, n11419, n11782, 
        n11781, n11780, n11779, n11778, n11777, n11776, n12867;
    wire [15:0]count;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(50[14:19])
    
    wire n16, n13248, n13, n13250, n13228, count_15__N_1457, n31, 
        n14125, n8412;
    wire [15:0]count_15__N_1441;
    
    wire n11903, n11904, n11902, n11901, n11775, n11774;
    wire [15:0]n375;
    
    wire n11773, n11772, n11771, n11770, n11767, n5406, n11766, 
        n11765, n11764, n11763, n11762, n11761, n11760, n11759, 
        n11758, n11757, n11756, n11755, n11754, n11753, n11752, 
        n11751, n11750, n11418, osc_clk_enable_833, osc_clk_enable_883, 
        osc_clk_enable_933, osc_clk_enable_983, osc_clk_enable_1033, osc_clk_enable_1083, 
        osc_clk_enable_1133, osc_clk_enable_1183, osc_clk_enable_1233, 
        osc_clk_enable_1283, osc_clk_enable_1333, osc_clk_enable_1383;
    wire [71:0]d10;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(47[26:29])
    wire [71:0]d10_71__N_1746;
    
    wire n11417, n11416, n11415, n11414, n11413, n11412, n7, n11332;
    wire [35:0]n6623;
    
    wire n11331, n11330, n11329, n11328, n11327, n11326, n11325, 
        n11324, n11323, n11322, n11321, n11320, n11319, n11318, 
        n11317, n11316, n11315, n11313, n6622, n11312, n11311, 
        n11310, n11309, n11308, n11307, n11306, n11305, n11304, 
        n11303, n11302, n11301, n11300, n11299, n11298, n11297, 
        n11296, n11292;
    wire [35:0]n6775;
    
    wire n11291, n11290, n11289, n11288, n11287, n11286, n11285, 
        n11284, n11283, n11282, n11281, n11280, n11279, n11278, 
        n11277, n11276, n11275, n11274;
    wire [35:0]n6813;
    
    wire n11273, n11272, n11271, n11270, n11269, n11268, n11267, 
        n11266, n11265, n11264, n11263, n11262, n11261, n11260, 
        n11259, n11258, n11257, n11900;
    wire [35:0]n4799;
    
    wire n11666;
    wire [35:0]n5863;
    
    wire n11665, n11664, n11663, n11662, n11661, n11660, n11659, 
        n11658, n11657, n11656, n11655, n11654, n11653, n11652, 
        n11651, n11650, n11150, n6774, n11149, n11148, n11147, 
        n11146, n11145, n11144, n11143, n11142, n11141, n11140, 
        n11139, n11138, n11137, n11136, n11135, n11134, n11133, 
        n11132, n11131, n11130, n11129, n11128, n11127, n11126, 
        n11125, n11124, n11123, n11122, n11121, n11120, n11119, 
        n11118, n11117, n11116, n11115, n11073, n11072, n11071, 
        n11070, n11069, n11068, n11067, n11066, n11065, n11064, 
        n11063, n11062, n11061, n11060, n11059, n11058, n11057, 
        n11056, n11055, n6014, n11054, n11053, n11052, n11051, 
        n11050, n11049, n11048, n11047, n11046, n11045, n11044, 
        n11043, n11042, n11041, n11040, n11039, n11038, n11037, 
        n5862, n11036, n11035, n11034, n11033, n11032, n11031, 
        n11030, n11029, n11028, n11027, n11026, n11025, n11024, 
        n11023, n11022, n11021, n11020, n10988, n10987, n10986, 
        n10985, n10984, n10983, n10982, n10981, n10962, n10961, 
        n10960, n10959, n10958, n10957, n10956, n10955, n10954, 
        n10953, n10952, n10951, n10950, n10949, n10948, n10947, 
        n10946, n10945, n10943, n10942, n10941, n10940, n10939, 
        n10938, n10937, n10936, n10935, n10934, n10933, n10932, 
        n10931, n10930, n10929, n10928, n10927, n10926, n10924, 
        n10923, n10922, n10921, n10920, n10919, n10918, n10917, 
        n10916, n10915, n10914, n10913, n10912, n10911, n10910, 
        n10909, n10908, n10907, n10905, n10904, n10903, n10902, 
        n10901, n10900, n10899, n10898, n10897, n10896, n10895, 
        n10894, n10893, n10892, n10891, n10890, n10889, n10888, 
        n10878, n4798, n10877, n10876, n10875, n10874, n10873, 
        n10872, n10871, n10870, n10869, n10868, n10867, n10866, 
        n10865, n10864, n10863, n10862, n10861, n11649, n11647, 
        n11646, n11645, n11644, n11643, n11642, n11641, n11640, 
        n11639, n11638, n11637, n11636, n11635, n11634, n11633, 
        n11632, n11631, n11630, n11488;
    wire [35:0]n6015;
    
    wire n11487, n11486, n11485, n11484, n11483, n11482, n11481, 
        n11480, n11479, n11478, n11477, n11476, n11475, n11474, 
        n11473, n11472, n11471, n11469, n11468, n11467, n11466, 
        n11465, n11464, n11463, n11462, n11461, n11460, n11459, 
        n11458, n11457, n11456, n11455, n11454, n11453, n11452, 
        n11448, n11447, n11446, n11445, n11444, n11443, n11442, 
        n11441, n11440, n11439, n11438, n11437, n13828, n13829, 
        n13826, n13825, n21, n19, n15, n11895, n11899, n11898, 
        n11847, n11848, n11849, n11852, n11867, n11868, n11865, 
        n11866, n11863, n11864, n11861, n11862, n11859, n11860, 
        n11857, n11858, n11855, n11856, n11854, n11897, n11917, 
        n11918, n11950, n11949, n11948, n11947, n11916, n11946, 
        n11915, n11945, n11944, n11943, n11914, n11942, n11941, 
        n11940, n11939, n11938, n11937, n11936, n11935, n11934, 
        n11896, n11931, n11930, n11929, n11928, n11927, n11926, 
        n11925, n11924, n11853, n11909, n11923, n11908, n11922, 
        n11907, n11921, n11906, n11920, n11905, n11919;
    
    CCU2D add_1019_29 (.A0(d3[62]), .B0(n5102), .C0(n5103[26]), .D0(d2[62]), 
          .A1(d3[63]), .B1(n5102), .C1(n5103[27]), .D1(d2[63]), .CIN(n11845), 
          .COUT(n11846), .S0(d3_71__N_561[62]), .S1(d3_71__N_561[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1019_29.INIT0 = 16'h74b8;
    defparam add_1019_29.INIT1 = 16'h74b8;
    defparam add_1019_29.INJECT1_0 = "NO";
    defparam add_1019_29.INJECT1_1 = "NO";
    CCU2D add_1019_23 (.A0(d3[56]), .B0(n5102), .C0(n5103[20]), .D0(d2[56]), 
          .A1(d3[57]), .B1(n5102), .C1(n5103[21]), .D1(d2[57]), .CIN(n11842), 
          .COUT(n11843), .S0(d3_71__N_561[56]), .S1(d3_71__N_561[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1019_23.INIT0 = 16'h74b8;
    defparam add_1019_23.INIT1 = 16'h74b8;
    defparam add_1019_23.INJECT1_0 = "NO";
    defparam add_1019_23.INJECT1_1 = "NO";
    CCU2D add_1019_17 (.A0(d3[50]), .B0(n5102), .C0(n5103[14]), .D0(d2[50]), 
          .A1(d3[51]), .B1(n5102), .C1(n5103[15]), .D1(d2[51]), .CIN(n11839), 
          .COUT(n11840), .S0(d3_71__N_561[50]), .S1(d3_71__N_561[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1019_17.INIT0 = 16'h74b8;
    defparam add_1019_17.INIT1 = 16'h74b8;
    defparam add_1019_17.INJECT1_0 = "NO";
    defparam add_1019_17.INJECT1_1 = "NO";
    CCU2D add_1019_21 (.A0(d3[54]), .B0(n5102), .C0(n5103[18]), .D0(d2[54]), 
          .A1(d3[55]), .B1(n5102), .C1(n5103[19]), .D1(d2[55]), .CIN(n11841), 
          .COUT(n11842), .S0(d3_71__N_561[54]), .S1(d3_71__N_561[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1019_21.INIT0 = 16'h74b8;
    defparam add_1019_21.INIT1 = 16'h74b8;
    defparam add_1019_21.INJECT1_0 = "NO";
    defparam add_1019_21.INJECT1_1 = "NO";
    CCU2D add_1019_27 (.A0(d3[60]), .B0(n5102), .C0(n5103[24]), .D0(d2[60]), 
          .A1(d3[61]), .B1(n5102), .C1(n5103[25]), .D1(d2[61]), .CIN(n11844), 
          .COUT(n11845), .S0(d3_71__N_561[60]), .S1(d3_71__N_561[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1019_27.INIT0 = 16'h74b8;
    defparam add_1019_27.INIT1 = 16'h74b8;
    defparam add_1019_27.INJECT1_0 = "NO";
    defparam add_1019_27.INJECT1_1 = "NO";
    CCU2D add_1019_19 (.A0(d3[52]), .B0(n5102), .C0(n5103[16]), .D0(d2[52]), 
          .A1(d3[53]), .B1(n5102), .C1(n5103[17]), .D1(d2[53]), .CIN(n11840), 
          .COUT(n11841), .S0(d3_71__N_561[52]), .S1(d3_71__N_561[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1019_19.INIT0 = 16'h74b8;
    defparam add_1019_19.INIT1 = 16'h74b8;
    defparam add_1019_19.INJECT1_0 = "NO";
    defparam add_1019_19.INJECT1_1 = "NO";
    CCU2D add_1013_4 (.A0(d1[38]), .B0(d2[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[39]), .B1(d2[39]), .C1(GND_net), .D1(GND_net), .CIN(n11893), 
          .COUT(n11894), .S0(n4951[2]), .S1(n4951[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1013_4.INIT0 = 16'h5666;
    defparam add_1013_4.INIT1 = 16'h5666;
    defparam add_1013_4.INJECT1_0 = "NO";
    defparam add_1013_4.INJECT1_1 = "NO";
    FD1P3AX d_tmp_i0_i0 (.D(d5[0]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i0 (.D(d_tmp[0]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i0.GSR = "ENABLED";
    FD1S3AX d2_i0 (.D(d2_71__N_489[0]), .CK(osc_clk), .Q(d2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i0.GSR = "ENABLED";
    FD1S3AX d3_i0 (.D(d3_71__N_561[0]), .CK(osc_clk), .Q(d3[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i0.GSR = "ENABLED";
    FD1S3AX d4_i0 (.D(d4_71__N_633[0]), .CK(osc_clk), .Q(d4[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i0.GSR = "ENABLED";
    FD1S3AX d5_i0 (.D(d5_71__N_705[0]), .CK(osc_clk), .Q(d5[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i0.GSR = "ENABLED";
    FD1P3AX d6_i0_i0 (.D(d6_71__N_1458[0]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i0 (.D(d6[0]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i0.GSR = "ENABLED";
    FD1S3AX v_comb_66 (.D(osc_clk_enable_743), .CK(osc_clk), .Q(v_comb)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66.GSR = "ENABLED";
    FD1P3AX d7_i0_i0 (.D(d7_71__N_1530[0]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i0 (.D(d7[0]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d8_i0_i0 (.D(d8_71__N_1602[0]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i0 (.D(d8[0]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d9_i0_i0 (.D(d9_71__N_1674[0]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i0 (.D(d9[0]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_out_i0_i0 (.D(d_out_11__N_1818[0]), .SP(osc_clk_enable_783), 
            .CK(osc_clk), .Q(CIC1_outCos[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i0.GSR = "ENABLED";
    FD1S3AX d1_i0 (.D(d1_71__N_417[0]), .CK(osc_clk), .Q(d1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i0.GSR = "ENABLED";
    CCU2D add_1013_2 (.A0(d1[36]), .B0(d2[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[37]), .B1(d2[37]), .C1(GND_net), .D1(GND_net), .COUT(n11893), 
          .S1(n4951[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1013_2.INIT0 = 16'h7000;
    defparam add_1013_2.INIT1 = 16'h5666;
    defparam add_1013_2.INJECT1_0 = "NO";
    defparam add_1013_2.INJECT1_1 = "NO";
    CCU2D add_1014_33 (.A0(d2[66]), .B0(n4950), .C0(n4951[30]), .D0(d1[66]), 
          .A1(d2[67]), .B1(n4950), .C1(n4951[31]), .D1(d1[67]), .CIN(n11888), 
          .COUT(n11889), .S0(d2_71__N_489[66]), .S1(d2_71__N_489[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1014_33.INIT0 = 16'h74b8;
    defparam add_1014_33.INIT1 = 16'h74b8;
    defparam add_1014_33.INJECT1_0 = "NO";
    defparam add_1014_33.INJECT1_1 = "NO";
    CCU2D add_1014_29 (.A0(d2[62]), .B0(n4950), .C0(n4951[26]), .D0(d1[62]), 
          .A1(d2[63]), .B1(n4950), .C1(n4951[27]), .D1(d1[63]), .CIN(n11886), 
          .COUT(n11887), .S0(d2_71__N_489[62]), .S1(d2_71__N_489[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1014_29.INIT0 = 16'h74b8;
    defparam add_1014_29.INIT1 = 16'h74b8;
    defparam add_1014_29.INJECT1_0 = "NO";
    defparam add_1014_29.INJECT1_1 = "NO";
    CCU2D add_1014_27 (.A0(d2[60]), .B0(n4950), .C0(n4951[24]), .D0(d1[60]), 
          .A1(d2[61]), .B1(n4950), .C1(n4951[25]), .D1(d1[61]), .CIN(n11885), 
          .COUT(n11886), .S0(d2_71__N_489[60]), .S1(d2_71__N_489[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1014_27.INIT0 = 16'h74b8;
    defparam add_1014_27.INIT1 = 16'h74b8;
    defparam add_1014_27.INJECT1_0 = "NO";
    defparam add_1014_27.INJECT1_1 = "NO";
    CCU2D add_1014_25 (.A0(d2[58]), .B0(n4950), .C0(n4951[22]), .D0(d1[58]), 
          .A1(d2[59]), .B1(n4950), .C1(n4951[23]), .D1(d1[59]), .CIN(n11884), 
          .COUT(n11885), .S0(d2_71__N_489[58]), .S1(d2_71__N_489[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1014_25.INIT0 = 16'h74b8;
    defparam add_1014_25.INIT1 = 16'h74b8;
    defparam add_1014_25.INJECT1_0 = "NO";
    defparam add_1014_25.INJECT1_1 = "NO";
    CCU2D add_1014_23 (.A0(d2[56]), .B0(n4950), .C0(n4951[20]), .D0(d1[56]), 
          .A1(d2[57]), .B1(n4950), .C1(n4951[21]), .D1(d1[57]), .CIN(n11883), 
          .COUT(n11884), .S0(d2_71__N_489[56]), .S1(d2_71__N_489[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1014_23.INIT0 = 16'h74b8;
    defparam add_1014_23.INIT1 = 16'h74b8;
    defparam add_1014_23.INJECT1_0 = "NO";
    defparam add_1014_23.INJECT1_1 = "NO";
    CCU2D add_1019_25 (.A0(d3[58]), .B0(n5102), .C0(n5103[22]), .D0(d2[58]), 
          .A1(d3[59]), .B1(n5102), .C1(n5103[23]), .D1(d2[59]), .CIN(n11843), 
          .COUT(n11844), .S0(d3_71__N_561[58]), .S1(d3_71__N_561[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1019_25.INIT0 = 16'h74b8;
    defparam add_1019_25.INIT1 = 16'h74b8;
    defparam add_1019_25.INJECT1_0 = "NO";
    defparam add_1019_25.INJECT1_1 = "NO";
    CCU2D add_1014_21 (.A0(d2[54]), .B0(n4950), .C0(n4951[18]), .D0(d1[54]), 
          .A1(d2[55]), .B1(n4950), .C1(n4951[19]), .D1(d1[55]), .CIN(n11882), 
          .COUT(n11883), .S0(d2_71__N_489[54]), .S1(d2_71__N_489[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1014_21.INIT0 = 16'h74b8;
    defparam add_1014_21.INIT1 = 16'h74b8;
    defparam add_1014_21.INJECT1_0 = "NO";
    defparam add_1014_21.INJECT1_1 = "NO";
    CCU2D add_1014_19 (.A0(d2[52]), .B0(n4950), .C0(n4951[16]), .D0(d1[52]), 
          .A1(d2[53]), .B1(n4950), .C1(n4951[17]), .D1(d1[53]), .CIN(n11881), 
          .COUT(n11882), .S0(d2_71__N_489[52]), .S1(d2_71__N_489[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1014_19.INIT0 = 16'h74b8;
    defparam add_1014_19.INIT1 = 16'h74b8;
    defparam add_1014_19.INJECT1_0 = "NO";
    defparam add_1014_19.INJECT1_1 = "NO";
    CCU2D add_1014_17 (.A0(d2[50]), .B0(n4950), .C0(n4951[14]), .D0(d1[50]), 
          .A1(d2[51]), .B1(n4950), .C1(n4951[15]), .D1(d1[51]), .CIN(n11880), 
          .COUT(n11881), .S0(d2_71__N_489[50]), .S1(d2_71__N_489[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1014_17.INIT0 = 16'h74b8;
    defparam add_1014_17.INIT1 = 16'h74b8;
    defparam add_1014_17.INJECT1_0 = "NO";
    defparam add_1014_17.INJECT1_1 = "NO";
    CCU2D add_1019_13 (.A0(d3[46]), .B0(n5102), .C0(n5103[10]), .D0(d2[46]), 
          .A1(d3[47]), .B1(n5102), .C1(n5103[11]), .D1(d2[47]), .CIN(n11837), 
          .COUT(n11838), .S0(d3_71__N_561[46]), .S1(d3_71__N_561[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1019_13.INIT0 = 16'h74b8;
    defparam add_1019_13.INIT1 = 16'h74b8;
    defparam add_1019_13.INJECT1_0 = "NO";
    defparam add_1019_13.INJECT1_1 = "NO";
    CCU2D add_1014_37 (.A0(d2[70]), .B0(n4950), .C0(n4951[34]), .D0(d1[70]), 
          .A1(d2[71]), .B1(n4950), .C1(n4951[35]), .D1(d1[71]), .CIN(n11890), 
          .S0(d2_71__N_489[70]), .S1(d2_71__N_489[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1014_37.INIT0 = 16'h74b8;
    defparam add_1014_37.INIT1 = 16'h74b8;
    defparam add_1014_37.INJECT1_0 = "NO";
    defparam add_1014_37.INJECT1_1 = "NO";
    CCU2D add_1014_35 (.A0(d2[68]), .B0(n4950), .C0(n4951[32]), .D0(d1[68]), 
          .A1(d2[69]), .B1(n4950), .C1(n4951[33]), .D1(d1[69]), .CIN(n11889), 
          .COUT(n11890), .S0(d2_71__N_489[68]), .S1(d2_71__N_489[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1014_35.INIT0 = 16'h74b8;
    defparam add_1014_35.INIT1 = 16'h74b8;
    defparam add_1014_35.INJECT1_0 = "NO";
    defparam add_1014_35.INJECT1_1 = "NO";
    CCU2D add_1014_31 (.A0(d2[64]), .B0(n4950), .C0(n4951[28]), .D0(d1[64]), 
          .A1(d2[65]), .B1(n4950), .C1(n4951[29]), .D1(d1[65]), .CIN(n11887), 
          .COUT(n11888), .S0(d2_71__N_489[64]), .S1(d2_71__N_489[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1014_31.INIT0 = 16'h74b8;
    defparam add_1014_31.INIT1 = 16'h74b8;
    defparam add_1014_31.INJECT1_0 = "NO";
    defparam add_1014_31.INJECT1_1 = "NO";
    CCU2D add_1019_5 (.A0(d3[38]), .B0(n5102), .C0(n5103[2]), .D0(d2[38]), 
          .A1(d3[39]), .B1(n5102), .C1(n5103[3]), .D1(d2[39]), .CIN(n11833), 
          .COUT(n11834), .S0(d3_71__N_561[38]), .S1(d3_71__N_561[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1019_5.INIT0 = 16'h74b8;
    defparam add_1019_5.INIT1 = 16'h74b8;
    defparam add_1019_5.INJECT1_0 = "NO";
    defparam add_1019_5.INJECT1_1 = "NO";
    CCU2D add_1023_32 (.A0(d3[66]), .B0(d4[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[67]), .B1(d4[67]), .C1(GND_net), .D1(GND_net), .CIN(n11825), 
          .COUT(n11826), .S0(n5255[30]), .S1(n5255[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1023_32.INIT0 = 16'h5666;
    defparam add_1023_32.INIT1 = 16'h5666;
    defparam add_1023_32.INJECT1_0 = "NO";
    defparam add_1023_32.INJECT1_1 = "NO";
    CCU2D add_1024_11 (.A0(d4[44]), .B0(n5254), .C0(n5255[8]), .D0(d3[44]), 
          .A1(d4[45]), .B1(n5254), .C1(n5255[9]), .D1(d3[45]), .CIN(n11795), 
          .COUT(n11796), .S0(d4_71__N_633[44]), .S1(d4_71__N_633[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1024_11.INIT0 = 16'h74b8;
    defparam add_1024_11.INIT1 = 16'h74b8;
    defparam add_1024_11.INJECT1_0 = "NO";
    defparam add_1024_11.INJECT1_1 = "NO";
    CCU2D add_1023_30 (.A0(d3[64]), .B0(d4[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[65]), .B1(d4[65]), .C1(GND_net), .D1(GND_net), .CIN(n11824), 
          .COUT(n11825), .S0(n5255[28]), .S1(n5255[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1023_30.INIT0 = 16'h5666;
    defparam add_1023_30.INIT1 = 16'h5666;
    defparam add_1023_30.INJECT1_0 = "NO";
    defparam add_1023_30.INJECT1_1 = "NO";
    CCU2D add_1019_3 (.A0(d3[36]), .B0(n5102), .C0(n5103[0]), .D0(d2[36]), 
          .A1(d3[37]), .B1(n5102), .C1(n5103[1]), .D1(d2[37]), .CIN(n11832), 
          .COUT(n11833), .S0(d3_71__N_561[36]), .S1(d3_71__N_561[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1019_3.INIT0 = 16'h74b8;
    defparam add_1019_3.INIT1 = 16'h74b8;
    defparam add_1019_3.INJECT1_0 = "NO";
    defparam add_1019_3.INJECT1_1 = "NO";
    CCU2D add_1053_11 (.A0(d_tmp[45]), .B0(d_d_tmp[45]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[46]), .B1(d_d_tmp[46]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11435), .COUT(n11436), .S0(n6167[9]), 
          .S1(n6167[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1053_11.INIT0 = 16'h5999;
    defparam add_1053_11.INIT1 = 16'h5999;
    defparam add_1053_11.INJECT1_0 = "NO";
    defparam add_1053_11.INJECT1_1 = "NO";
    CCU2D add_1023_28 (.A0(d3[62]), .B0(d4[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[63]), .B1(d4[63]), .C1(GND_net), .D1(GND_net), .CIN(n11823), 
          .COUT(n11824), .S0(n5255[26]), .S1(n5255[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1023_28.INIT0 = 16'h5666;
    defparam add_1023_28.INIT1 = 16'h5666;
    defparam add_1023_28.INJECT1_0 = "NO";
    defparam add_1023_28.INJECT1_1 = "NO";
    CCU2D add_1019_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5102), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11832));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1019_1.INIT0 = 16'hF000;
    defparam add_1019_1.INIT1 = 16'h0555;
    defparam add_1019_1.INJECT1_0 = "NO";
    defparam add_1019_1.INJECT1_1 = "NO";
    CCU2D add_1019_11 (.A0(d3[44]), .B0(n5102), .C0(n5103[8]), .D0(d2[44]), 
          .A1(d3[45]), .B1(n5102), .C1(n5103[9]), .D1(d2[45]), .CIN(n11836), 
          .COUT(n11837), .S0(d3_71__N_561[44]), .S1(d3_71__N_561[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1019_11.INIT0 = 16'h74b8;
    defparam add_1019_11.INIT1 = 16'h74b8;
    defparam add_1019_11.INJECT1_0 = "NO";
    defparam add_1019_11.INJECT1_1 = "NO";
    CCU2D add_1023_24 (.A0(d3[58]), .B0(d4[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[59]), .B1(d4[59]), .C1(GND_net), .D1(GND_net), .CIN(n11821), 
          .COUT(n11822), .S0(n5255[22]), .S1(n5255[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1023_24.INIT0 = 16'h5666;
    defparam add_1023_24.INIT1 = 16'h5666;
    defparam add_1023_24.INJECT1_0 = "NO";
    defparam add_1023_24.INJECT1_1 = "NO";
    CCU2D add_1023_22 (.A0(d3[56]), .B0(d4[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[57]), .B1(d4[57]), .C1(GND_net), .D1(GND_net), .CIN(n11820), 
          .COUT(n11821), .S0(n5255[20]), .S1(n5255[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1023_22.INIT0 = 16'h5666;
    defparam add_1023_22.INIT1 = 16'h5666;
    defparam add_1023_22.INJECT1_0 = "NO";
    defparam add_1023_22.INJECT1_1 = "NO";
    CCU2D add_1023_20 (.A0(d3[54]), .B0(d4[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[55]), .B1(d4[55]), .C1(GND_net), .D1(GND_net), .CIN(n11819), 
          .COUT(n11820), .S0(n5255[18]), .S1(n5255[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1023_20.INIT0 = 16'h5666;
    defparam add_1023_20.INIT1 = 16'h5666;
    defparam add_1023_20.INJECT1_0 = "NO";
    defparam add_1023_20.INJECT1_1 = "NO";
    CCU2D add_1023_18 (.A0(d3[52]), .B0(d4[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[53]), .B1(d4[53]), .C1(GND_net), .D1(GND_net), .CIN(n11818), 
          .COUT(n11819), .S0(n5255[16]), .S1(n5255[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1023_18.INIT0 = 16'h5666;
    defparam add_1023_18.INIT1 = 16'h5666;
    defparam add_1023_18.INJECT1_0 = "NO";
    defparam add_1023_18.INJECT1_1 = "NO";
    CCU2D add_1023_12 (.A0(d3[46]), .B0(d4[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[47]), .B1(d4[47]), .C1(GND_net), .D1(GND_net), .CIN(n11815), 
          .COUT(n11816), .S0(n5255[10]), .S1(n5255[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1023_12.INIT0 = 16'h5666;
    defparam add_1023_12.INIT1 = 16'h5666;
    defparam add_1023_12.INJECT1_0 = "NO";
    defparam add_1023_12.INJECT1_1 = "NO";
    CCU2D add_1023_6 (.A0(d3[40]), .B0(d4[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[41]), .B1(d4[41]), .C1(GND_net), .D1(GND_net), .CIN(n11812), 
          .COUT(n11813), .S0(n5255[4]), .S1(n5255[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1023_6.INIT0 = 16'h5666;
    defparam add_1023_6.INIT1 = 16'h5666;
    defparam add_1023_6.INJECT1_0 = "NO";
    defparam add_1023_6.INJECT1_1 = "NO";
    CCU2D add_1024_9 (.A0(d4[42]), .B0(n5254), .C0(n5255[6]), .D0(d3[42]), 
          .A1(d4[43]), .B1(n5254), .C1(n5255[7]), .D1(d3[43]), .CIN(n11794), 
          .COUT(n11795), .S0(d4_71__N_633[42]), .S1(d4_71__N_633[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1024_9.INIT0 = 16'h74b8;
    defparam add_1024_9.INIT1 = 16'h74b8;
    defparam add_1024_9.INJECT1_0 = "NO";
    defparam add_1024_9.INJECT1_1 = "NO";
    CCU2D add_1023_10 (.A0(d3[44]), .B0(d4[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[45]), .B1(d4[45]), .C1(GND_net), .D1(GND_net), .CIN(n11814), 
          .COUT(n11815), .S0(n5255[8]), .S1(n5255[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1023_10.INIT0 = 16'h5666;
    defparam add_1023_10.INIT1 = 16'h5666;
    defparam add_1023_10.INJECT1_0 = "NO";
    defparam add_1023_10.INJECT1_1 = "NO";
    CCU2D add_1023_16 (.A0(d3[50]), .B0(d4[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[51]), .B1(d4[51]), .C1(GND_net), .D1(GND_net), .CIN(n11817), 
          .COUT(n11818), .S0(n5255[14]), .S1(n5255[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1023_16.INIT0 = 16'h5666;
    defparam add_1023_16.INIT1 = 16'h5666;
    defparam add_1023_16.INJECT1_0 = "NO";
    defparam add_1023_16.INJECT1_1 = "NO";
    CCU2D add_1023_8 (.A0(d3[42]), .B0(d4[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[43]), .B1(d4[43]), .C1(GND_net), .D1(GND_net), .CIN(n11813), 
          .COUT(n11814), .S0(n5255[6]), .S1(n5255[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1023_8.INIT0 = 16'h5666;
    defparam add_1023_8.INIT1 = 16'h5666;
    defparam add_1023_8.INJECT1_0 = "NO";
    defparam add_1023_8.INJECT1_1 = "NO";
    CCU2D add_1023_4 (.A0(d3[38]), .B0(d4[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[39]), .B1(d4[39]), .C1(GND_net), .D1(GND_net), .CIN(n11811), 
          .COUT(n11812), .S0(n5255[2]), .S1(n5255[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1023_4.INIT0 = 16'h5666;
    defparam add_1023_4.INIT1 = 16'h5666;
    defparam add_1023_4.INJECT1_0 = "NO";
    defparam add_1023_4.INJECT1_1 = "NO";
    CCU2D add_1023_14 (.A0(d3[48]), .B0(d4[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[49]), .B1(d4[49]), .C1(GND_net), .D1(GND_net), .CIN(n11816), 
          .COUT(n11817), .S0(n5255[12]), .S1(n5255[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1023_14.INIT0 = 16'h5666;
    defparam add_1023_14.INIT1 = 16'h5666;
    defparam add_1023_14.INJECT1_0 = "NO";
    defparam add_1023_14.INJECT1_1 = "NO";
    CCU2D add_1024_7 (.A0(d4[40]), .B0(n5254), .C0(n5255[4]), .D0(d3[40]), 
          .A1(d4[41]), .B1(n5254), .C1(n5255[5]), .D1(d3[41]), .CIN(n11793), 
          .COUT(n11794), .S0(d4_71__N_633[40]), .S1(d4_71__N_633[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1024_7.INIT0 = 16'h74b8;
    defparam add_1024_7.INIT1 = 16'h74b8;
    defparam add_1024_7.INJECT1_0 = "NO";
    defparam add_1024_7.INJECT1_1 = "NO";
    CCU2D add_1023_26 (.A0(d3[60]), .B0(d4[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[61]), .B1(d4[61]), .C1(GND_net), .D1(GND_net), .CIN(n11822), 
          .COUT(n11823), .S0(n5255[24]), .S1(n5255[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1023_26.INIT0 = 16'h5666;
    defparam add_1023_26.INIT1 = 16'h5666;
    defparam add_1023_26.INJECT1_0 = "NO";
    defparam add_1023_26.INJECT1_1 = "NO";
    CCU2D add_1023_36 (.A0(d3[70]), .B0(d4[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[71]), .B1(d4[71]), .C1(GND_net), .D1(GND_net), .CIN(n11827), 
          .S0(n5255[34]), .S1(n5255[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1023_36.INIT0 = 16'h5666;
    defparam add_1023_36.INIT1 = 16'h5666;
    defparam add_1023_36.INJECT1_0 = "NO";
    defparam add_1023_36.INJECT1_1 = "NO";
    CCU2D add_1024_5 (.A0(d4[38]), .B0(n5254), .C0(n5255[2]), .D0(d3[38]), 
          .A1(d4[39]), .B1(n5254), .C1(n5255[3]), .D1(d3[39]), .CIN(n11792), 
          .COUT(n11793), .S0(d4_71__N_633[38]), .S1(d4_71__N_633[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1024_5.INIT0 = 16'h74b8;
    defparam add_1024_5.INIT1 = 16'h74b8;
    defparam add_1024_5.INJECT1_0 = "NO";
    defparam add_1024_5.INJECT1_1 = "NO";
    CCU2D add_1019_9 (.A0(d3[42]), .B0(n5102), .C0(n5103[6]), .D0(d2[42]), 
          .A1(d3[43]), .B1(n5102), .C1(n5103[7]), .D1(d2[43]), .CIN(n11835), 
          .COUT(n11836), .S0(d3_71__N_561[42]), .S1(d3_71__N_561[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1019_9.INIT0 = 16'h74b8;
    defparam add_1019_9.INIT1 = 16'h74b8;
    defparam add_1019_9.INJECT1_0 = "NO";
    defparam add_1019_9.INJECT1_1 = "NO";
    CCU2D add_1053_9 (.A0(d_tmp[43]), .B0(d_d_tmp[43]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[44]), .B1(d_d_tmp[44]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11434), .COUT(n11435), .S0(n6167[7]), 
          .S1(n6167[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1053_9.INIT0 = 16'h5999;
    defparam add_1053_9.INIT1 = 16'h5999;
    defparam add_1053_9.INJECT1_0 = "NO";
    defparam add_1053_9.INJECT1_1 = "NO";
    CCU2D add_1053_7 (.A0(d_tmp[41]), .B0(d_d_tmp[41]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[42]), .B1(d_d_tmp[42]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11433), .COUT(n11434), .S0(n6167[5]), 
          .S1(n6167[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1053_7.INIT0 = 16'h5999;
    defparam add_1053_7.INIT1 = 16'h5999;
    defparam add_1053_7.INJECT1_0 = "NO";
    defparam add_1053_7.INJECT1_1 = "NO";
    CCU2D add_1023_34 (.A0(d3[68]), .B0(d4[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[69]), .B1(d4[69]), .C1(GND_net), .D1(GND_net), .CIN(n11826), 
          .COUT(n11827), .S0(n5255[32]), .S1(n5255[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1023_34.INIT0 = 16'h5666;
    defparam add_1023_34.INIT1 = 16'h5666;
    defparam add_1023_34.INJECT1_0 = "NO";
    defparam add_1023_34.INJECT1_1 = "NO";
    CCU2D add_1019_7 (.A0(d3[40]), .B0(n5102), .C0(n5103[4]), .D0(d2[40]), 
          .A1(d3[41]), .B1(n5102), .C1(n5103[5]), .D1(d2[41]), .CIN(n11834), 
          .COUT(n11835), .S0(d3_71__N_561[40]), .S1(d3_71__N_561[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1019_7.INIT0 = 16'h74b8;
    defparam add_1019_7.INIT1 = 16'h74b8;
    defparam add_1019_7.INJECT1_0 = "NO";
    defparam add_1019_7.INJECT1_1 = "NO";
    CCU2D add_1053_5 (.A0(d_tmp[39]), .B0(d_d_tmp[39]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[40]), .B1(d_d_tmp[40]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11432), .COUT(n11433), .S0(n6167[3]), 
          .S1(n6167[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1053_5.INIT0 = 16'h5999;
    defparam add_1053_5.INIT1 = 16'h5999;
    defparam add_1053_5.INJECT1_0 = "NO";
    defparam add_1053_5.INJECT1_1 = "NO";
    CCU2D add_1053_3 (.A0(d_tmp[37]), .B0(d_d_tmp[37]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[38]), .B1(d_d_tmp[38]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11431), .COUT(n11432), .S0(n6167[1]), 
          .S1(n6167[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1053_3.INIT0 = 16'h5999;
    defparam add_1053_3.INIT1 = 16'h5999;
    defparam add_1053_3.INJECT1_0 = "NO";
    defparam add_1053_3.INJECT1_1 = "NO";
    CCU2D add_1023_2 (.A0(d3[36]), .B0(d4[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[37]), .B1(d4[37]), .C1(GND_net), .D1(GND_net), .COUT(n11811), 
          .S1(n5255[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1023_2.INIT0 = 16'h7000;
    defparam add_1023_2.INIT1 = 16'h5666;
    defparam add_1023_2.INJECT1_0 = "NO";
    defparam add_1023_2.INJECT1_1 = "NO";
    CCU2D add_1024_3 (.A0(d4[36]), .B0(n5254), .C0(n5255[0]), .D0(d3[36]), 
          .A1(d4[37]), .B1(n5254), .C1(n5255[1]), .D1(d3[37]), .CIN(n11791), 
          .COUT(n11792), .S0(d4_71__N_633[36]), .S1(d4_71__N_633[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1024_3.INIT0 = 16'h74b8;
    defparam add_1024_3.INIT1 = 16'h74b8;
    defparam add_1024_3.INJECT1_0 = "NO";
    defparam add_1024_3.INJECT1_1 = "NO";
    CCU2D add_1024_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5254), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11791));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1024_1.INIT0 = 16'hF000;
    defparam add_1024_1.INIT1 = 16'h0555;
    defparam add_1024_1.INJECT1_0 = "NO";
    defparam add_1024_1.INJECT1_1 = "NO";
    CCU2D add_1028_36 (.A0(d4[70]), .B0(d5[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[71]), .B1(d5[71]), .C1(GND_net), .D1(GND_net), .CIN(n11786), 
          .S0(n5407[34]), .S1(n5407[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1028_36.INIT0 = 16'h5666;
    defparam add_1028_36.INIT1 = 16'h5666;
    defparam add_1028_36.INJECT1_0 = "NO";
    defparam add_1028_36.INJECT1_1 = "NO";
    CCU2D add_1028_34 (.A0(d4[68]), .B0(d5[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[69]), .B1(d5[69]), .C1(GND_net), .D1(GND_net), .CIN(n11785), 
          .COUT(n11786), .S0(n5407[32]), .S1(n5407[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1028_34.INIT0 = 16'h5666;
    defparam add_1028_34.INIT1 = 16'h5666;
    defparam add_1028_34.INJECT1_0 = "NO";
    defparam add_1028_34.INJECT1_1 = "NO";
    CCU2D add_1024_31 (.A0(d4[64]), .B0(n5254), .C0(n5255[28]), .D0(d3[64]), 
          .A1(d4[65]), .B1(n5254), .C1(n5255[29]), .D1(d3[65]), .CIN(n11805), 
          .COUT(n11806), .S0(d4_71__N_633[64]), .S1(d4_71__N_633[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1024_31.INIT0 = 16'h74b8;
    defparam add_1024_31.INIT1 = 16'h74b8;
    defparam add_1024_31.INJECT1_0 = "NO";
    defparam add_1024_31.INJECT1_1 = "NO";
    CCU2D add_1024_19 (.A0(d4[52]), .B0(n5254), .C0(n5255[16]), .D0(d3[52]), 
          .A1(d4[53]), .B1(n5254), .C1(n5255[17]), .D1(d3[53]), .CIN(n11799), 
          .COUT(n11800), .S0(d4_71__N_633[52]), .S1(d4_71__N_633[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1024_19.INIT0 = 16'h74b8;
    defparam add_1024_19.INIT1 = 16'h74b8;
    defparam add_1024_19.INJECT1_0 = "NO";
    defparam add_1024_19.INJECT1_1 = "NO";
    CCU2D add_1028_32 (.A0(d4[66]), .B0(d5[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[67]), .B1(d5[67]), .C1(GND_net), .D1(GND_net), .CIN(n11784), 
          .COUT(n11785), .S0(n5407[30]), .S1(n5407[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1028_32.INIT0 = 16'h5666;
    defparam add_1028_32.INIT1 = 16'h5666;
    defparam add_1028_32.INJECT1_0 = "NO";
    defparam add_1028_32.INJECT1_1 = "NO";
    CCU2D add_1024_17 (.A0(d4[50]), .B0(n5254), .C0(n5255[14]), .D0(d3[50]), 
          .A1(d4[51]), .B1(n5254), .C1(n5255[15]), .D1(d3[51]), .CIN(n11798), 
          .COUT(n11799), .S0(d4_71__N_633[50]), .S1(d4_71__N_633[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1024_17.INIT0 = 16'h74b8;
    defparam add_1024_17.INIT1 = 16'h74b8;
    defparam add_1024_17.INJECT1_0 = "NO";
    defparam add_1024_17.INJECT1_1 = "NO";
    CCU2D add_1024_29 (.A0(d4[62]), .B0(n5254), .C0(n5255[26]), .D0(d3[62]), 
          .A1(d4[63]), .B1(n5254), .C1(n5255[27]), .D1(d3[63]), .CIN(n11804), 
          .COUT(n11805), .S0(d4_71__N_633[62]), .S1(d4_71__N_633[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1024_29.INIT0 = 16'h74b8;
    defparam add_1024_29.INIT1 = 16'h74b8;
    defparam add_1024_29.INJECT1_0 = "NO";
    defparam add_1024_29.INJECT1_1 = "NO";
    CCU2D add_1024_15 (.A0(d4[48]), .B0(n5254), .C0(n5255[12]), .D0(d3[48]), 
          .A1(d4[49]), .B1(n5254), .C1(n5255[13]), .D1(d3[49]), .CIN(n11797), 
          .COUT(n11798), .S0(d4_71__N_633[48]), .S1(d4_71__N_633[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1024_15.INIT0 = 16'h74b8;
    defparam add_1024_15.INIT1 = 16'h74b8;
    defparam add_1024_15.INJECT1_0 = "NO";
    defparam add_1024_15.INJECT1_1 = "NO";
    CCU2D add_1024_27 (.A0(d4[60]), .B0(n5254), .C0(n5255[24]), .D0(d3[60]), 
          .A1(d4[61]), .B1(n5254), .C1(n5255[25]), .D1(d3[61]), .CIN(n11803), 
          .COUT(n11804), .S0(d4_71__N_633[60]), .S1(d4_71__N_633[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1024_27.INIT0 = 16'h74b8;
    defparam add_1024_27.INIT1 = 16'h74b8;
    defparam add_1024_27.INJECT1_0 = "NO";
    defparam add_1024_27.INJECT1_1 = "NO";
    CCU2D add_1024_37 (.A0(d4[70]), .B0(n5254), .C0(n5255[34]), .D0(d3[70]), 
          .A1(d4[71]), .B1(n5254), .C1(n5255[35]), .D1(d3[71]), .CIN(n11808), 
          .S0(d4_71__N_633[70]), .S1(d4_71__N_633[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1024_37.INIT0 = 16'h74b8;
    defparam add_1024_37.INIT1 = 16'h74b8;
    defparam add_1024_37.INJECT1_0 = "NO";
    defparam add_1024_37.INJECT1_1 = "NO";
    CCU2D add_1024_25 (.A0(d4[58]), .B0(n5254), .C0(n5255[22]), .D0(d3[58]), 
          .A1(d4[59]), .B1(n5254), .C1(n5255[23]), .D1(d3[59]), .CIN(n11802), 
          .COUT(n11803), .S0(d4_71__N_633[58]), .S1(d4_71__N_633[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1024_25.INIT0 = 16'h74b8;
    defparam add_1024_25.INIT1 = 16'h74b8;
    defparam add_1024_25.INJECT1_0 = "NO";
    defparam add_1024_25.INJECT1_1 = "NO";
    CCU2D add_1024_13 (.A0(d4[46]), .B0(n5254), .C0(n5255[10]), .D0(d3[46]), 
          .A1(d4[47]), .B1(n5254), .C1(n5255[11]), .D1(d3[47]), .CIN(n11796), 
          .COUT(n11797), .S0(d4_71__N_633[46]), .S1(d4_71__N_633[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1024_13.INIT0 = 16'h74b8;
    defparam add_1024_13.INIT1 = 16'h74b8;
    defparam add_1024_13.INJECT1_0 = "NO";
    defparam add_1024_13.INJECT1_1 = "NO";
    CCU2D add_1024_23 (.A0(d4[56]), .B0(n5254), .C0(n5255[20]), .D0(d3[56]), 
          .A1(d4[57]), .B1(n5254), .C1(n5255[21]), .D1(d3[57]), .CIN(n11801), 
          .COUT(n11802), .S0(d4_71__N_633[56]), .S1(d4_71__N_633[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1024_23.INIT0 = 16'h74b8;
    defparam add_1024_23.INIT1 = 16'h74b8;
    defparam add_1024_23.INJECT1_0 = "NO";
    defparam add_1024_23.INJECT1_1 = "NO";
    CCU2D add_1024_35 (.A0(d4[68]), .B0(n5254), .C0(n5255[32]), .D0(d3[68]), 
          .A1(d4[69]), .B1(n5254), .C1(n5255[33]), .D1(d3[69]), .CIN(n11807), 
          .COUT(n11808), .S0(d4_71__N_633[68]), .S1(d4_71__N_633[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1024_35.INIT0 = 16'h74b8;
    defparam add_1024_35.INIT1 = 16'h74b8;
    defparam add_1024_35.INJECT1_0 = "NO";
    defparam add_1024_35.INJECT1_1 = "NO";
    CCU2D add_1024_21 (.A0(d4[54]), .B0(n5254), .C0(n5255[18]), .D0(d3[54]), 
          .A1(d4[55]), .B1(n5254), .C1(n5255[19]), .D1(d3[55]), .CIN(n11800), 
          .COUT(n11801), .S0(d4_71__N_633[54]), .S1(d4_71__N_633[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1024_21.INIT0 = 16'h74b8;
    defparam add_1024_21.INIT1 = 16'h74b8;
    defparam add_1024_21.INJECT1_0 = "NO";
    defparam add_1024_21.INJECT1_1 = "NO";
    CCU2D add_1024_33 (.A0(d4[66]), .B0(n5254), .C0(n5255[30]), .D0(d3[66]), 
          .A1(d4[67]), .B1(n5254), .C1(n5255[31]), .D1(d3[67]), .CIN(n11806), 
          .COUT(n11807), .S0(d4_71__N_633[66]), .S1(d4_71__N_633[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1024_33.INIT0 = 16'h74b8;
    defparam add_1024_33.INIT1 = 16'h74b8;
    defparam add_1024_33.INJECT1_0 = "NO";
    defparam add_1024_33.INJECT1_1 = "NO";
    CCU2D add_1014_15 (.A0(d2[48]), .B0(n4950), .C0(n4951[12]), .D0(d1[48]), 
          .A1(d2[49]), .B1(n4950), .C1(n4951[13]), .D1(d1[49]), .CIN(n11879), 
          .COUT(n11880), .S0(d2_71__N_489[48]), .S1(d2_71__N_489[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1014_15.INIT0 = 16'h74b8;
    defparam add_1014_15.INIT1 = 16'h74b8;
    defparam add_1014_15.INJECT1_0 = "NO";
    defparam add_1014_15.INJECT1_1 = "NO";
    CCU2D add_1014_13 (.A0(d2[46]), .B0(n4950), .C0(n4951[10]), .D0(d1[46]), 
          .A1(d2[47]), .B1(n4950), .C1(n4951[11]), .D1(d1[47]), .CIN(n11878), 
          .COUT(n11879), .S0(d2_71__N_489[46]), .S1(d2_71__N_489[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1014_13.INIT0 = 16'h74b8;
    defparam add_1014_13.INIT1 = 16'h74b8;
    defparam add_1014_13.INJECT1_0 = "NO";
    defparam add_1014_13.INJECT1_1 = "NO";
    CCU2D add_1028_30 (.A0(d4[64]), .B0(d5[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[65]), .B1(d5[65]), .C1(GND_net), .D1(GND_net), .CIN(n11783), 
          .COUT(n11784), .S0(n5407[28]), .S1(n5407[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1028_30.INIT0 = 16'h5666;
    defparam add_1028_30.INIT1 = 16'h5666;
    defparam add_1028_30.INJECT1_0 = "NO";
    defparam add_1028_30.INJECT1_1 = "NO";
    CCU2D add_1014_11 (.A0(d2[44]), .B0(n4950), .C0(n4951[8]), .D0(d1[44]), 
          .A1(d2[45]), .B1(n4950), .C1(n4951[9]), .D1(d1[45]), .CIN(n11877), 
          .COUT(n11878), .S0(d2_71__N_489[44]), .S1(d2_71__N_489[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1014_11.INIT0 = 16'h74b8;
    defparam add_1014_11.INIT1 = 16'h74b8;
    defparam add_1014_11.INJECT1_0 = "NO";
    defparam add_1014_11.INJECT1_1 = "NO";
    CCU2D add_1019_15 (.A0(d3[48]), .B0(n5102), .C0(n5103[12]), .D0(d2[48]), 
          .A1(d3[49]), .B1(n5102), .C1(n5103[13]), .D1(d2[49]), .CIN(n11838), 
          .COUT(n11839), .S0(d3_71__N_561[48]), .S1(d3_71__N_561[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1019_15.INIT0 = 16'h74b8;
    defparam add_1019_15.INIT1 = 16'h74b8;
    defparam add_1019_15.INJECT1_0 = "NO";
    defparam add_1019_15.INJECT1_1 = "NO";
    CCU2D add_1014_7 (.A0(d2[40]), .B0(n4950), .C0(n4951[4]), .D0(d1[40]), 
          .A1(d2[41]), .B1(n4950), .C1(n4951[5]), .D1(d1[41]), .CIN(n11875), 
          .COUT(n11876), .S0(d2_71__N_489[40]), .S1(d2_71__N_489[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1014_7.INIT0 = 16'h74b8;
    defparam add_1014_7.INIT1 = 16'h74b8;
    defparam add_1014_7.INJECT1_0 = "NO";
    defparam add_1014_7.INJECT1_1 = "NO";
    CCU2D add_1014_3 (.A0(d2[36]), .B0(n4950), .C0(n4951[0]), .D0(d1[36]), 
          .A1(d2[37]), .B1(n4950), .C1(n4951[1]), .D1(d1[37]), .CIN(n11873), 
          .COUT(n11874), .S0(d2_71__N_489[36]), .S1(d2_71__N_489[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1014_3.INIT0 = 16'h74b8;
    defparam add_1014_3.INIT1 = 16'h74b8;
    defparam add_1014_3.INJECT1_0 = "NO";
    defparam add_1014_3.INJECT1_1 = "NO";
    CCU2D add_1053_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[36]), .B1(d_d_tmp[36]), .C1(GND_net), .D1(GND_net), 
          .COUT(n11431), .S1(n6167[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1053_1.INIT0 = 16'hF000;
    defparam add_1053_1.INIT1 = 16'h5999;
    defparam add_1053_1.INJECT1_0 = "NO";
    defparam add_1053_1.INJECT1_1 = "NO";
    CCU2D add_1054_37 (.A0(d_d_tmp[70]), .B0(n6166), .C0(n6167[34]), .D0(d_tmp[70]), 
          .A1(d_d_tmp[71]), .B1(n6166), .C1(n6167[35]), .D1(d_tmp[71]), 
          .CIN(n11429), .S0(d6_71__N_1458[70]), .S1(d6_71__N_1458[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1054_37.INIT0 = 16'hb874;
    defparam add_1054_37.INIT1 = 16'hb874;
    defparam add_1054_37.INJECT1_0 = "NO";
    defparam add_1054_37.INJECT1_1 = "NO";
    CCU2D add_1054_35 (.A0(d_d_tmp[68]), .B0(n6166), .C0(n6167[32]), .D0(d_tmp[68]), 
          .A1(d_d_tmp[69]), .B1(n6166), .C1(n6167[33]), .D1(d_tmp[69]), 
          .CIN(n11428), .COUT(n11429), .S0(d6_71__N_1458[68]), .S1(d6_71__N_1458[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1054_35.INIT0 = 16'hb874;
    defparam add_1054_35.INIT1 = 16'hb874;
    defparam add_1054_35.INJECT1_0 = "NO";
    defparam add_1054_35.INJECT1_1 = "NO";
    CCU2D add_1054_33 (.A0(d_d_tmp[66]), .B0(n6166), .C0(n6167[30]), .D0(d_tmp[66]), 
          .A1(d_d_tmp[67]), .B1(n6166), .C1(n6167[31]), .D1(d_tmp[67]), 
          .CIN(n11427), .COUT(n11428), .S0(d6_71__N_1458[66]), .S1(d6_71__N_1458[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1054_33.INIT0 = 16'hb874;
    defparam add_1054_33.INIT1 = 16'hb874;
    defparam add_1054_33.INJECT1_0 = "NO";
    defparam add_1054_33.INJECT1_1 = "NO";
    CCU2D add_1054_31 (.A0(d_d_tmp[64]), .B0(n6166), .C0(n6167[28]), .D0(d_tmp[64]), 
          .A1(d_d_tmp[65]), .B1(n6166), .C1(n6167[29]), .D1(d_tmp[65]), 
          .CIN(n11426), .COUT(n11427), .S0(d6_71__N_1458[64]), .S1(d6_71__N_1458[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1054_31.INIT0 = 16'hb874;
    defparam add_1054_31.INIT1 = 16'hb874;
    defparam add_1054_31.INJECT1_0 = "NO";
    defparam add_1054_31.INJECT1_1 = "NO";
    CCU2D add_1054_29 (.A0(d_d_tmp[62]), .B0(n6166), .C0(n6167[26]), .D0(d_tmp[62]), 
          .A1(d_d_tmp[63]), .B1(n6166), .C1(n6167[27]), .D1(d_tmp[63]), 
          .CIN(n11425), .COUT(n11426), .S0(d6_71__N_1458[62]), .S1(d6_71__N_1458[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1054_29.INIT0 = 16'hb874;
    defparam add_1054_29.INIT1 = 16'hb874;
    defparam add_1054_29.INJECT1_0 = "NO";
    defparam add_1054_29.INJECT1_1 = "NO";
    CCU2D add_1054_27 (.A0(d_d_tmp[60]), .B0(n6166), .C0(n6167[24]), .D0(d_tmp[60]), 
          .A1(d_d_tmp[61]), .B1(n6166), .C1(n6167[25]), .D1(d_tmp[61]), 
          .CIN(n11424), .COUT(n11425), .S0(d6_71__N_1458[60]), .S1(d6_71__N_1458[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1054_27.INIT0 = 16'hb874;
    defparam add_1054_27.INIT1 = 16'hb874;
    defparam add_1054_27.INJECT1_0 = "NO";
    defparam add_1054_27.INJECT1_1 = "NO";
    CCU2D add_1054_25 (.A0(d_d_tmp[58]), .B0(n6166), .C0(n6167[22]), .D0(d_tmp[58]), 
          .A1(d_d_tmp[59]), .B1(n6166), .C1(n6167[23]), .D1(d_tmp[59]), 
          .CIN(n11423), .COUT(n11424), .S0(d6_71__N_1458[58]), .S1(d6_71__N_1458[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1054_25.INIT0 = 16'hb874;
    defparam add_1054_25.INIT1 = 16'hb874;
    defparam add_1054_25.INJECT1_0 = "NO";
    defparam add_1054_25.INJECT1_1 = "NO";
    CCU2D add_1054_23 (.A0(d_d_tmp[56]), .B0(n6166), .C0(n6167[20]), .D0(d_tmp[56]), 
          .A1(d_d_tmp[57]), .B1(n6166), .C1(n6167[21]), .D1(d_tmp[57]), 
          .CIN(n11422), .COUT(n11423), .S0(d6_71__N_1458[56]), .S1(d6_71__N_1458[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1054_23.INIT0 = 16'hb874;
    defparam add_1054_23.INIT1 = 16'hb874;
    defparam add_1054_23.INJECT1_0 = "NO";
    defparam add_1054_23.INJECT1_1 = "NO";
    CCU2D add_1054_21 (.A0(d_d_tmp[54]), .B0(n6166), .C0(n6167[18]), .D0(d_tmp[54]), 
          .A1(d_d_tmp[55]), .B1(n6166), .C1(n6167[19]), .D1(d_tmp[55]), 
          .CIN(n11421), .COUT(n11422), .S0(d6_71__N_1458[54]), .S1(d6_71__N_1458[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1054_21.INIT0 = 16'hb874;
    defparam add_1054_21.INIT1 = 16'hb874;
    defparam add_1054_21.INJECT1_0 = "NO";
    defparam add_1054_21.INJECT1_1 = "NO";
    CCU2D add_1054_19 (.A0(d_d_tmp[52]), .B0(n6166), .C0(n6167[16]), .D0(d_tmp[52]), 
          .A1(d_d_tmp[53]), .B1(n6166), .C1(n6167[17]), .D1(d_tmp[53]), 
          .CIN(n11420), .COUT(n11421), .S0(d6_71__N_1458[52]), .S1(d6_71__N_1458[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1054_19.INIT0 = 16'hb874;
    defparam add_1054_19.INIT1 = 16'hb874;
    defparam add_1054_19.INJECT1_0 = "NO";
    defparam add_1054_19.INJECT1_1 = "NO";
    CCU2D add_1054_17 (.A0(d_d_tmp[50]), .B0(n6166), .C0(n6167[14]), .D0(d_tmp[50]), 
          .A1(d_d_tmp[51]), .B1(n6166), .C1(n6167[15]), .D1(d_tmp[51]), 
          .CIN(n11419), .COUT(n11420), .S0(d6_71__N_1458[50]), .S1(d6_71__N_1458[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1054_17.INIT0 = 16'hb874;
    defparam add_1054_17.INIT1 = 16'hb874;
    defparam add_1054_17.INJECT1_0 = "NO";
    defparam add_1054_17.INJECT1_1 = "NO";
    CCU2D add_1028_28 (.A0(d4[62]), .B0(d5[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[63]), .B1(d5[63]), .C1(GND_net), .D1(GND_net), .CIN(n11782), 
          .COUT(n11783), .S0(n5407[26]), .S1(n5407[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1028_28.INIT0 = 16'h5666;
    defparam add_1028_28.INIT1 = 16'h5666;
    defparam add_1028_28.INJECT1_0 = "NO";
    defparam add_1028_28.INJECT1_1 = "NO";
    CCU2D add_1028_26 (.A0(d4[60]), .B0(d5[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[61]), .B1(d5[61]), .C1(GND_net), .D1(GND_net), .CIN(n11781), 
          .COUT(n11782), .S0(n5407[24]), .S1(n5407[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1028_26.INIT0 = 16'h5666;
    defparam add_1028_26.INIT1 = 16'h5666;
    defparam add_1028_26.INJECT1_0 = "NO";
    defparam add_1028_26.INJECT1_1 = "NO";
    CCU2D add_1028_24 (.A0(d4[58]), .B0(d5[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[59]), .B1(d5[59]), .C1(GND_net), .D1(GND_net), .CIN(n11780), 
          .COUT(n11781), .S0(n5407[22]), .S1(n5407[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1028_24.INIT0 = 16'h5666;
    defparam add_1028_24.INIT1 = 16'h5666;
    defparam add_1028_24.INJECT1_0 = "NO";
    defparam add_1028_24.INJECT1_1 = "NO";
    CCU2D add_1028_22 (.A0(d4[56]), .B0(d5[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[57]), .B1(d5[57]), .C1(GND_net), .D1(GND_net), .CIN(n11779), 
          .COUT(n11780), .S0(n5407[20]), .S1(n5407[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1028_22.INIT0 = 16'h5666;
    defparam add_1028_22.INIT1 = 16'h5666;
    defparam add_1028_22.INJECT1_0 = "NO";
    defparam add_1028_22.INJECT1_1 = "NO";
    CCU2D add_1028_20 (.A0(d4[54]), .B0(d5[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[55]), .B1(d5[55]), .C1(GND_net), .D1(GND_net), .CIN(n11778), 
          .COUT(n11779), .S0(n5407[18]), .S1(n5407[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1028_20.INIT0 = 16'h5666;
    defparam add_1028_20.INIT1 = 16'h5666;
    defparam add_1028_20.INJECT1_0 = "NO";
    defparam add_1028_20.INJECT1_1 = "NO";
    CCU2D add_1028_18 (.A0(d4[52]), .B0(d5[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[53]), .B1(d5[53]), .C1(GND_net), .D1(GND_net), .CIN(n11777), 
          .COUT(n11778), .S0(n5407[16]), .S1(n5407[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1028_18.INIT0 = 16'h5666;
    defparam add_1028_18.INIT1 = 16'h5666;
    defparam add_1028_18.INJECT1_0 = "NO";
    defparam add_1028_18.INJECT1_1 = "NO";
    CCU2D add_1028_16 (.A0(d4[50]), .B0(d5[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[51]), .B1(d5[51]), .C1(GND_net), .D1(GND_net), .CIN(n11776), 
          .COUT(n11777), .S0(n5407[14]), .S1(n5407[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1028_16.INIT0 = 16'h5666;
    defparam add_1028_16.INIT1 = 16'h5666;
    defparam add_1028_16.INJECT1_0 = "NO";
    defparam add_1028_16.INJECT1_1 = "NO";
    CCU2D add_1014_5 (.A0(d2[38]), .B0(n4950), .C0(n4951[2]), .D0(d1[38]), 
          .A1(d2[39]), .B1(n4950), .C1(n4951[3]), .D1(d1[39]), .CIN(n11874), 
          .COUT(n11875), .S0(d2_71__N_489[38]), .S1(d2_71__N_489[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1014_5.INIT0 = 16'h74b8;
    defparam add_1014_5.INIT1 = 16'h74b8;
    defparam add_1014_5.INJECT1_0 = "NO";
    defparam add_1014_5.INJECT1_1 = "NO";
    CCU2D add_1014_9 (.A0(d2[42]), .B0(n4950), .C0(n4951[6]), .D0(d1[42]), 
          .A1(d2[43]), .B1(n4950), .C1(n4951[7]), .D1(d1[43]), .CIN(n11876), 
          .COUT(n11877), .S0(d2_71__N_489[42]), .S1(d2_71__N_489[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1014_9.INIT0 = 16'h74b8;
    defparam add_1014_9.INIT1 = 16'h74b8;
    defparam add_1014_9.INJECT1_0 = "NO";
    defparam add_1014_9.INJECT1_1 = "NO";
    LUT4 i4_2_lut (.A(n12867), .B(count[2]), .Z(n16)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i4_2_lut.init = 16'heeee;
    LUT4 i5849_4_lut (.A(n13248), .B(n13), .C(n13250), .D(n13228), .Z(count_15__N_1457)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i5849_4_lut.init = 16'h2000;
    LUT4 i5799_4_lut (.A(count[0]), .B(count[8]), .C(count[1]), .D(count[7]), 
         .Z(n13248)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5799_4_lut.init = 16'h8000;
    LUT4 i5901_2_lut (.A(n31), .B(n14125), .Z(n8412)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam i5901_2_lut.init = 16'hdddd;
    FD1S3IX count__i0 (.D(count_15__N_1441[0]), .CK(osc_clk), .CD(osc_clk_enable_743), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i0.GSR = "ENABLED";
    CCU2D add_1013_24 (.A0(d1[58]), .B0(d2[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[59]), .B1(d2[59]), .C1(GND_net), .D1(GND_net), .CIN(n11903), 
          .COUT(n11904), .S0(n4951[22]), .S1(n4951[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1013_24.INIT0 = 16'h5666;
    defparam add_1013_24.INIT1 = 16'h5666;
    defparam add_1013_24.INJECT1_0 = "NO";
    defparam add_1013_24.INJECT1_1 = "NO";
    CCU2D add_1013_22 (.A0(d1[56]), .B0(d2[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[57]), .B1(d2[57]), .C1(GND_net), .D1(GND_net), .CIN(n11902), 
          .COUT(n11903), .S0(n4951[20]), .S1(n4951[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1013_22.INIT0 = 16'h5666;
    defparam add_1013_22.INIT1 = 16'h5666;
    defparam add_1013_22.INJECT1_0 = "NO";
    defparam add_1013_22.INJECT1_1 = "NO";
    CCU2D add_1013_20 (.A0(d1[54]), .B0(d2[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[55]), .B1(d2[55]), .C1(GND_net), .D1(GND_net), .CIN(n11901), 
          .COUT(n11902), .S0(n4951[18]), .S1(n4951[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1013_20.INIT0 = 16'h5666;
    defparam add_1013_20.INIT1 = 16'h5666;
    defparam add_1013_20.INJECT1_0 = "NO";
    defparam add_1013_20.INJECT1_1 = "NO";
    LUT4 i1_2_lut (.A(n12867), .B(count[3]), .Z(n13)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut.init = 16'hbbbb;
    CCU2D add_1028_14 (.A0(d4[48]), .B0(d5[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[49]), .B1(d5[49]), .C1(GND_net), .D1(GND_net), .CIN(n11775), 
          .COUT(n11776), .S0(n5407[12]), .S1(n5407[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1028_14.INIT0 = 16'h5666;
    defparam add_1028_14.INIT1 = 16'h5666;
    defparam add_1028_14.INJECT1_0 = "NO";
    defparam add_1028_14.INJECT1_1 = "NO";
    CCU2D add_1028_12 (.A0(d4[46]), .B0(d5[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[47]), .B1(d5[47]), .C1(GND_net), .D1(GND_net), .CIN(n11774), 
          .COUT(n11775), .S0(n5407[10]), .S1(n5407[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1028_12.INIT0 = 16'h5666;
    defparam add_1028_12.INIT1 = 16'h5666;
    defparam add_1028_12.INJECT1_0 = "NO";
    defparam add_1028_12.INJECT1_1 = "NO";
    FD1S3IX count__i1 (.D(n375[1]), .CK(osc_clk), .CD(n8412), .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i1.GSR = "ENABLED";
    CCU2D add_1028_10 (.A0(d4[44]), .B0(d5[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[45]), .B1(d5[45]), .C1(GND_net), .D1(GND_net), .CIN(n11773), 
          .COUT(n11774), .S0(n5407[8]), .S1(n5407[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1028_10.INIT0 = 16'h5666;
    defparam add_1028_10.INIT1 = 16'h5666;
    defparam add_1028_10.INJECT1_0 = "NO";
    defparam add_1028_10.INJECT1_1 = "NO";
    CCU2D add_1028_8 (.A0(d4[42]), .B0(d5[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[43]), .B1(d5[43]), .C1(GND_net), .D1(GND_net), .CIN(n11772), 
          .COUT(n11773), .S0(n5407[6]), .S1(n5407[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1028_8.INIT0 = 16'h5666;
    defparam add_1028_8.INIT1 = 16'h5666;
    defparam add_1028_8.INJECT1_0 = "NO";
    defparam add_1028_8.INJECT1_1 = "NO";
    CCU2D add_1028_6 (.A0(d4[40]), .B0(d5[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[41]), .B1(d5[41]), .C1(GND_net), .D1(GND_net), .CIN(n11771), 
          .COUT(n11772), .S0(n5407[4]), .S1(n5407[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1028_6.INIT0 = 16'h5666;
    defparam add_1028_6.INIT1 = 16'h5666;
    defparam add_1028_6.INJECT1_0 = "NO";
    defparam add_1028_6.INJECT1_1 = "NO";
    CCU2D add_1028_4 (.A0(d4[38]), .B0(d5[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[39]), .B1(d5[39]), .C1(GND_net), .D1(GND_net), .CIN(n11770), 
          .COUT(n11771), .S0(n5407[2]), .S1(n5407[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1028_4.INIT0 = 16'h5666;
    defparam add_1028_4.INIT1 = 16'h5666;
    defparam add_1028_4.INJECT1_0 = "NO";
    defparam add_1028_4.INJECT1_1 = "NO";
    CCU2D add_1028_2 (.A0(d4[36]), .B0(d5[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[37]), .B1(d5[37]), .C1(GND_net), .D1(GND_net), .COUT(n11770), 
          .S1(n5407[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1028_2.INIT0 = 16'h7000;
    defparam add_1028_2.INIT1 = 16'h5666;
    defparam add_1028_2.INJECT1_0 = "NO";
    defparam add_1028_2.INJECT1_1 = "NO";
    CCU2D add_1029_37 (.A0(d5[70]), .B0(n5406), .C0(n5407[34]), .D0(d4[70]), 
          .A1(d5[71]), .B1(n5406), .C1(n5407[35]), .D1(d4[71]), .CIN(n11767), 
          .S0(d5_71__N_705[70]), .S1(d5_71__N_705[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1029_37.INIT0 = 16'h74b8;
    defparam add_1029_37.INIT1 = 16'h74b8;
    defparam add_1029_37.INJECT1_0 = "NO";
    defparam add_1029_37.INJECT1_1 = "NO";
    CCU2D add_1029_35 (.A0(d5[68]), .B0(n5406), .C0(n5407[32]), .D0(d4[68]), 
          .A1(d5[69]), .B1(n5406), .C1(n5407[33]), .D1(d4[69]), .CIN(n11766), 
          .COUT(n11767), .S0(d5_71__N_705[68]), .S1(d5_71__N_705[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1029_35.INIT0 = 16'h74b8;
    defparam add_1029_35.INIT1 = 16'h74b8;
    defparam add_1029_35.INJECT1_0 = "NO";
    defparam add_1029_35.INJECT1_1 = "NO";
    CCU2D add_1029_33 (.A0(d5[66]), .B0(n5406), .C0(n5407[30]), .D0(d4[66]), 
          .A1(d5[67]), .B1(n5406), .C1(n5407[31]), .D1(d4[67]), .CIN(n11765), 
          .COUT(n11766), .S0(d5_71__N_705[66]), .S1(d5_71__N_705[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1029_33.INIT0 = 16'h74b8;
    defparam add_1029_33.INIT1 = 16'h74b8;
    defparam add_1029_33.INJECT1_0 = "NO";
    defparam add_1029_33.INJECT1_1 = "NO";
    CCU2D add_1029_31 (.A0(d5[64]), .B0(n5406), .C0(n5407[28]), .D0(d4[64]), 
          .A1(d5[65]), .B1(n5406), .C1(n5407[29]), .D1(d4[65]), .CIN(n11764), 
          .COUT(n11765), .S0(d5_71__N_705[64]), .S1(d5_71__N_705[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1029_31.INIT0 = 16'h74b8;
    defparam add_1029_31.INIT1 = 16'h74b8;
    defparam add_1029_31.INJECT1_0 = "NO";
    defparam add_1029_31.INJECT1_1 = "NO";
    CCU2D add_1029_29 (.A0(d5[62]), .B0(n5406), .C0(n5407[26]), .D0(d4[62]), 
          .A1(d5[63]), .B1(n5406), .C1(n5407[27]), .D1(d4[63]), .CIN(n11763), 
          .COUT(n11764), .S0(d5_71__N_705[62]), .S1(d5_71__N_705[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1029_29.INIT0 = 16'h74b8;
    defparam add_1029_29.INIT1 = 16'h74b8;
    defparam add_1029_29.INJECT1_0 = "NO";
    defparam add_1029_29.INJECT1_1 = "NO";
    CCU2D add_1029_27 (.A0(d5[60]), .B0(n5406), .C0(n5407[24]), .D0(d4[60]), 
          .A1(d5[61]), .B1(n5406), .C1(n5407[25]), .D1(d4[61]), .CIN(n11762), 
          .COUT(n11763), .S0(d5_71__N_705[60]), .S1(d5_71__N_705[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1029_27.INIT0 = 16'h74b8;
    defparam add_1029_27.INIT1 = 16'h74b8;
    defparam add_1029_27.INJECT1_0 = "NO";
    defparam add_1029_27.INJECT1_1 = "NO";
    CCU2D add_1029_25 (.A0(d5[58]), .B0(n5406), .C0(n5407[22]), .D0(d4[58]), 
          .A1(d5[59]), .B1(n5406), .C1(n5407[23]), .D1(d4[59]), .CIN(n11761), 
          .COUT(n11762), .S0(d5_71__N_705[58]), .S1(d5_71__N_705[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1029_25.INIT0 = 16'h74b8;
    defparam add_1029_25.INIT1 = 16'h74b8;
    defparam add_1029_25.INJECT1_0 = "NO";
    defparam add_1029_25.INJECT1_1 = "NO";
    CCU2D add_1029_23 (.A0(d5[56]), .B0(n5406), .C0(n5407[20]), .D0(d4[56]), 
          .A1(d5[57]), .B1(n5406), .C1(n5407[21]), .D1(d4[57]), .CIN(n11760), 
          .COUT(n11761), .S0(d5_71__N_705[56]), .S1(d5_71__N_705[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1029_23.INIT0 = 16'h74b8;
    defparam add_1029_23.INIT1 = 16'h74b8;
    defparam add_1029_23.INJECT1_0 = "NO";
    defparam add_1029_23.INJECT1_1 = "NO";
    LUT4 i4791_2_lut (.A(d4[36]), .B(d5[36]), .Z(n5407[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4791_2_lut.init = 16'h6666;
    CCU2D add_1029_21 (.A0(d5[54]), .B0(n5406), .C0(n5407[18]), .D0(d4[54]), 
          .A1(d5[55]), .B1(n5406), .C1(n5407[19]), .D1(d4[55]), .CIN(n11759), 
          .COUT(n11760), .S0(d5_71__N_705[54]), .S1(d5_71__N_705[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1029_21.INIT0 = 16'h74b8;
    defparam add_1029_21.INIT1 = 16'h74b8;
    defparam add_1029_21.INJECT1_0 = "NO";
    defparam add_1029_21.INJECT1_1 = "NO";
    CCU2D add_1029_19 (.A0(d5[52]), .B0(n5406), .C0(n5407[16]), .D0(d4[52]), 
          .A1(d5[53]), .B1(n5406), .C1(n5407[17]), .D1(d4[53]), .CIN(n11758), 
          .COUT(n11759), .S0(d5_71__N_705[52]), .S1(d5_71__N_705[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1029_19.INIT0 = 16'h74b8;
    defparam add_1029_19.INIT1 = 16'h74b8;
    defparam add_1029_19.INJECT1_0 = "NO";
    defparam add_1029_19.INJECT1_1 = "NO";
    CCU2D add_1029_17 (.A0(d5[50]), .B0(n5406), .C0(n5407[14]), .D0(d4[50]), 
          .A1(d5[51]), .B1(n5406), .C1(n5407[15]), .D1(d4[51]), .CIN(n11757), 
          .COUT(n11758), .S0(d5_71__N_705[50]), .S1(d5_71__N_705[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1029_17.INIT0 = 16'h74b8;
    defparam add_1029_17.INIT1 = 16'h74b8;
    defparam add_1029_17.INJECT1_0 = "NO";
    defparam add_1029_17.INJECT1_1 = "NO";
    LUT4 i2723_2_lut (.A(n375[11]), .B(n31), .Z(count_15__N_1441[11])) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(86[13] 89[16])
    defparam i2723_2_lut.init = 16'hbbbb;
    CCU2D add_1029_15 (.A0(d5[48]), .B0(n5406), .C0(n5407[12]), .D0(d4[48]), 
          .A1(d5[49]), .B1(n5406), .C1(n5407[13]), .D1(d4[49]), .CIN(n11756), 
          .COUT(n11757), .S0(d5_71__N_705[48]), .S1(d5_71__N_705[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1029_15.INIT0 = 16'h74b8;
    defparam add_1029_15.INIT1 = 16'h74b8;
    defparam add_1029_15.INJECT1_0 = "NO";
    defparam add_1029_15.INJECT1_1 = "NO";
    CCU2D add_1029_13 (.A0(d5[46]), .B0(n5406), .C0(n5407[10]), .D0(d4[46]), 
          .A1(d5[47]), .B1(n5406), .C1(n5407[11]), .D1(d4[47]), .CIN(n11755), 
          .COUT(n11756), .S0(d5_71__N_705[46]), .S1(d5_71__N_705[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1029_13.INIT0 = 16'h74b8;
    defparam add_1029_13.INIT1 = 16'h74b8;
    defparam add_1029_13.INJECT1_0 = "NO";
    defparam add_1029_13.INJECT1_1 = "NO";
    CCU2D add_1029_11 (.A0(d5[44]), .B0(n5406), .C0(n5407[8]), .D0(d4[44]), 
          .A1(d5[45]), .B1(n5406), .C1(n5407[9]), .D1(d4[45]), .CIN(n11754), 
          .COUT(n11755), .S0(d5_71__N_705[44]), .S1(d5_71__N_705[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1029_11.INIT0 = 16'h74b8;
    defparam add_1029_11.INIT1 = 16'h74b8;
    defparam add_1029_11.INJECT1_0 = "NO";
    defparam add_1029_11.INJECT1_1 = "NO";
    CCU2D add_1029_9 (.A0(d5[42]), .B0(n5406), .C0(n5407[6]), .D0(d4[42]), 
          .A1(d5[43]), .B1(n5406), .C1(n5407[7]), .D1(d4[43]), .CIN(n11753), 
          .COUT(n11754), .S0(d5_71__N_705[42]), .S1(d5_71__N_705[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1029_9.INIT0 = 16'h74b8;
    defparam add_1029_9.INIT1 = 16'h74b8;
    defparam add_1029_9.INJECT1_0 = "NO";
    defparam add_1029_9.INJECT1_1 = "NO";
    CCU2D add_1029_7 (.A0(d5[40]), .B0(n5406), .C0(n5407[4]), .D0(d4[40]), 
          .A1(d5[41]), .B1(n5406), .C1(n5407[5]), .D1(d4[41]), .CIN(n11752), 
          .COUT(n11753), .S0(d5_71__N_705[40]), .S1(d5_71__N_705[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1029_7.INIT0 = 16'h74b8;
    defparam add_1029_7.INIT1 = 16'h74b8;
    defparam add_1029_7.INJECT1_0 = "NO";
    defparam add_1029_7.INJECT1_1 = "NO";
    CCU2D add_1029_5 (.A0(d5[38]), .B0(n5406), .C0(n5407[2]), .D0(d4[38]), 
          .A1(d5[39]), .B1(n5406), .C1(n5407[3]), .D1(d4[39]), .CIN(n11751), 
          .COUT(n11752), .S0(d5_71__N_705[38]), .S1(d5_71__N_705[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1029_5.INIT0 = 16'h74b8;
    defparam add_1029_5.INIT1 = 16'h74b8;
    defparam add_1029_5.INJECT1_0 = "NO";
    defparam add_1029_5.INJECT1_1 = "NO";
    CCU2D add_1029_3 (.A0(d5[36]), .B0(n5406), .C0(n5407[0]), .D0(d4[36]), 
          .A1(d5[37]), .B1(n5406), .C1(n5407[1]), .D1(d4[37]), .CIN(n11750), 
          .COUT(n11751), .S0(d5_71__N_705[36]), .S1(d5_71__N_705[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1029_3.INIT0 = 16'h74b8;
    defparam add_1029_3.INIT1 = 16'h74b8;
    defparam add_1029_3.INJECT1_0 = "NO";
    defparam add_1029_3.INJECT1_1 = "NO";
    CCU2D add_1029_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5406), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11750));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1029_1.INIT0 = 16'hF000;
    defparam add_1029_1.INIT1 = 16'h0555;
    defparam add_1029_1.INJECT1_0 = "NO";
    defparam add_1029_1.INJECT1_1 = "NO";
    LUT4 i5801_4_lut (.A(count[9]), .B(count[2]), .C(count[4]), .D(count[6]), 
         .Z(n13250)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5801_4_lut.init = 16'h8000;
    CCU2D add_1054_15 (.A0(d_d_tmp[48]), .B0(n6166), .C0(n6167[12]), .D0(d_tmp[48]), 
          .A1(d_d_tmp[49]), .B1(n6166), .C1(n6167[13]), .D1(d_tmp[49]), 
          .CIN(n11418), .COUT(n11419), .S0(d6_71__N_1458[48]), .S1(d6_71__N_1458[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1054_15.INIT0 = 16'hb874;
    defparam add_1054_15.INIT1 = 16'hb874;
    defparam add_1054_15.INJECT1_0 = "NO";
    defparam add_1054_15.INJECT1_1 = "NO";
    FD1P3AX d_tmp_i0_i1 (.D(d5[1]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i2 (.D(d5[2]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i3 (.D(d5[3]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i4 (.D(d5[4]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i5 (.D(d5[5]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i6 (.D(d5[6]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i7 (.D(d5[7]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i8 (.D(d5[8]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i9 (.D(d5[9]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i10 (.D(d5[10]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i11 (.D(d5[11]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i12 (.D(d5[12]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i13 (.D(d5[13]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i14 (.D(d5[14]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i15 (.D(d5[15]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i16 (.D(d5[16]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i17 (.D(d5[17]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i18 (.D(d5[18]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i19 (.D(d5[19]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i20 (.D(d5[20]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i21 (.D(d5[21]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i22 (.D(d5[22]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i23 (.D(d5[23]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i24 (.D(d5[24]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i25 (.D(d5[25]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i26 (.D(d5[26]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i27 (.D(d5[27]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i28 (.D(d5[28]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i29 (.D(d5[29]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i30 (.D(d5[30]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i31 (.D(d5[31]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i32 (.D(d5[32]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i33 (.D(d5[33]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i34 (.D(d5[34]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i35 (.D(d5[35]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i36 (.D(d5[36]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i37 (.D(d5[37]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i38 (.D(d5[38]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i39 (.D(d5[39]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i40 (.D(d5[40]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i41 (.D(d5[41]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i42 (.D(d5[42]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i43 (.D(d5[43]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i44 (.D(d5[44]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i45 (.D(d5[45]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i46 (.D(d5[46]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i47 (.D(d5[47]), .SP(osc_clk_enable_743), .CK(osc_clk), 
            .Q(d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i48 (.D(d5[48]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i49 (.D(d5[49]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i50 (.D(d5[50]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i51 (.D(d5[51]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i52 (.D(d5[52]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i53 (.D(d5[53]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i54 (.D(d5[54]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i55 (.D(d5[55]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i56 (.D(d5[56]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i57 (.D(d5[57]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i58 (.D(d5[58]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i59 (.D(d5[59]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i60 (.D(d5[60]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i61 (.D(d5[61]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i62 (.D(d5[62]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i63 (.D(d5[63]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i64 (.D(d5[64]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i65 (.D(d5[65]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i66 (.D(d5[66]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i67 (.D(d5[67]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i68 (.D(d5[68]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i69 (.D(d5[69]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i70 (.D(d5[70]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i71 (.D(d5[71]), .SP(count_15__N_1457), .CK(osc_clk), 
            .Q(d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i1 (.D(d_tmp[1]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i2 (.D(d_tmp[2]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i3 (.D(d_tmp[3]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i4 (.D(d_tmp[4]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i5 (.D(d_tmp[5]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i6 (.D(d_tmp[6]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i7 (.D(d_tmp[7]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i8 (.D(d_tmp[8]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i9 (.D(d_tmp[9]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i10 (.D(d_tmp[10]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i11 (.D(d_tmp[11]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i12 (.D(d_tmp[12]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i13 (.D(d_tmp[13]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i14 (.D(d_tmp[14]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i15 (.D(d_tmp[15]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i16 (.D(d_tmp[16]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i17 (.D(d_tmp[17]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i18 (.D(d_tmp[18]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i19 (.D(d_tmp[19]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i20 (.D(d_tmp[20]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i21 (.D(d_tmp[21]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i22 (.D(d_tmp[22]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i23 (.D(d_tmp[23]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i24 (.D(d_tmp[24]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i25 (.D(d_tmp[25]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i26 (.D(d_tmp[26]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i27 (.D(d_tmp[27]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i28 (.D(d_tmp[28]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i29 (.D(d_tmp[29]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i30 (.D(d_tmp[30]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i31 (.D(d_tmp[31]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i32 (.D(d_tmp[32]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i33 (.D(d_tmp[33]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i34 (.D(d_tmp[34]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i35 (.D(d_tmp[35]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i36 (.D(d_tmp[36]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i37 (.D(d_tmp[37]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i38 (.D(d_tmp[38]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i39 (.D(d_tmp[39]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i40 (.D(d_tmp[40]), .SP(osc_clk_enable_783), .CK(osc_clk), 
            .Q(d_d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i41 (.D(d_tmp[41]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i42 (.D(d_tmp[42]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i43 (.D(d_tmp[43]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i44 (.D(d_tmp[44]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i45 (.D(d_tmp[45]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i46 (.D(d_tmp[46]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i47 (.D(d_tmp[47]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i48 (.D(d_tmp[48]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i49 (.D(d_tmp[49]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i50 (.D(d_tmp[50]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i51 (.D(d_tmp[51]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i52 (.D(d_tmp[52]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i53 (.D(d_tmp[53]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i54 (.D(d_tmp[54]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i55 (.D(d_tmp[55]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i56 (.D(d_tmp[56]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i57 (.D(d_tmp[57]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i58 (.D(d_tmp[58]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i59 (.D(d_tmp[59]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i60 (.D(d_tmp[60]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i61 (.D(d_tmp[61]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i62 (.D(d_tmp[62]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i63 (.D(d_tmp[63]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i64 (.D(d_tmp[64]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i65 (.D(d_tmp[65]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i66 (.D(d_tmp[66]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i67 (.D(d_tmp[67]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i68 (.D(d_tmp[68]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i69 (.D(d_tmp[69]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i70 (.D(d_tmp[70]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i71 (.D(d_tmp[71]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d_d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d_tmp_i0_i71.GSR = "ENABLED";
    FD1S3AX d2_i1 (.D(d2_71__N_489[1]), .CK(osc_clk), .Q(d2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i1.GSR = "ENABLED";
    FD1S3AX d2_i2 (.D(d2_71__N_489[2]), .CK(osc_clk), .Q(d2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i2.GSR = "ENABLED";
    FD1S3AX d2_i3 (.D(d2_71__N_489[3]), .CK(osc_clk), .Q(d2[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i3.GSR = "ENABLED";
    FD1S3AX d2_i4 (.D(d2_71__N_489[4]), .CK(osc_clk), .Q(d2[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i4.GSR = "ENABLED";
    FD1S3AX d2_i5 (.D(d2_71__N_489[5]), .CK(osc_clk), .Q(d2[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i5.GSR = "ENABLED";
    FD1S3AX d2_i6 (.D(d2_71__N_489[6]), .CK(osc_clk), .Q(d2[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i6.GSR = "ENABLED";
    FD1S3AX d2_i7 (.D(d2_71__N_489[7]), .CK(osc_clk), .Q(d2[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i7.GSR = "ENABLED";
    FD1S3AX d2_i8 (.D(d2_71__N_489[8]), .CK(osc_clk), .Q(d2[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i8.GSR = "ENABLED";
    FD1S3AX d2_i9 (.D(d2_71__N_489[9]), .CK(osc_clk), .Q(d2[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i9.GSR = "ENABLED";
    FD1S3AX d2_i10 (.D(d2_71__N_489[10]), .CK(osc_clk), .Q(d2[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i10.GSR = "ENABLED";
    FD1S3AX d2_i11 (.D(d2_71__N_489[11]), .CK(osc_clk), .Q(d2[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i11.GSR = "ENABLED";
    FD1S3AX d2_i12 (.D(d2_71__N_489[12]), .CK(osc_clk), .Q(d2[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i12.GSR = "ENABLED";
    FD1S3AX d2_i13 (.D(d2_71__N_489[13]), .CK(osc_clk), .Q(d2[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i13.GSR = "ENABLED";
    FD1S3AX d2_i14 (.D(d2_71__N_489[14]), .CK(osc_clk), .Q(d2[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i14.GSR = "ENABLED";
    FD1S3AX d2_i15 (.D(d2_71__N_489[15]), .CK(osc_clk), .Q(d2[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i15.GSR = "ENABLED";
    FD1S3AX d2_i16 (.D(d2_71__N_489[16]), .CK(osc_clk), .Q(d2[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i16.GSR = "ENABLED";
    FD1S3AX d2_i17 (.D(d2_71__N_489[17]), .CK(osc_clk), .Q(d2[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i17.GSR = "ENABLED";
    FD1S3AX d2_i18 (.D(d2_71__N_489[18]), .CK(osc_clk), .Q(d2[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i18.GSR = "ENABLED";
    FD1S3AX d2_i19 (.D(d2_71__N_489[19]), .CK(osc_clk), .Q(d2[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i19.GSR = "ENABLED";
    FD1S3AX d2_i20 (.D(d2_71__N_489[20]), .CK(osc_clk), .Q(d2[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i20.GSR = "ENABLED";
    FD1S3AX d2_i21 (.D(d2_71__N_489[21]), .CK(osc_clk), .Q(d2[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i21.GSR = "ENABLED";
    FD1S3AX d2_i22 (.D(d2_71__N_489[22]), .CK(osc_clk), .Q(d2[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i22.GSR = "ENABLED";
    FD1S3AX d2_i23 (.D(d2_71__N_489[23]), .CK(osc_clk), .Q(d2[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i23.GSR = "ENABLED";
    FD1S3AX d2_i24 (.D(d2_71__N_489[24]), .CK(osc_clk), .Q(d2[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i24.GSR = "ENABLED";
    FD1S3AX d2_i25 (.D(d2_71__N_489[25]), .CK(osc_clk), .Q(d2[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i25.GSR = "ENABLED";
    FD1S3AX d2_i26 (.D(d2_71__N_489[26]), .CK(osc_clk), .Q(d2[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i26.GSR = "ENABLED";
    FD1S3AX d2_i27 (.D(d2_71__N_489[27]), .CK(osc_clk), .Q(d2[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i27.GSR = "ENABLED";
    FD1S3AX d2_i28 (.D(d2_71__N_489[28]), .CK(osc_clk), .Q(d2[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i28.GSR = "ENABLED";
    FD1S3AX d2_i29 (.D(d2_71__N_489[29]), .CK(osc_clk), .Q(d2[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i29.GSR = "ENABLED";
    FD1S3AX d2_i30 (.D(d2_71__N_489[30]), .CK(osc_clk), .Q(d2[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i30.GSR = "ENABLED";
    FD1S3AX d2_i31 (.D(d2_71__N_489[31]), .CK(osc_clk), .Q(d2[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i31.GSR = "ENABLED";
    FD1S3AX d2_i32 (.D(d2_71__N_489[32]), .CK(osc_clk), .Q(d2[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i32.GSR = "ENABLED";
    FD1S3AX d2_i33 (.D(d2_71__N_489[33]), .CK(osc_clk), .Q(d2[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i33.GSR = "ENABLED";
    FD1S3AX d2_i34 (.D(d2_71__N_489[34]), .CK(osc_clk), .Q(d2[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i34.GSR = "ENABLED";
    FD1S3AX d2_i35 (.D(d2_71__N_489[35]), .CK(osc_clk), .Q(d2[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i35.GSR = "ENABLED";
    FD1S3AX d2_i36 (.D(d2_71__N_489[36]), .CK(osc_clk), .Q(d2[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i36.GSR = "ENABLED";
    FD1S3AX d2_i37 (.D(d2_71__N_489[37]), .CK(osc_clk), .Q(d2[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i37.GSR = "ENABLED";
    FD1S3AX d2_i38 (.D(d2_71__N_489[38]), .CK(osc_clk), .Q(d2[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i38.GSR = "ENABLED";
    FD1S3AX d2_i39 (.D(d2_71__N_489[39]), .CK(osc_clk), .Q(d2[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i39.GSR = "ENABLED";
    FD1S3AX d2_i40 (.D(d2_71__N_489[40]), .CK(osc_clk), .Q(d2[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i40.GSR = "ENABLED";
    FD1S3AX d2_i41 (.D(d2_71__N_489[41]), .CK(osc_clk), .Q(d2[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i41.GSR = "ENABLED";
    FD1S3AX d2_i42 (.D(d2_71__N_489[42]), .CK(osc_clk), .Q(d2[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i42.GSR = "ENABLED";
    FD1S3AX d2_i43 (.D(d2_71__N_489[43]), .CK(osc_clk), .Q(d2[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i43.GSR = "ENABLED";
    FD1S3AX d2_i44 (.D(d2_71__N_489[44]), .CK(osc_clk), .Q(d2[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i44.GSR = "ENABLED";
    FD1S3AX d2_i45 (.D(d2_71__N_489[45]), .CK(osc_clk), .Q(d2[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i45.GSR = "ENABLED";
    FD1S3AX d2_i46 (.D(d2_71__N_489[46]), .CK(osc_clk), .Q(d2[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i46.GSR = "ENABLED";
    FD1S3AX d2_i47 (.D(d2_71__N_489[47]), .CK(osc_clk), .Q(d2[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i47.GSR = "ENABLED";
    FD1S3AX d2_i48 (.D(d2_71__N_489[48]), .CK(osc_clk), .Q(d2[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i48.GSR = "ENABLED";
    FD1S3AX d2_i49 (.D(d2_71__N_489[49]), .CK(osc_clk), .Q(d2[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i49.GSR = "ENABLED";
    FD1S3AX d2_i50 (.D(d2_71__N_489[50]), .CK(osc_clk), .Q(d2[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i50.GSR = "ENABLED";
    FD1S3AX d2_i51 (.D(d2_71__N_489[51]), .CK(osc_clk), .Q(d2[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i51.GSR = "ENABLED";
    FD1S3AX d2_i52 (.D(d2_71__N_489[52]), .CK(osc_clk), .Q(d2[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i52.GSR = "ENABLED";
    FD1S3AX d2_i53 (.D(d2_71__N_489[53]), .CK(osc_clk), .Q(d2[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i53.GSR = "ENABLED";
    FD1S3AX d2_i54 (.D(d2_71__N_489[54]), .CK(osc_clk), .Q(d2[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i54.GSR = "ENABLED";
    FD1S3AX d2_i55 (.D(d2_71__N_489[55]), .CK(osc_clk), .Q(d2[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i55.GSR = "ENABLED";
    FD1S3AX d2_i56 (.D(d2_71__N_489[56]), .CK(osc_clk), .Q(d2[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i56.GSR = "ENABLED";
    FD1S3AX d2_i57 (.D(d2_71__N_489[57]), .CK(osc_clk), .Q(d2[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i57.GSR = "ENABLED";
    FD1S3AX d2_i58 (.D(d2_71__N_489[58]), .CK(osc_clk), .Q(d2[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i58.GSR = "ENABLED";
    FD1S3AX d2_i59 (.D(d2_71__N_489[59]), .CK(osc_clk), .Q(d2[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i59.GSR = "ENABLED";
    FD1S3AX d2_i60 (.D(d2_71__N_489[60]), .CK(osc_clk), .Q(d2[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i60.GSR = "ENABLED";
    FD1S3AX d2_i61 (.D(d2_71__N_489[61]), .CK(osc_clk), .Q(d2[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i61.GSR = "ENABLED";
    FD1S3AX d2_i62 (.D(d2_71__N_489[62]), .CK(osc_clk), .Q(d2[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i62.GSR = "ENABLED";
    FD1S3AX d2_i63 (.D(d2_71__N_489[63]), .CK(osc_clk), .Q(d2[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i63.GSR = "ENABLED";
    FD1S3AX d2_i64 (.D(d2_71__N_489[64]), .CK(osc_clk), .Q(d2[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i64.GSR = "ENABLED";
    FD1S3AX d2_i65 (.D(d2_71__N_489[65]), .CK(osc_clk), .Q(d2[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i65.GSR = "ENABLED";
    FD1S3AX d2_i66 (.D(d2_71__N_489[66]), .CK(osc_clk), .Q(d2[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i66.GSR = "ENABLED";
    FD1S3AX d2_i67 (.D(d2_71__N_489[67]), .CK(osc_clk), .Q(d2[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i67.GSR = "ENABLED";
    FD1S3AX d2_i68 (.D(d2_71__N_489[68]), .CK(osc_clk), .Q(d2[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i68.GSR = "ENABLED";
    FD1S3AX d2_i69 (.D(d2_71__N_489[69]), .CK(osc_clk), .Q(d2[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i69.GSR = "ENABLED";
    FD1S3AX d2_i70 (.D(d2_71__N_489[70]), .CK(osc_clk), .Q(d2[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i70.GSR = "ENABLED";
    FD1S3AX d2_i71 (.D(d2_71__N_489[71]), .CK(osc_clk), .Q(d2[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d2_i71.GSR = "ENABLED";
    FD1S3AX d3_i1 (.D(d3_71__N_561[1]), .CK(osc_clk), .Q(d3[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i1.GSR = "ENABLED";
    FD1S3AX d3_i2 (.D(d3_71__N_561[2]), .CK(osc_clk), .Q(d3[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i2.GSR = "ENABLED";
    FD1S3AX d3_i3 (.D(d3_71__N_561[3]), .CK(osc_clk), .Q(d3[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i3.GSR = "ENABLED";
    FD1S3AX d3_i4 (.D(d3_71__N_561[4]), .CK(osc_clk), .Q(d3[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i4.GSR = "ENABLED";
    FD1S3AX d3_i5 (.D(d3_71__N_561[5]), .CK(osc_clk), .Q(d3[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i5.GSR = "ENABLED";
    FD1S3AX d3_i6 (.D(d3_71__N_561[6]), .CK(osc_clk), .Q(d3[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i6.GSR = "ENABLED";
    FD1S3AX d3_i7 (.D(d3_71__N_561[7]), .CK(osc_clk), .Q(d3[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i7.GSR = "ENABLED";
    FD1S3AX d3_i8 (.D(d3_71__N_561[8]), .CK(osc_clk), .Q(d3[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i8.GSR = "ENABLED";
    FD1S3AX d3_i9 (.D(d3_71__N_561[9]), .CK(osc_clk), .Q(d3[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i9.GSR = "ENABLED";
    FD1S3AX d3_i10 (.D(d3_71__N_561[10]), .CK(osc_clk), .Q(d3[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i10.GSR = "ENABLED";
    FD1S3AX d3_i11 (.D(d3_71__N_561[11]), .CK(osc_clk), .Q(d3[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i11.GSR = "ENABLED";
    FD1S3AX d3_i12 (.D(d3_71__N_561[12]), .CK(osc_clk), .Q(d3[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i12.GSR = "ENABLED";
    FD1S3AX d3_i13 (.D(d3_71__N_561[13]), .CK(osc_clk), .Q(d3[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i13.GSR = "ENABLED";
    FD1S3AX d3_i14 (.D(d3_71__N_561[14]), .CK(osc_clk), .Q(d3[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i14.GSR = "ENABLED";
    FD1S3AX d3_i15 (.D(d3_71__N_561[15]), .CK(osc_clk), .Q(d3[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i15.GSR = "ENABLED";
    FD1S3AX d3_i16 (.D(d3_71__N_561[16]), .CK(osc_clk), .Q(d3[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i16.GSR = "ENABLED";
    FD1S3AX d3_i17 (.D(d3_71__N_561[17]), .CK(osc_clk), .Q(d3[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i17.GSR = "ENABLED";
    FD1S3AX d3_i18 (.D(d3_71__N_561[18]), .CK(osc_clk), .Q(d3[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i18.GSR = "ENABLED";
    FD1S3AX d3_i19 (.D(d3_71__N_561[19]), .CK(osc_clk), .Q(d3[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i19.GSR = "ENABLED";
    FD1S3AX d3_i20 (.D(d3_71__N_561[20]), .CK(osc_clk), .Q(d3[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i20.GSR = "ENABLED";
    FD1S3AX d3_i21 (.D(d3_71__N_561[21]), .CK(osc_clk), .Q(d3[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i21.GSR = "ENABLED";
    FD1S3AX d3_i22 (.D(d3_71__N_561[22]), .CK(osc_clk), .Q(d3[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i22.GSR = "ENABLED";
    FD1S3AX d3_i23 (.D(d3_71__N_561[23]), .CK(osc_clk), .Q(d3[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i23.GSR = "ENABLED";
    FD1S3AX d3_i24 (.D(d3_71__N_561[24]), .CK(osc_clk), .Q(d3[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i24.GSR = "ENABLED";
    FD1S3AX d3_i25 (.D(d3_71__N_561[25]), .CK(osc_clk), .Q(d3[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i25.GSR = "ENABLED";
    FD1S3AX d3_i26 (.D(d3_71__N_561[26]), .CK(osc_clk), .Q(d3[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i26.GSR = "ENABLED";
    FD1S3AX d3_i27 (.D(d3_71__N_561[27]), .CK(osc_clk), .Q(d3[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i27.GSR = "ENABLED";
    FD1S3AX d3_i28 (.D(d3_71__N_561[28]), .CK(osc_clk), .Q(d3[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i28.GSR = "ENABLED";
    FD1S3AX d3_i29 (.D(d3_71__N_561[29]), .CK(osc_clk), .Q(d3[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i29.GSR = "ENABLED";
    FD1S3AX d3_i30 (.D(d3_71__N_561[30]), .CK(osc_clk), .Q(d3[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i30.GSR = "ENABLED";
    FD1S3AX d3_i31 (.D(d3_71__N_561[31]), .CK(osc_clk), .Q(d3[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i31.GSR = "ENABLED";
    FD1S3AX d3_i32 (.D(d3_71__N_561[32]), .CK(osc_clk), .Q(d3[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i32.GSR = "ENABLED";
    FD1S3AX d3_i33 (.D(d3_71__N_561[33]), .CK(osc_clk), .Q(d3[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i33.GSR = "ENABLED";
    FD1S3AX d3_i34 (.D(d3_71__N_561[34]), .CK(osc_clk), .Q(d3[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i34.GSR = "ENABLED";
    FD1S3AX d3_i35 (.D(d3_71__N_561[35]), .CK(osc_clk), .Q(d3[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i35.GSR = "ENABLED";
    FD1S3AX d3_i36 (.D(d3_71__N_561[36]), .CK(osc_clk), .Q(d3[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i36.GSR = "ENABLED";
    FD1S3AX d3_i37 (.D(d3_71__N_561[37]), .CK(osc_clk), .Q(d3[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i37.GSR = "ENABLED";
    FD1S3AX d3_i38 (.D(d3_71__N_561[38]), .CK(osc_clk), .Q(d3[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i38.GSR = "ENABLED";
    FD1S3AX d3_i39 (.D(d3_71__N_561[39]), .CK(osc_clk), .Q(d3[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i39.GSR = "ENABLED";
    FD1S3AX d3_i40 (.D(d3_71__N_561[40]), .CK(osc_clk), .Q(d3[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i40.GSR = "ENABLED";
    FD1S3AX d3_i41 (.D(d3_71__N_561[41]), .CK(osc_clk), .Q(d3[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i41.GSR = "ENABLED";
    FD1S3AX d3_i42 (.D(d3_71__N_561[42]), .CK(osc_clk), .Q(d3[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i42.GSR = "ENABLED";
    FD1S3AX d3_i43 (.D(d3_71__N_561[43]), .CK(osc_clk), .Q(d3[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i43.GSR = "ENABLED";
    FD1S3AX d3_i44 (.D(d3_71__N_561[44]), .CK(osc_clk), .Q(d3[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i44.GSR = "ENABLED";
    FD1S3AX d3_i45 (.D(d3_71__N_561[45]), .CK(osc_clk), .Q(d3[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i45.GSR = "ENABLED";
    FD1S3AX d3_i46 (.D(d3_71__N_561[46]), .CK(osc_clk), .Q(d3[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i46.GSR = "ENABLED";
    FD1S3AX d3_i47 (.D(d3_71__N_561[47]), .CK(osc_clk), .Q(d3[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i47.GSR = "ENABLED";
    FD1S3AX d3_i48 (.D(d3_71__N_561[48]), .CK(osc_clk), .Q(d3[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i48.GSR = "ENABLED";
    FD1S3AX d3_i49 (.D(d3_71__N_561[49]), .CK(osc_clk), .Q(d3[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i49.GSR = "ENABLED";
    FD1S3AX d3_i50 (.D(d3_71__N_561[50]), .CK(osc_clk), .Q(d3[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i50.GSR = "ENABLED";
    FD1S3AX d3_i51 (.D(d3_71__N_561[51]), .CK(osc_clk), .Q(d3[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i51.GSR = "ENABLED";
    FD1S3AX d3_i52 (.D(d3_71__N_561[52]), .CK(osc_clk), .Q(d3[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i52.GSR = "ENABLED";
    FD1S3AX d3_i53 (.D(d3_71__N_561[53]), .CK(osc_clk), .Q(d3[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i53.GSR = "ENABLED";
    FD1S3AX d3_i54 (.D(d3_71__N_561[54]), .CK(osc_clk), .Q(d3[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i54.GSR = "ENABLED";
    FD1S3AX d3_i55 (.D(d3_71__N_561[55]), .CK(osc_clk), .Q(d3[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i55.GSR = "ENABLED";
    FD1S3AX d3_i56 (.D(d3_71__N_561[56]), .CK(osc_clk), .Q(d3[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i56.GSR = "ENABLED";
    FD1S3AX d3_i57 (.D(d3_71__N_561[57]), .CK(osc_clk), .Q(d3[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i57.GSR = "ENABLED";
    FD1S3AX d3_i58 (.D(d3_71__N_561[58]), .CK(osc_clk), .Q(d3[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i58.GSR = "ENABLED";
    FD1S3AX d3_i59 (.D(d3_71__N_561[59]), .CK(osc_clk), .Q(d3[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i59.GSR = "ENABLED";
    FD1S3AX d3_i60 (.D(d3_71__N_561[60]), .CK(osc_clk), .Q(d3[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i60.GSR = "ENABLED";
    FD1S3AX d3_i61 (.D(d3_71__N_561[61]), .CK(osc_clk), .Q(d3[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i61.GSR = "ENABLED";
    FD1S3AX d3_i62 (.D(d3_71__N_561[62]), .CK(osc_clk), .Q(d3[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i62.GSR = "ENABLED";
    FD1S3AX d3_i63 (.D(d3_71__N_561[63]), .CK(osc_clk), .Q(d3[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i63.GSR = "ENABLED";
    FD1S3AX d3_i64 (.D(d3_71__N_561[64]), .CK(osc_clk), .Q(d3[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i64.GSR = "ENABLED";
    FD1S3AX d3_i65 (.D(d3_71__N_561[65]), .CK(osc_clk), .Q(d3[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i65.GSR = "ENABLED";
    FD1S3AX d3_i66 (.D(d3_71__N_561[66]), .CK(osc_clk), .Q(d3[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i66.GSR = "ENABLED";
    FD1S3AX d3_i67 (.D(d3_71__N_561[67]), .CK(osc_clk), .Q(d3[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i67.GSR = "ENABLED";
    FD1S3AX d3_i68 (.D(d3_71__N_561[68]), .CK(osc_clk), .Q(d3[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i68.GSR = "ENABLED";
    FD1S3AX d3_i69 (.D(d3_71__N_561[69]), .CK(osc_clk), .Q(d3[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i69.GSR = "ENABLED";
    FD1S3AX d3_i70 (.D(d3_71__N_561[70]), .CK(osc_clk), .Q(d3[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i70.GSR = "ENABLED";
    FD1S3AX d3_i71 (.D(d3_71__N_561[71]), .CK(osc_clk), .Q(d3[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d3_i71.GSR = "ENABLED";
    FD1S3AX d4_i1 (.D(d4_71__N_633[1]), .CK(osc_clk), .Q(d4[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i1.GSR = "ENABLED";
    FD1S3AX d4_i2 (.D(d4_71__N_633[2]), .CK(osc_clk), .Q(d4[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i2.GSR = "ENABLED";
    FD1S3AX d4_i3 (.D(d4_71__N_633[3]), .CK(osc_clk), .Q(d4[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i3.GSR = "ENABLED";
    FD1S3AX d4_i4 (.D(d4_71__N_633[4]), .CK(osc_clk), .Q(d4[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i4.GSR = "ENABLED";
    FD1S3AX d4_i5 (.D(d4_71__N_633[5]), .CK(osc_clk), .Q(d4[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i5.GSR = "ENABLED";
    FD1S3AX d4_i6 (.D(d4_71__N_633[6]), .CK(osc_clk), .Q(d4[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i6.GSR = "ENABLED";
    FD1S3AX d4_i7 (.D(d4_71__N_633[7]), .CK(osc_clk), .Q(d4[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i7.GSR = "ENABLED";
    FD1S3AX d4_i8 (.D(d4_71__N_633[8]), .CK(osc_clk), .Q(d4[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i8.GSR = "ENABLED";
    FD1S3AX d4_i9 (.D(d4_71__N_633[9]), .CK(osc_clk), .Q(d4[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i9.GSR = "ENABLED";
    FD1S3AX d4_i10 (.D(d4_71__N_633[10]), .CK(osc_clk), .Q(d4[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i10.GSR = "ENABLED";
    FD1S3AX d4_i11 (.D(d4_71__N_633[11]), .CK(osc_clk), .Q(d4[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i11.GSR = "ENABLED";
    FD1S3AX d4_i12 (.D(d4_71__N_633[12]), .CK(osc_clk), .Q(d4[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i12.GSR = "ENABLED";
    FD1S3AX d4_i13 (.D(d4_71__N_633[13]), .CK(osc_clk), .Q(d4[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i13.GSR = "ENABLED";
    FD1S3AX d4_i14 (.D(d4_71__N_633[14]), .CK(osc_clk), .Q(d4[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i14.GSR = "ENABLED";
    FD1S3AX d4_i15 (.D(d4_71__N_633[15]), .CK(osc_clk), .Q(d4[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i15.GSR = "ENABLED";
    FD1S3AX d4_i16 (.D(d4_71__N_633[16]), .CK(osc_clk), .Q(d4[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i16.GSR = "ENABLED";
    FD1S3AX d4_i17 (.D(d4_71__N_633[17]), .CK(osc_clk), .Q(d4[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i17.GSR = "ENABLED";
    FD1S3AX d4_i18 (.D(d4_71__N_633[18]), .CK(osc_clk), .Q(d4[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i18.GSR = "ENABLED";
    FD1S3AX d4_i19 (.D(d4_71__N_633[19]), .CK(osc_clk), .Q(d4[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i19.GSR = "ENABLED";
    FD1S3AX d4_i20 (.D(d4_71__N_633[20]), .CK(osc_clk), .Q(d4[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i20.GSR = "ENABLED";
    FD1S3AX d4_i21 (.D(d4_71__N_633[21]), .CK(osc_clk), .Q(d4[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i21.GSR = "ENABLED";
    FD1S3AX d4_i22 (.D(d4_71__N_633[22]), .CK(osc_clk), .Q(d4[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i22.GSR = "ENABLED";
    FD1S3AX d4_i23 (.D(d4_71__N_633[23]), .CK(osc_clk), .Q(d4[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i23.GSR = "ENABLED";
    FD1S3AX d4_i24 (.D(d4_71__N_633[24]), .CK(osc_clk), .Q(d4[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i24.GSR = "ENABLED";
    FD1S3AX d4_i25 (.D(d4_71__N_633[25]), .CK(osc_clk), .Q(d4[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i25.GSR = "ENABLED";
    FD1S3AX d4_i26 (.D(d4_71__N_633[26]), .CK(osc_clk), .Q(d4[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i26.GSR = "ENABLED";
    FD1S3AX d4_i27 (.D(d4_71__N_633[27]), .CK(osc_clk), .Q(d4[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i27.GSR = "ENABLED";
    FD1S3AX d4_i28 (.D(d4_71__N_633[28]), .CK(osc_clk), .Q(d4[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i28.GSR = "ENABLED";
    FD1S3AX d4_i29 (.D(d4_71__N_633[29]), .CK(osc_clk), .Q(d4[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i29.GSR = "ENABLED";
    FD1S3AX d4_i30 (.D(d4_71__N_633[30]), .CK(osc_clk), .Q(d4[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i30.GSR = "ENABLED";
    FD1S3AX d4_i31 (.D(d4_71__N_633[31]), .CK(osc_clk), .Q(d4[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i31.GSR = "ENABLED";
    FD1S3AX d4_i32 (.D(d4_71__N_633[32]), .CK(osc_clk), .Q(d4[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i32.GSR = "ENABLED";
    FD1S3AX d4_i33 (.D(d4_71__N_633[33]), .CK(osc_clk), .Q(d4[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i33.GSR = "ENABLED";
    FD1S3AX d4_i34 (.D(d4_71__N_633[34]), .CK(osc_clk), .Q(d4[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i34.GSR = "ENABLED";
    FD1S3AX d4_i35 (.D(d4_71__N_633[35]), .CK(osc_clk), .Q(d4[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i35.GSR = "ENABLED";
    FD1S3AX d4_i36 (.D(d4_71__N_633[36]), .CK(osc_clk), .Q(d4[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i36.GSR = "ENABLED";
    FD1S3AX d4_i37 (.D(d4_71__N_633[37]), .CK(osc_clk), .Q(d4[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i37.GSR = "ENABLED";
    FD1S3AX d4_i38 (.D(d4_71__N_633[38]), .CK(osc_clk), .Q(d4[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i38.GSR = "ENABLED";
    FD1S3AX d4_i39 (.D(d4_71__N_633[39]), .CK(osc_clk), .Q(d4[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i39.GSR = "ENABLED";
    FD1S3AX d4_i40 (.D(d4_71__N_633[40]), .CK(osc_clk), .Q(d4[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i40.GSR = "ENABLED";
    FD1S3AX d4_i41 (.D(d4_71__N_633[41]), .CK(osc_clk), .Q(d4[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i41.GSR = "ENABLED";
    FD1S3AX d4_i42 (.D(d4_71__N_633[42]), .CK(osc_clk), .Q(d4[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i42.GSR = "ENABLED";
    FD1S3AX d4_i43 (.D(d4_71__N_633[43]), .CK(osc_clk), .Q(d4[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i43.GSR = "ENABLED";
    FD1S3AX d4_i44 (.D(d4_71__N_633[44]), .CK(osc_clk), .Q(d4[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i44.GSR = "ENABLED";
    FD1S3AX d4_i45 (.D(d4_71__N_633[45]), .CK(osc_clk), .Q(d4[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i45.GSR = "ENABLED";
    FD1S3AX d4_i46 (.D(d4_71__N_633[46]), .CK(osc_clk), .Q(d4[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i46.GSR = "ENABLED";
    FD1S3AX d4_i47 (.D(d4_71__N_633[47]), .CK(osc_clk), .Q(d4[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i47.GSR = "ENABLED";
    FD1S3AX d4_i48 (.D(d4_71__N_633[48]), .CK(osc_clk), .Q(d4[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i48.GSR = "ENABLED";
    FD1S3AX d4_i49 (.D(d4_71__N_633[49]), .CK(osc_clk), .Q(d4[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i49.GSR = "ENABLED";
    FD1S3AX d4_i50 (.D(d4_71__N_633[50]), .CK(osc_clk), .Q(d4[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i50.GSR = "ENABLED";
    FD1S3AX d4_i51 (.D(d4_71__N_633[51]), .CK(osc_clk), .Q(d4[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i51.GSR = "ENABLED";
    FD1S3AX d4_i52 (.D(d4_71__N_633[52]), .CK(osc_clk), .Q(d4[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i52.GSR = "ENABLED";
    FD1S3AX d4_i53 (.D(d4_71__N_633[53]), .CK(osc_clk), .Q(d4[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i53.GSR = "ENABLED";
    FD1S3AX d4_i54 (.D(d4_71__N_633[54]), .CK(osc_clk), .Q(d4[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i54.GSR = "ENABLED";
    FD1S3AX d4_i55 (.D(d4_71__N_633[55]), .CK(osc_clk), .Q(d4[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i55.GSR = "ENABLED";
    FD1S3AX d4_i56 (.D(d4_71__N_633[56]), .CK(osc_clk), .Q(d4[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i56.GSR = "ENABLED";
    FD1S3AX d4_i57 (.D(d4_71__N_633[57]), .CK(osc_clk), .Q(d4[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i57.GSR = "ENABLED";
    FD1S3AX d4_i58 (.D(d4_71__N_633[58]), .CK(osc_clk), .Q(d4[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i58.GSR = "ENABLED";
    FD1S3AX d4_i59 (.D(d4_71__N_633[59]), .CK(osc_clk), .Q(d4[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i59.GSR = "ENABLED";
    FD1S3AX d4_i60 (.D(d4_71__N_633[60]), .CK(osc_clk), .Q(d4[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i60.GSR = "ENABLED";
    FD1S3AX d4_i61 (.D(d4_71__N_633[61]), .CK(osc_clk), .Q(d4[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i61.GSR = "ENABLED";
    FD1S3AX d4_i62 (.D(d4_71__N_633[62]), .CK(osc_clk), .Q(d4[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i62.GSR = "ENABLED";
    FD1S3AX d4_i63 (.D(d4_71__N_633[63]), .CK(osc_clk), .Q(d4[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i63.GSR = "ENABLED";
    FD1S3AX d4_i64 (.D(d4_71__N_633[64]), .CK(osc_clk), .Q(d4[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i64.GSR = "ENABLED";
    FD1S3AX d4_i65 (.D(d4_71__N_633[65]), .CK(osc_clk), .Q(d4[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i65.GSR = "ENABLED";
    FD1S3AX d4_i66 (.D(d4_71__N_633[66]), .CK(osc_clk), .Q(d4[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i66.GSR = "ENABLED";
    FD1S3AX d4_i67 (.D(d4_71__N_633[67]), .CK(osc_clk), .Q(d4[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i67.GSR = "ENABLED";
    FD1S3AX d4_i68 (.D(d4_71__N_633[68]), .CK(osc_clk), .Q(d4[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i68.GSR = "ENABLED";
    FD1S3AX d4_i69 (.D(d4_71__N_633[69]), .CK(osc_clk), .Q(d4[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i69.GSR = "ENABLED";
    FD1S3AX d4_i70 (.D(d4_71__N_633[70]), .CK(osc_clk), .Q(d4[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i70.GSR = "ENABLED";
    FD1S3AX d4_i71 (.D(d4_71__N_633[71]), .CK(osc_clk), .Q(d4[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d4_i71.GSR = "ENABLED";
    FD1S3AX d5_i1 (.D(d5_71__N_705[1]), .CK(osc_clk), .Q(d5[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i1.GSR = "ENABLED";
    FD1S3AX d5_i2 (.D(d5_71__N_705[2]), .CK(osc_clk), .Q(d5[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i2.GSR = "ENABLED";
    FD1S3AX d5_i3 (.D(d5_71__N_705[3]), .CK(osc_clk), .Q(d5[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i3.GSR = "ENABLED";
    FD1S3AX d5_i4 (.D(d5_71__N_705[4]), .CK(osc_clk), .Q(d5[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i4.GSR = "ENABLED";
    FD1S3AX d5_i5 (.D(d5_71__N_705[5]), .CK(osc_clk), .Q(d5[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i5.GSR = "ENABLED";
    FD1S3AX d5_i6 (.D(d5_71__N_705[6]), .CK(osc_clk), .Q(d5[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i6.GSR = "ENABLED";
    FD1S3AX d5_i7 (.D(d5_71__N_705[7]), .CK(osc_clk), .Q(d5[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i7.GSR = "ENABLED";
    FD1S3AX d5_i8 (.D(d5_71__N_705[8]), .CK(osc_clk), .Q(d5[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i8.GSR = "ENABLED";
    FD1S3AX d5_i9 (.D(d5_71__N_705[9]), .CK(osc_clk), .Q(d5[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i9.GSR = "ENABLED";
    FD1S3AX d5_i10 (.D(d5_71__N_705[10]), .CK(osc_clk), .Q(d5[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i10.GSR = "ENABLED";
    FD1S3AX d5_i11 (.D(d5_71__N_705[11]), .CK(osc_clk), .Q(d5[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i11.GSR = "ENABLED";
    FD1S3AX d5_i12 (.D(d5_71__N_705[12]), .CK(osc_clk), .Q(d5[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i12.GSR = "ENABLED";
    FD1S3AX d5_i13 (.D(d5_71__N_705[13]), .CK(osc_clk), .Q(d5[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i13.GSR = "ENABLED";
    FD1S3AX d5_i14 (.D(d5_71__N_705[14]), .CK(osc_clk), .Q(d5[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i14.GSR = "ENABLED";
    FD1S3AX d5_i15 (.D(d5_71__N_705[15]), .CK(osc_clk), .Q(d5[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i15.GSR = "ENABLED";
    FD1S3AX d5_i16 (.D(d5_71__N_705[16]), .CK(osc_clk), .Q(d5[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i16.GSR = "ENABLED";
    FD1S3AX d5_i17 (.D(d5_71__N_705[17]), .CK(osc_clk), .Q(d5[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i17.GSR = "ENABLED";
    FD1S3AX d5_i18 (.D(d5_71__N_705[18]), .CK(osc_clk), .Q(d5[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i18.GSR = "ENABLED";
    FD1S3AX d5_i19 (.D(d5_71__N_705[19]), .CK(osc_clk), .Q(d5[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i19.GSR = "ENABLED";
    FD1S3AX d5_i20 (.D(d5_71__N_705[20]), .CK(osc_clk), .Q(d5[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i20.GSR = "ENABLED";
    FD1S3AX d5_i21 (.D(d5_71__N_705[21]), .CK(osc_clk), .Q(d5[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i21.GSR = "ENABLED";
    FD1S3AX d5_i22 (.D(d5_71__N_705[22]), .CK(osc_clk), .Q(d5[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i22.GSR = "ENABLED";
    FD1S3AX d5_i23 (.D(d5_71__N_705[23]), .CK(osc_clk), .Q(d5[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i23.GSR = "ENABLED";
    FD1S3AX d5_i24 (.D(d5_71__N_705[24]), .CK(osc_clk), .Q(d5[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i24.GSR = "ENABLED";
    FD1S3AX d5_i25 (.D(d5_71__N_705[25]), .CK(osc_clk), .Q(d5[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i25.GSR = "ENABLED";
    FD1S3AX d5_i26 (.D(d5_71__N_705[26]), .CK(osc_clk), .Q(d5[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i26.GSR = "ENABLED";
    FD1S3AX d5_i27 (.D(d5_71__N_705[27]), .CK(osc_clk), .Q(d5[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i27.GSR = "ENABLED";
    FD1S3AX d5_i28 (.D(d5_71__N_705[28]), .CK(osc_clk), .Q(d5[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i28.GSR = "ENABLED";
    FD1S3AX d5_i29 (.D(d5_71__N_705[29]), .CK(osc_clk), .Q(d5[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i29.GSR = "ENABLED";
    FD1S3AX d5_i30 (.D(d5_71__N_705[30]), .CK(osc_clk), .Q(d5[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i30.GSR = "ENABLED";
    FD1S3AX d5_i31 (.D(d5_71__N_705[31]), .CK(osc_clk), .Q(d5[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i31.GSR = "ENABLED";
    FD1S3AX d5_i32 (.D(d5_71__N_705[32]), .CK(osc_clk), .Q(d5[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i32.GSR = "ENABLED";
    FD1S3AX d5_i33 (.D(d5_71__N_705[33]), .CK(osc_clk), .Q(d5[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i33.GSR = "ENABLED";
    FD1S3AX d5_i34 (.D(d5_71__N_705[34]), .CK(osc_clk), .Q(d5[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i34.GSR = "ENABLED";
    FD1S3AX d5_i35 (.D(d5_71__N_705[35]), .CK(osc_clk), .Q(d5[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i35.GSR = "ENABLED";
    FD1S3AX d5_i36 (.D(d5_71__N_705[36]), .CK(osc_clk), .Q(d5[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i36.GSR = "ENABLED";
    FD1S3AX d5_i37 (.D(d5_71__N_705[37]), .CK(osc_clk), .Q(d5[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i37.GSR = "ENABLED";
    FD1S3AX d5_i38 (.D(d5_71__N_705[38]), .CK(osc_clk), .Q(d5[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i38.GSR = "ENABLED";
    FD1S3AX d5_i39 (.D(d5_71__N_705[39]), .CK(osc_clk), .Q(d5[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i39.GSR = "ENABLED";
    FD1S3AX d5_i40 (.D(d5_71__N_705[40]), .CK(osc_clk), .Q(d5[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i40.GSR = "ENABLED";
    FD1S3AX d5_i41 (.D(d5_71__N_705[41]), .CK(osc_clk), .Q(d5[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i41.GSR = "ENABLED";
    FD1S3AX d5_i42 (.D(d5_71__N_705[42]), .CK(osc_clk), .Q(d5[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i42.GSR = "ENABLED";
    FD1S3AX d5_i43 (.D(d5_71__N_705[43]), .CK(osc_clk), .Q(d5[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i43.GSR = "ENABLED";
    FD1S3AX d5_i44 (.D(d5_71__N_705[44]), .CK(osc_clk), .Q(d5[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i44.GSR = "ENABLED";
    FD1S3AX d5_i45 (.D(d5_71__N_705[45]), .CK(osc_clk), .Q(d5[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i45.GSR = "ENABLED";
    FD1S3AX d5_i46 (.D(d5_71__N_705[46]), .CK(osc_clk), .Q(d5[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i46.GSR = "ENABLED";
    FD1S3AX d5_i47 (.D(d5_71__N_705[47]), .CK(osc_clk), .Q(d5[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i47.GSR = "ENABLED";
    FD1S3AX d5_i48 (.D(d5_71__N_705[48]), .CK(osc_clk), .Q(d5[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i48.GSR = "ENABLED";
    FD1S3AX d5_i49 (.D(d5_71__N_705[49]), .CK(osc_clk), .Q(d5[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i49.GSR = "ENABLED";
    FD1S3AX d5_i50 (.D(d5_71__N_705[50]), .CK(osc_clk), .Q(d5[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i50.GSR = "ENABLED";
    FD1S3AX d5_i51 (.D(d5_71__N_705[51]), .CK(osc_clk), .Q(d5[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i51.GSR = "ENABLED";
    FD1S3AX d5_i52 (.D(d5_71__N_705[52]), .CK(osc_clk), .Q(d5[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i52.GSR = "ENABLED";
    FD1S3AX d5_i53 (.D(d5_71__N_705[53]), .CK(osc_clk), .Q(d5[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i53.GSR = "ENABLED";
    FD1S3AX d5_i54 (.D(d5_71__N_705[54]), .CK(osc_clk), .Q(d5[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i54.GSR = "ENABLED";
    FD1S3AX d5_i55 (.D(d5_71__N_705[55]), .CK(osc_clk), .Q(d5[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i55.GSR = "ENABLED";
    FD1S3AX d5_i56 (.D(d5_71__N_705[56]), .CK(osc_clk), .Q(d5[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i56.GSR = "ENABLED";
    FD1S3AX d5_i57 (.D(d5_71__N_705[57]), .CK(osc_clk), .Q(d5[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i57.GSR = "ENABLED";
    FD1S3AX d5_i58 (.D(d5_71__N_705[58]), .CK(osc_clk), .Q(d5[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i58.GSR = "ENABLED";
    FD1S3AX d5_i59 (.D(d5_71__N_705[59]), .CK(osc_clk), .Q(d5[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i59.GSR = "ENABLED";
    FD1S3AX d5_i60 (.D(d5_71__N_705[60]), .CK(osc_clk), .Q(d5[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i60.GSR = "ENABLED";
    FD1S3AX d5_i61 (.D(d5_71__N_705[61]), .CK(osc_clk), .Q(d5[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i61.GSR = "ENABLED";
    FD1S3AX d5_i62 (.D(d5_71__N_705[62]), .CK(osc_clk), .Q(d5[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i62.GSR = "ENABLED";
    FD1S3AX d5_i63 (.D(d5_71__N_705[63]), .CK(osc_clk), .Q(d5[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i63.GSR = "ENABLED";
    FD1S3AX d5_i64 (.D(d5_71__N_705[64]), .CK(osc_clk), .Q(d5[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i64.GSR = "ENABLED";
    FD1S3AX d5_i65 (.D(d5_71__N_705[65]), .CK(osc_clk), .Q(d5[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i65.GSR = "ENABLED";
    FD1S3AX d5_i66 (.D(d5_71__N_705[66]), .CK(osc_clk), .Q(d5[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i66.GSR = "ENABLED";
    FD1S3AX d5_i67 (.D(d5_71__N_705[67]), .CK(osc_clk), .Q(d5[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i67.GSR = "ENABLED";
    FD1S3AX d5_i68 (.D(d5_71__N_705[68]), .CK(osc_clk), .Q(d5[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i68.GSR = "ENABLED";
    FD1S3AX d5_i69 (.D(d5_71__N_705[69]), .CK(osc_clk), .Q(d5[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i69.GSR = "ENABLED";
    FD1S3AX d5_i70 (.D(d5_71__N_705[70]), .CK(osc_clk), .Q(d5[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i70.GSR = "ENABLED";
    FD1S3AX d5_i71 (.D(d5_71__N_705[71]), .CK(osc_clk), .Q(d5[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d5_i71.GSR = "ENABLED";
    FD1P3AX d6_i0_i1 (.D(d6_71__N_1458[1]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d6_i0_i2 (.D(d6_71__N_1458[2]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d6_i0_i3 (.D(d6_71__N_1458[3]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d6_i0_i4 (.D(d6_71__N_1458[4]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d6_i0_i5 (.D(d6_71__N_1458[5]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d6_i0_i6 (.D(d6_71__N_1458[6]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d6_i0_i7 (.D(d6_71__N_1458[7]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d6_i0_i8 (.D(d6_71__N_1458[8]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d6_i0_i9 (.D(d6_71__N_1458[9]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d6_i0_i10 (.D(d6_71__N_1458[10]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d6_i0_i11 (.D(d6_71__N_1458[11]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d6_i0_i12 (.D(d6_71__N_1458[12]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d6_i0_i13 (.D(d6_71__N_1458[13]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d6_i0_i14 (.D(d6_71__N_1458[14]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d6_i0_i15 (.D(d6_71__N_1458[15]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d6_i0_i16 (.D(d6_71__N_1458[16]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d6_i0_i17 (.D(d6_71__N_1458[17]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d6_i0_i18 (.D(d6_71__N_1458[18]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d6_i0_i19 (.D(d6_71__N_1458[19]), .SP(osc_clk_enable_833), .CK(osc_clk), 
            .Q(d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d6_i0_i20 (.D(d6_71__N_1458[20]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d6_i0_i21 (.D(d6_71__N_1458[21]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d6_i0_i22 (.D(d6_71__N_1458[22]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d6_i0_i23 (.D(d6_71__N_1458[23]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d6_i0_i24 (.D(d6_71__N_1458[24]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d6_i0_i25 (.D(d6_71__N_1458[25]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d6_i0_i26 (.D(d6_71__N_1458[26]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d6_i0_i27 (.D(d6_71__N_1458[27]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d6_i0_i28 (.D(d6_71__N_1458[28]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d6_i0_i29 (.D(d6_71__N_1458[29]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d6_i0_i30 (.D(d6_71__N_1458[30]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d6_i0_i31 (.D(d6_71__N_1458[31]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d6_i0_i32 (.D(d6_71__N_1458[32]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d6_i0_i33 (.D(d6_71__N_1458[33]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d6_i0_i34 (.D(d6_71__N_1458[34]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d6_i0_i35 (.D(d6_71__N_1458[35]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d6_i0_i36 (.D(d6_71__N_1458[36]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d6_i0_i37 (.D(d6_71__N_1458[37]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d6_i0_i38 (.D(d6_71__N_1458[38]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d6_i0_i39 (.D(d6_71__N_1458[39]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d6_i0_i40 (.D(d6_71__N_1458[40]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d6_i0_i41 (.D(d6_71__N_1458[41]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d6_i0_i42 (.D(d6_71__N_1458[42]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d6_i0_i43 (.D(d6_71__N_1458[43]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d6_i0_i44 (.D(d6_71__N_1458[44]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d6_i0_i45 (.D(d6_71__N_1458[45]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d6_i0_i46 (.D(d6_71__N_1458[46]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d6_i0_i47 (.D(d6_71__N_1458[47]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d6_i0_i48 (.D(d6_71__N_1458[48]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d6_i0_i49 (.D(d6_71__N_1458[49]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d6_i0_i50 (.D(d6_71__N_1458[50]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d6_i0_i51 (.D(d6_71__N_1458[51]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d6_i0_i52 (.D(d6_71__N_1458[52]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d6_i0_i53 (.D(d6_71__N_1458[53]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d6_i0_i54 (.D(d6_71__N_1458[54]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d6_i0_i55 (.D(d6_71__N_1458[55]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d6_i0_i56 (.D(d6_71__N_1458[56]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d6_i0_i57 (.D(d6_71__N_1458[57]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d6_i0_i58 (.D(d6_71__N_1458[58]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d6_i0_i59 (.D(d6_71__N_1458[59]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d6_i0_i60 (.D(d6_71__N_1458[60]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d6_i0_i61 (.D(d6_71__N_1458[61]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d6_i0_i62 (.D(d6_71__N_1458[62]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d6_i0_i63 (.D(d6_71__N_1458[63]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d6_i0_i64 (.D(d6_71__N_1458[64]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d6_i0_i65 (.D(d6_71__N_1458[65]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d6_i0_i66 (.D(d6_71__N_1458[66]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d6_i0_i67 (.D(d6_71__N_1458[67]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d6_i0_i68 (.D(d6_71__N_1458[68]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d6_i0_i69 (.D(d6_71__N_1458[69]), .SP(osc_clk_enable_883), .CK(osc_clk), 
            .Q(d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d6_i0_i70 (.D(d6_71__N_1458[70]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d6_i0_i71 (.D(d6_71__N_1458[71]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i1 (.D(d6[1]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i2 (.D(d6[2]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i3 (.D(d6[3]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i4 (.D(d6[4]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i5 (.D(d6[5]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i6 (.D(d6[6]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i7 (.D(d6[7]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i8 (.D(d6[8]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i9 (.D(d6[9]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i10 (.D(d6[10]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i11 (.D(d6[11]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i12 (.D(d6[12]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i13 (.D(d6[13]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i14 (.D(d6[14]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i15 (.D(d6[15]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i16 (.D(d6[16]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i17 (.D(d6[17]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i18 (.D(d6[18]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i19 (.D(d6[19]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i20 (.D(d6[20]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i21 (.D(d6[21]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i22 (.D(d6[22]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i23 (.D(d6[23]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i24 (.D(d6[24]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i25 (.D(d6[25]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i26 (.D(d6[26]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i27 (.D(d6[27]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i28 (.D(d6[28]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i29 (.D(d6[29]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i30 (.D(d6[30]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i31 (.D(d6[31]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i32 (.D(d6[32]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i33 (.D(d6[33]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i34 (.D(d6[34]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i35 (.D(d6[35]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i36 (.D(d6[36]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i37 (.D(d6[37]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i38 (.D(d6[38]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i39 (.D(d6[39]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i40 (.D(d6[40]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i41 (.D(d6[41]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i42 (.D(d6[42]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i43 (.D(d6[43]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i44 (.D(d6[44]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i45 (.D(d6[45]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i46 (.D(d6[46]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i47 (.D(d6[47]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i48 (.D(d6[48]), .SP(osc_clk_enable_933), .CK(osc_clk), 
            .Q(d_d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i49 (.D(d6[49]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d_d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i50 (.D(d6[50]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d_d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i51 (.D(d6[51]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d_d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i52 (.D(d6[52]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d_d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i53 (.D(d6[53]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d_d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i54 (.D(d6[54]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d_d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i55 (.D(d6[55]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d_d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i56 (.D(d6[56]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d_d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i57 (.D(d6[57]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d_d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i58 (.D(d6[58]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d_d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i59 (.D(d6[59]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d_d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i60 (.D(d6[60]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d_d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i61 (.D(d6[61]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d_d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i62 (.D(d6[62]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d_d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i63 (.D(d6[63]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d_d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i64 (.D(d6[64]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d_d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i65 (.D(d6[65]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d_d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i66 (.D(d6[66]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d_d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i67 (.D(d6[67]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d_d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i68 (.D(d6[68]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d_d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i69 (.D(d6[69]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d_d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i70 (.D(d6[70]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d_d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i71 (.D(d6[71]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d_d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d7_i0_i1 (.D(d7_71__N_1530[1]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d7_i0_i2 (.D(d7_71__N_1530[2]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d7_i0_i3 (.D(d7_71__N_1530[3]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d7_i0_i4 (.D(d7_71__N_1530[4]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d7_i0_i5 (.D(d7_71__N_1530[5]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d7_i0_i6 (.D(d7_71__N_1530[6]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d7_i0_i7 (.D(d7_71__N_1530[7]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d7_i0_i8 (.D(d7_71__N_1530[8]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d7_i0_i9 (.D(d7_71__N_1530[9]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d7_i0_i10 (.D(d7_71__N_1530[10]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d7_i0_i11 (.D(d7_71__N_1530[11]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d7_i0_i12 (.D(d7_71__N_1530[12]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d7_i0_i13 (.D(d7_71__N_1530[13]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d7_i0_i14 (.D(d7_71__N_1530[14]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d7_i0_i15 (.D(d7_71__N_1530[15]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d7_i0_i16 (.D(d7_71__N_1530[16]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d7_i0_i17 (.D(d7_71__N_1530[17]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d7_i0_i18 (.D(d7_71__N_1530[18]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d7_i0_i19 (.D(d7_71__N_1530[19]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d7_i0_i20 (.D(d7_71__N_1530[20]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d7_i0_i21 (.D(d7_71__N_1530[21]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d7_i0_i22 (.D(d7_71__N_1530[22]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d7_i0_i23 (.D(d7_71__N_1530[23]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d7_i0_i24 (.D(d7_71__N_1530[24]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d7_i0_i25 (.D(d7_71__N_1530[25]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d7_i0_i26 (.D(d7_71__N_1530[26]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d7_i0_i27 (.D(d7_71__N_1530[27]), .SP(osc_clk_enable_983), .CK(osc_clk), 
            .Q(d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d7_i0_i28 (.D(d7_71__N_1530[28]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d7_i0_i29 (.D(d7_71__N_1530[29]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d7_i0_i30 (.D(d7_71__N_1530[30]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d7_i0_i31 (.D(d7_71__N_1530[31]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d7_i0_i32 (.D(d7_71__N_1530[32]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d7_i0_i33 (.D(d7_71__N_1530[33]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d7_i0_i34 (.D(d7_71__N_1530[34]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d7_i0_i35 (.D(d7_71__N_1530[35]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d7_i0_i36 (.D(d7_71__N_1530[36]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d7_i0_i37 (.D(d7_71__N_1530[37]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d7_i0_i38 (.D(d7_71__N_1530[38]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d7_i0_i39 (.D(d7_71__N_1530[39]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d7_i0_i40 (.D(d7_71__N_1530[40]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d7_i0_i41 (.D(d7_71__N_1530[41]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d7_i0_i42 (.D(d7_71__N_1530[42]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d7_i0_i43 (.D(d7_71__N_1530[43]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d7_i0_i44 (.D(d7_71__N_1530[44]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d7_i0_i45 (.D(d7_71__N_1530[45]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d7_i0_i46 (.D(d7_71__N_1530[46]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d7_i0_i47 (.D(d7_71__N_1530[47]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d7_i0_i48 (.D(d7_71__N_1530[48]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d7_i0_i49 (.D(d7_71__N_1530[49]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d7_i0_i50 (.D(d7_71__N_1530[50]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d7_i0_i51 (.D(d7_71__N_1530[51]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d7_i0_i52 (.D(d7_71__N_1530[52]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d7_i0_i53 (.D(d7_71__N_1530[53]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d7_i0_i54 (.D(d7_71__N_1530[54]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d7_i0_i55 (.D(d7_71__N_1530[55]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d7_i0_i56 (.D(d7_71__N_1530[56]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d7_i0_i57 (.D(d7_71__N_1530[57]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d7_i0_i58 (.D(d7_71__N_1530[58]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d7_i0_i59 (.D(d7_71__N_1530[59]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d7_i0_i60 (.D(d7_71__N_1530[60]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d7_i0_i61 (.D(d7_71__N_1530[61]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d7_i0_i62 (.D(d7_71__N_1530[62]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d7_i0_i63 (.D(d7_71__N_1530[63]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d7_i0_i64 (.D(d7_71__N_1530[64]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d7_i0_i65 (.D(d7_71__N_1530[65]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d7_i0_i66 (.D(d7_71__N_1530[66]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d7_i0_i67 (.D(d7_71__N_1530[67]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d7_i0_i68 (.D(d7_71__N_1530[68]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d7_i0_i69 (.D(d7_71__N_1530[69]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d7_i0_i70 (.D(d7_71__N_1530[70]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d7_i0_i71 (.D(d7_71__N_1530[71]), .SP(osc_clk_enable_1033), 
            .CK(osc_clk), .Q(d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i1 (.D(d7[1]), .SP(osc_clk_enable_1033), .CK(osc_clk), 
            .Q(d_d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i2 (.D(d7[2]), .SP(osc_clk_enable_1033), .CK(osc_clk), 
            .Q(d_d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i3 (.D(d7[3]), .SP(osc_clk_enable_1033), .CK(osc_clk), 
            .Q(d_d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i4 (.D(d7[4]), .SP(osc_clk_enable_1033), .CK(osc_clk), 
            .Q(d_d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i5 (.D(d7[5]), .SP(osc_clk_enable_1033), .CK(osc_clk), 
            .Q(d_d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i6 (.D(d7[6]), .SP(osc_clk_enable_1033), .CK(osc_clk), 
            .Q(d_d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i7 (.D(d7[7]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i8 (.D(d7[8]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i9 (.D(d7[9]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i10 (.D(d7[10]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i11 (.D(d7[11]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i12 (.D(d7[12]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i13 (.D(d7[13]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i14 (.D(d7[14]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i15 (.D(d7[15]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i16 (.D(d7[16]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i17 (.D(d7[17]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i18 (.D(d7[18]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i19 (.D(d7[19]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i20 (.D(d7[20]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i21 (.D(d7[21]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i22 (.D(d7[22]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i23 (.D(d7[23]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i24 (.D(d7[24]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i25 (.D(d7[25]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i26 (.D(d7[26]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i27 (.D(d7[27]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i28 (.D(d7[28]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i29 (.D(d7[29]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i30 (.D(d7[30]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i31 (.D(d7[31]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i32 (.D(d7[32]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i33 (.D(d7[33]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i34 (.D(d7[34]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i35 (.D(d7[35]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i36 (.D(d7[36]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i37 (.D(d7[37]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i38 (.D(d7[38]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i39 (.D(d7[39]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i40 (.D(d7[40]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i41 (.D(d7[41]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i42 (.D(d7[42]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i43 (.D(d7[43]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i44 (.D(d7[44]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i45 (.D(d7[45]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i46 (.D(d7[46]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i47 (.D(d7[47]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i48 (.D(d7[48]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i49 (.D(d7[49]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i50 (.D(d7[50]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i51 (.D(d7[51]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i52 (.D(d7[52]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i53 (.D(d7[53]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i54 (.D(d7[54]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i55 (.D(d7[55]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i56 (.D(d7[56]), .SP(osc_clk_enable_1083), .CK(osc_clk), 
            .Q(d_d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i57 (.D(d7[57]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d_d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i58 (.D(d7[58]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d_d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i59 (.D(d7[59]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d_d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i60 (.D(d7[60]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d_d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i61 (.D(d7[61]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d_d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i62 (.D(d7[62]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d_d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i63 (.D(d7[63]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d_d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i64 (.D(d7[64]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d_d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i65 (.D(d7[65]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d_d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i66 (.D(d7[66]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d_d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i67 (.D(d7[67]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d_d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i68 (.D(d7[68]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d_d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i69 (.D(d7[69]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d_d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i70 (.D(d7[70]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d_d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i71 (.D(d7[71]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d_d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d8_i0_i1 (.D(d8_71__N_1602[1]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d8_i0_i2 (.D(d8_71__N_1602[2]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d8_i0_i3 (.D(d8_71__N_1602[3]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d8_i0_i4 (.D(d8_71__N_1602[4]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d8_i0_i5 (.D(d8_71__N_1602[5]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d8_i0_i6 (.D(d8_71__N_1602[6]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d8_i0_i7 (.D(d8_71__N_1602[7]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d8_i0_i8 (.D(d8_71__N_1602[8]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d8_i0_i9 (.D(d8_71__N_1602[9]), .SP(osc_clk_enable_1133), .CK(osc_clk), 
            .Q(d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d8_i0_i10 (.D(d8_71__N_1602[10]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d8_i0_i11 (.D(d8_71__N_1602[11]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d8_i0_i12 (.D(d8_71__N_1602[12]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d8_i0_i13 (.D(d8_71__N_1602[13]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d8_i0_i14 (.D(d8_71__N_1602[14]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d8_i0_i15 (.D(d8_71__N_1602[15]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d8_i0_i16 (.D(d8_71__N_1602[16]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d8_i0_i17 (.D(d8_71__N_1602[17]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d8_i0_i18 (.D(d8_71__N_1602[18]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d8_i0_i19 (.D(d8_71__N_1602[19]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d8_i0_i20 (.D(d8_71__N_1602[20]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d8_i0_i21 (.D(d8_71__N_1602[21]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d8_i0_i22 (.D(d8_71__N_1602[22]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d8_i0_i23 (.D(d8_71__N_1602[23]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d8_i0_i24 (.D(d8_71__N_1602[24]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d8_i0_i25 (.D(d8_71__N_1602[25]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d8_i0_i26 (.D(d8_71__N_1602[26]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d8_i0_i27 (.D(d8_71__N_1602[27]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d8_i0_i28 (.D(d8_71__N_1602[28]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d8_i0_i29 (.D(d8_71__N_1602[29]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d8_i0_i30 (.D(d8_71__N_1602[30]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d8_i0_i31 (.D(d8_71__N_1602[31]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d8_i0_i32 (.D(d8_71__N_1602[32]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d8_i0_i33 (.D(d8_71__N_1602[33]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d8_i0_i34 (.D(d8_71__N_1602[34]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d8_i0_i35 (.D(d8_71__N_1602[35]), .SP(osc_clk_enable_1133), 
            .CK(osc_clk), .Q(d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d8_i0_i36 (.D(d8_71__N_1602[36]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d8_i0_i37 (.D(d8_71__N_1602[37]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d8_i0_i38 (.D(d8_71__N_1602[38]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d8_i0_i39 (.D(d8_71__N_1602[39]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d8_i0_i40 (.D(d8_71__N_1602[40]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d8_i0_i41 (.D(d8_71__N_1602[41]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d8_i0_i42 (.D(d8_71__N_1602[42]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d8_i0_i43 (.D(d8_71__N_1602[43]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d8_i0_i44 (.D(d8_71__N_1602[44]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d8_i0_i45 (.D(d8_71__N_1602[45]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d8_i0_i46 (.D(d8_71__N_1602[46]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d8_i0_i47 (.D(d8_71__N_1602[47]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d8_i0_i48 (.D(d8_71__N_1602[48]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d8_i0_i49 (.D(d8_71__N_1602[49]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d8_i0_i50 (.D(d8_71__N_1602[50]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d8_i0_i51 (.D(d8_71__N_1602[51]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d8_i0_i52 (.D(d8_71__N_1602[52]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d8_i0_i53 (.D(d8_71__N_1602[53]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d8_i0_i54 (.D(d8_71__N_1602[54]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d8_i0_i55 (.D(d8_71__N_1602[55]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d8_i0_i56 (.D(d8_71__N_1602[56]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d8_i0_i57 (.D(d8_71__N_1602[57]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d8_i0_i58 (.D(d8_71__N_1602[58]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d8_i0_i59 (.D(d8_71__N_1602[59]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d8_i0_i60 (.D(d8_71__N_1602[60]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d8_i0_i61 (.D(d8_71__N_1602[61]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d8_i0_i62 (.D(d8_71__N_1602[62]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d8_i0_i63 (.D(d8_71__N_1602[63]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d8_i0_i64 (.D(d8_71__N_1602[64]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d8_i0_i65 (.D(d8_71__N_1602[65]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d8_i0_i66 (.D(d8_71__N_1602[66]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d8_i0_i67 (.D(d8_71__N_1602[67]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d8_i0_i68 (.D(d8_71__N_1602[68]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d8_i0_i69 (.D(d8_71__N_1602[69]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d8_i0_i70 (.D(d8_71__N_1602[70]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d8_i0_i71 (.D(d8_71__N_1602[71]), .SP(osc_clk_enable_1183), 
            .CK(osc_clk), .Q(d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i1 (.D(d8[1]), .SP(osc_clk_enable_1183), .CK(osc_clk), 
            .Q(d_d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i2 (.D(d8[2]), .SP(osc_clk_enable_1183), .CK(osc_clk), 
            .Q(d_d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i3 (.D(d8[3]), .SP(osc_clk_enable_1183), .CK(osc_clk), 
            .Q(d_d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i4 (.D(d8[4]), .SP(osc_clk_enable_1183), .CK(osc_clk), 
            .Q(d_d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i5 (.D(d8[5]), .SP(osc_clk_enable_1183), .CK(osc_clk), 
            .Q(d_d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i6 (.D(d8[6]), .SP(osc_clk_enable_1183), .CK(osc_clk), 
            .Q(d_d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i7 (.D(d8[7]), .SP(osc_clk_enable_1183), .CK(osc_clk), 
            .Q(d_d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i8 (.D(d8[8]), .SP(osc_clk_enable_1183), .CK(osc_clk), 
            .Q(d_d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i9 (.D(d8[9]), .SP(osc_clk_enable_1183), .CK(osc_clk), 
            .Q(d_d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i10 (.D(d8[10]), .SP(osc_clk_enable_1183), .CK(osc_clk), 
            .Q(d_d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i11 (.D(d8[11]), .SP(osc_clk_enable_1183), .CK(osc_clk), 
            .Q(d_d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i12 (.D(d8[12]), .SP(osc_clk_enable_1183), .CK(osc_clk), 
            .Q(d_d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i13 (.D(d8[13]), .SP(osc_clk_enable_1183), .CK(osc_clk), 
            .Q(d_d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i14 (.D(d8[14]), .SP(osc_clk_enable_1183), .CK(osc_clk), 
            .Q(d_d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i15 (.D(d8[15]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i16 (.D(d8[16]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i17 (.D(d8[17]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i18 (.D(d8[18]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i19 (.D(d8[19]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i20 (.D(d8[20]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i21 (.D(d8[21]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i22 (.D(d8[22]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i23 (.D(d8[23]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i24 (.D(d8[24]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i25 (.D(d8[25]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i26 (.D(d8[26]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i27 (.D(d8[27]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i28 (.D(d8[28]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i29 (.D(d8[29]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i30 (.D(d8[30]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i31 (.D(d8[31]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i32 (.D(d8[32]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i33 (.D(d8[33]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i34 (.D(d8[34]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i35 (.D(d8[35]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i36 (.D(d8[36]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i37 (.D(d8[37]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i38 (.D(d8[38]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i39 (.D(d8[39]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i40 (.D(d8[40]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i41 (.D(d8[41]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i42 (.D(d8[42]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i43 (.D(d8[43]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i44 (.D(d8[44]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i45 (.D(d8[45]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i46 (.D(d8[46]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i47 (.D(d8[47]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i48 (.D(d8[48]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i49 (.D(d8[49]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i50 (.D(d8[50]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i51 (.D(d8[51]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i52 (.D(d8[52]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i53 (.D(d8[53]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i54 (.D(d8[54]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i55 (.D(d8[55]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i56 (.D(d8[56]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i57 (.D(d8[57]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i58 (.D(d8[58]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i59 (.D(d8[59]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i60 (.D(d8[60]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i61 (.D(d8[61]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i62 (.D(d8[62]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i63 (.D(d8[63]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i64 (.D(d8[64]), .SP(osc_clk_enable_1233), .CK(osc_clk), 
            .Q(d_d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i65 (.D(d8[65]), .SP(osc_clk_enable_1283), .CK(osc_clk), 
            .Q(d_d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i66 (.D(d8[66]), .SP(osc_clk_enable_1283), .CK(osc_clk), 
            .Q(d_d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i67 (.D(d8[67]), .SP(osc_clk_enable_1283), .CK(osc_clk), 
            .Q(d_d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i68 (.D(d8[68]), .SP(osc_clk_enable_1283), .CK(osc_clk), 
            .Q(d_d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i69 (.D(d8[69]), .SP(osc_clk_enable_1283), .CK(osc_clk), 
            .Q(d_d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i70 (.D(d8[70]), .SP(osc_clk_enable_1283), .CK(osc_clk), 
            .Q(d_d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i71 (.D(d8[71]), .SP(osc_clk_enable_1283), .CK(osc_clk), 
            .Q(d_d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d9_i0_i1 (.D(d9_71__N_1674[1]), .SP(osc_clk_enable_1283), .CK(osc_clk), 
            .Q(d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d9_i0_i2 (.D(d9_71__N_1674[2]), .SP(osc_clk_enable_1283), .CK(osc_clk), 
            .Q(d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d9_i0_i3 (.D(d9_71__N_1674[3]), .SP(osc_clk_enable_1283), .CK(osc_clk), 
            .Q(d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d9_i0_i4 (.D(d9_71__N_1674[4]), .SP(osc_clk_enable_1283), .CK(osc_clk), 
            .Q(d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d9_i0_i5 (.D(d9_71__N_1674[5]), .SP(osc_clk_enable_1283), .CK(osc_clk), 
            .Q(d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d9_i0_i6 (.D(d9_71__N_1674[6]), .SP(osc_clk_enable_1283), .CK(osc_clk), 
            .Q(d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d9_i0_i7 (.D(d9_71__N_1674[7]), .SP(osc_clk_enable_1283), .CK(osc_clk), 
            .Q(d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d9_i0_i8 (.D(d9_71__N_1674[8]), .SP(osc_clk_enable_1283), .CK(osc_clk), 
            .Q(d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d9_i0_i9 (.D(d9_71__N_1674[9]), .SP(osc_clk_enable_1283), .CK(osc_clk), 
            .Q(d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d9_i0_i10 (.D(d9_71__N_1674[10]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d9_i0_i11 (.D(d9_71__N_1674[11]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d9_i0_i12 (.D(d9_71__N_1674[12]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d9_i0_i13 (.D(d9_71__N_1674[13]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d9_i0_i14 (.D(d9_71__N_1674[14]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d9_i0_i15 (.D(d9_71__N_1674[15]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d9_i0_i16 (.D(d9_71__N_1674[16]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d9_i0_i17 (.D(d9_71__N_1674[17]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d9_i0_i18 (.D(d9_71__N_1674[18]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d9_i0_i19 (.D(d9_71__N_1674[19]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d9_i0_i20 (.D(d9_71__N_1674[20]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d9_i0_i21 (.D(d9_71__N_1674[21]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d9_i0_i22 (.D(d9_71__N_1674[22]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d9_i0_i23 (.D(d9_71__N_1674[23]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d9_i0_i24 (.D(d9_71__N_1674[24]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d9_i0_i25 (.D(d9_71__N_1674[25]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d9_i0_i26 (.D(d9_71__N_1674[26]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d9_i0_i27 (.D(d9_71__N_1674[27]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d9_i0_i28 (.D(d9_71__N_1674[28]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d9_i0_i29 (.D(d9_71__N_1674[29]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d9_i0_i30 (.D(d9_71__N_1674[30]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d9_i0_i31 (.D(d9_71__N_1674[31]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d9_i0_i32 (.D(d9_71__N_1674[32]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d9_i0_i33 (.D(d9_71__N_1674[33]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d9_i0_i34 (.D(d9_71__N_1674[34]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d9_i0_i35 (.D(d9_71__N_1674[35]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d9_i0_i36 (.D(d9_71__N_1674[36]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d9_i0_i37 (.D(d9_71__N_1674[37]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d9_i0_i38 (.D(d9_71__N_1674[38]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d9_i0_i39 (.D(d9_71__N_1674[39]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d9_i0_i40 (.D(d9_71__N_1674[40]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d9_i0_i41 (.D(d9_71__N_1674[41]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d9_i0_i42 (.D(d9_71__N_1674[42]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d9_i0_i43 (.D(d9_71__N_1674[43]), .SP(osc_clk_enable_1283), 
            .CK(osc_clk), .Q(d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d9_i0_i44 (.D(d9_71__N_1674[44]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d9_i0_i45 (.D(d9_71__N_1674[45]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d9_i0_i46 (.D(d9_71__N_1674[46]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d9_i0_i47 (.D(d9_71__N_1674[47]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d9_i0_i48 (.D(d9_71__N_1674[48]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d9_i0_i49 (.D(d9_71__N_1674[49]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d9_i0_i50 (.D(d9_71__N_1674[50]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d9_i0_i51 (.D(d9_71__N_1674[51]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d9_i0_i52 (.D(d9_71__N_1674[52]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d9_i0_i53 (.D(d9_71__N_1674[53]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d9_i0_i54 (.D(d9_71__N_1674[54]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d9_i0_i55 (.D(d9_71__N_1674[55]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d9_i0_i56 (.D(d9_71__N_1674[56]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d9_i0_i57 (.D(d9_71__N_1674[57]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d9_i0_i58 (.D(d9_71__N_1674[58]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d9_i0_i59 (.D(d9_71__N_1674[59]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d9_i0_i60 (.D(d9_71__N_1674[60]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d9_i0_i61 (.D(d9_71__N_1674[61]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d9_i0_i62 (.D(d9_71__N_1674[62]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d9_i0_i63 (.D(d9_71__N_1674[63]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d9_i0_i64 (.D(d9_71__N_1674[64]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d9_i0_i65 (.D(d9_71__N_1674[65]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d9_i0_i66 (.D(d9_71__N_1674[66]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d9_i0_i67 (.D(d9_71__N_1674[67]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d9_i0_i68 (.D(d9_71__N_1674[68]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d9_i0_i69 (.D(d9_71__N_1674[69]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d9_i0_i70 (.D(d9_71__N_1674[70]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d9_i0_i71 (.D(d9_71__N_1674[71]), .SP(osc_clk_enable_1333), 
            .CK(osc_clk), .Q(d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i1 (.D(d9[1]), .SP(osc_clk_enable_1333), .CK(osc_clk), 
            .Q(d_d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i2 (.D(d9[2]), .SP(osc_clk_enable_1333), .CK(osc_clk), 
            .Q(d_d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i3 (.D(d9[3]), .SP(osc_clk_enable_1333), .CK(osc_clk), 
            .Q(d_d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i4 (.D(d9[4]), .SP(osc_clk_enable_1333), .CK(osc_clk), 
            .Q(d_d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i5 (.D(d9[5]), .SP(osc_clk_enable_1333), .CK(osc_clk), 
            .Q(d_d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i6 (.D(d9[6]), .SP(osc_clk_enable_1333), .CK(osc_clk), 
            .Q(d_d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i7 (.D(d9[7]), .SP(osc_clk_enable_1333), .CK(osc_clk), 
            .Q(d_d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i8 (.D(d9[8]), .SP(osc_clk_enable_1333), .CK(osc_clk), 
            .Q(d_d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i9 (.D(d9[9]), .SP(osc_clk_enable_1333), .CK(osc_clk), 
            .Q(d_d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i10 (.D(d9[10]), .SP(osc_clk_enable_1333), .CK(osc_clk), 
            .Q(d_d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i11 (.D(d9[11]), .SP(osc_clk_enable_1333), .CK(osc_clk), 
            .Q(d_d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i12 (.D(d9[12]), .SP(osc_clk_enable_1333), .CK(osc_clk), 
            .Q(d_d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i13 (.D(d9[13]), .SP(osc_clk_enable_1333), .CK(osc_clk), 
            .Q(d_d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i14 (.D(d9[14]), .SP(osc_clk_enable_1333), .CK(osc_clk), 
            .Q(d_d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i15 (.D(d9[15]), .SP(osc_clk_enable_1333), .CK(osc_clk), 
            .Q(d_d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i16 (.D(d9[16]), .SP(osc_clk_enable_1333), .CK(osc_clk), 
            .Q(d_d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i17 (.D(d9[17]), .SP(osc_clk_enable_1333), .CK(osc_clk), 
            .Q(d_d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i18 (.D(d9[18]), .SP(osc_clk_enable_1333), .CK(osc_clk), 
            .Q(d_d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i19 (.D(d9[19]), .SP(osc_clk_enable_1333), .CK(osc_clk), 
            .Q(d_d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i20 (.D(d9[20]), .SP(osc_clk_enable_1333), .CK(osc_clk), 
            .Q(d_d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i21 (.D(d9[21]), .SP(osc_clk_enable_1333), .CK(osc_clk), 
            .Q(d_d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i22 (.D(d9[22]), .SP(osc_clk_enable_1333), .CK(osc_clk), 
            .Q(d_d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i23 (.D(d9[23]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i24 (.D(d9[24]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i25 (.D(d9[25]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i26 (.D(d9[26]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i27 (.D(d9[27]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i28 (.D(d9[28]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i29 (.D(d9[29]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i30 (.D(d9[30]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i31 (.D(d9[31]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i32 (.D(d9[32]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i33 (.D(d9[33]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i34 (.D(d9[34]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i35 (.D(d9[35]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i36 (.D(d9[36]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i37 (.D(d9[37]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i38 (.D(d9[38]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i39 (.D(d9[39]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i40 (.D(d9[40]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i41 (.D(d9[41]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i42 (.D(d9[42]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i43 (.D(d9[43]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i44 (.D(d9[44]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i45 (.D(d9[45]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i46 (.D(d9[46]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i47 (.D(d9[47]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i48 (.D(d9[48]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i49 (.D(d9[49]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i50 (.D(d9[50]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i51 (.D(d9[51]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i52 (.D(d9[52]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i53 (.D(d9[53]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i54 (.D(d9[54]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i55 (.D(d9[55]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i56 (.D(d9[56]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i57 (.D(d9[57]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i58 (.D(d9[58]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i59 (.D(d9[59]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i60 (.D(d9[60]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i61 (.D(d9[61]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i62 (.D(d9[62]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i63 (.D(d9[63]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i64 (.D(d9[64]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i65 (.D(d9[65]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i66 (.D(d9[66]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i67 (.D(d9[67]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i68 (.D(d9[68]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i69 (.D(d9[69]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i70 (.D(d9[70]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i71 (.D(d9[71]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d_d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d10__i2 (.D(d10_71__N_1746[57]), .SP(osc_clk_enable_1383), .CK(osc_clk), 
            .Q(d10[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i2.GSR = "ENABLED";
    FD1P3AX d10__i3 (.D(d10_71__N_1746[58]), .SP(v_comb), .CK(osc_clk), 
            .Q(d10[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i3.GSR = "ENABLED";
    FD1P3AX d10__i4 (.D(d10_71__N_1746[59]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[59] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i4.GSR = "ENABLED";
    FD1P3AX d10__i5 (.D(d10_71__N_1746[60]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[60] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i5.GSR = "ENABLED";
    FD1P3AX d10__i6 (.D(d10_71__N_1746[61]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[61] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i6.GSR = "ENABLED";
    FD1P3AX d10__i7 (.D(d10_71__N_1746[62]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[62] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i7.GSR = "ENABLED";
    FD1P3AX d10__i8 (.D(d10_71__N_1746[63]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[63] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i8.GSR = "ENABLED";
    FD1P3AX d10__i9 (.D(d10_71__N_1746[64]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[64] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i9.GSR = "ENABLED";
    FD1P3AX d10__i10 (.D(d10_71__N_1746[65]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[65] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i10.GSR = "ENABLED";
    FD1P3AX d10__i11 (.D(d10_71__N_1746[66]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[66] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i11.GSR = "ENABLED";
    FD1P3AX d10__i12 (.D(d10_71__N_1746[67]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[67] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i12.GSR = "ENABLED";
    FD1P3AX d10__i13 (.D(d10_71__N_1746[68]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[68] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i13.GSR = "ENABLED";
    FD1P3AX d10__i14 (.D(d10_71__N_1746[69]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[69] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i14.GSR = "ENABLED";
    FD1P3AX d10__i15 (.D(d10_71__N_1746[70]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[70] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i15.GSR = "ENABLED";
    FD1P3AX d10__i16 (.D(d10_71__N_1746[71]), .SP(v_comb), .CK(osc_clk), 
            .Q(\d10[71] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d10__i16.GSR = "ENABLED";
    FD1P3AX d_out_i0_i1 (.D(d_out_11__N_1818[1]), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i1.GSR = "ENABLED";
    FD1P3AX d_out_i0_i2 (.D(\d_out_11__N_1818[2] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i2.GSR = "ENABLED";
    FD1P3AX d_out_i0_i3 (.D(\d_out_11__N_1818[3] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i3.GSR = "ENABLED";
    FD1P3AX d_out_i0_i4 (.D(\d_out_11__N_1818[4] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i4.GSR = "ENABLED";
    FD1P3AX d_out_i0_i5 (.D(\d_out_11__N_1818[5] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i5.GSR = "ENABLED";
    FD1P3AX d_out_i0_i6 (.D(\d_out_11__N_1818[6] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i6.GSR = "ENABLED";
    FD1P3AX d_out_i0_i7 (.D(\d_out_11__N_1818[7] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i7.GSR = "ENABLED";
    FD1P3AX d_out_i0_i8 (.D(\d_out_11__N_1818[8] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i8.GSR = "ENABLED";
    FD1P3AX d_out_i0_i9 (.D(\d_out_11__N_1818[9] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i9.GSR = "ENABLED";
    FD1P3AX d_out_i0_i10 (.D(\d_out_11__N_1818[10] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i10.GSR = "ENABLED";
    FD1P3AX d_out_i0_i11 (.D(\d_out_11__N_1818[11] ), .SP(v_comb), .CK(osc_clk), 
            .Q(CIC1_outCos[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(93[10] 121[8])
    defparam d_out_i0_i11.GSR = "ENABLED";
    FD1S3AX d1_i1 (.D(d1_71__N_417[1]), .CK(osc_clk), .Q(d1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i1.GSR = "ENABLED";
    FD1S3AX d1_i2 (.D(d1_71__N_417[2]), .CK(osc_clk), .Q(d1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i2.GSR = "ENABLED";
    FD1S3AX d1_i3 (.D(d1_71__N_417[3]), .CK(osc_clk), .Q(d1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i3.GSR = "ENABLED";
    FD1S3AX d1_i4 (.D(d1_71__N_417[4]), .CK(osc_clk), .Q(d1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i4.GSR = "ENABLED";
    FD1S3AX d1_i5 (.D(d1_71__N_417[5]), .CK(osc_clk), .Q(d1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i5.GSR = "ENABLED";
    FD1S3AX d1_i6 (.D(d1_71__N_417[6]), .CK(osc_clk), .Q(d1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i6.GSR = "ENABLED";
    FD1S3AX d1_i7 (.D(d1_71__N_417[7]), .CK(osc_clk), .Q(d1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i7.GSR = "ENABLED";
    FD1S3AX d1_i8 (.D(d1_71__N_417[8]), .CK(osc_clk), .Q(d1[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i8.GSR = "ENABLED";
    FD1S3AX d1_i9 (.D(d1_71__N_417[9]), .CK(osc_clk), .Q(d1[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i9.GSR = "ENABLED";
    FD1S3AX d1_i10 (.D(d1_71__N_417[10]), .CK(osc_clk), .Q(d1[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i10.GSR = "ENABLED";
    FD1S3AX d1_i11 (.D(d1_71__N_417[11]), .CK(osc_clk), .Q(d1[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i11.GSR = "ENABLED";
    FD1S3AX d1_i12 (.D(d1_71__N_417[12]), .CK(osc_clk), .Q(d1[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i12.GSR = "ENABLED";
    FD1S3AX d1_i13 (.D(d1_71__N_417[13]), .CK(osc_clk), .Q(d1[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i13.GSR = "ENABLED";
    FD1S3AX d1_i14 (.D(d1_71__N_417[14]), .CK(osc_clk), .Q(d1[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i14.GSR = "ENABLED";
    FD1S3AX d1_i15 (.D(d1_71__N_417[15]), .CK(osc_clk), .Q(d1[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i15.GSR = "ENABLED";
    FD1S3AX d1_i16 (.D(d1_71__N_417[16]), .CK(osc_clk), .Q(d1[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i16.GSR = "ENABLED";
    FD1S3AX d1_i17 (.D(d1_71__N_417[17]), .CK(osc_clk), .Q(d1[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i17.GSR = "ENABLED";
    FD1S3AX d1_i18 (.D(d1_71__N_417[18]), .CK(osc_clk), .Q(d1[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i18.GSR = "ENABLED";
    FD1S3AX d1_i19 (.D(d1_71__N_417[19]), .CK(osc_clk), .Q(d1[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i19.GSR = "ENABLED";
    FD1S3AX d1_i20 (.D(d1_71__N_417[20]), .CK(osc_clk), .Q(d1[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i20.GSR = "ENABLED";
    FD1S3AX d1_i21 (.D(d1_71__N_417[21]), .CK(osc_clk), .Q(d1[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i21.GSR = "ENABLED";
    FD1S3AX d1_i22 (.D(d1_71__N_417[22]), .CK(osc_clk), .Q(d1[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i22.GSR = "ENABLED";
    FD1S3AX d1_i23 (.D(d1_71__N_417[23]), .CK(osc_clk), .Q(d1[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i23.GSR = "ENABLED";
    FD1S3AX d1_i24 (.D(d1_71__N_417[24]), .CK(osc_clk), .Q(d1[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i24.GSR = "ENABLED";
    FD1S3AX d1_i25 (.D(d1_71__N_417[25]), .CK(osc_clk), .Q(d1[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i25.GSR = "ENABLED";
    FD1S3AX d1_i26 (.D(d1_71__N_417[26]), .CK(osc_clk), .Q(d1[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i26.GSR = "ENABLED";
    FD1S3AX d1_i27 (.D(d1_71__N_417[27]), .CK(osc_clk), .Q(d1[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i27.GSR = "ENABLED";
    FD1S3AX d1_i28 (.D(d1_71__N_417[28]), .CK(osc_clk), .Q(d1[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i28.GSR = "ENABLED";
    FD1S3AX d1_i29 (.D(d1_71__N_417[29]), .CK(osc_clk), .Q(d1[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i29.GSR = "ENABLED";
    FD1S3AX d1_i30 (.D(d1_71__N_417[30]), .CK(osc_clk), .Q(d1[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i30.GSR = "ENABLED";
    FD1S3AX d1_i31 (.D(d1_71__N_417[31]), .CK(osc_clk), .Q(d1[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i31.GSR = "ENABLED";
    FD1S3AX d1_i32 (.D(d1_71__N_417[32]), .CK(osc_clk), .Q(d1[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i32.GSR = "ENABLED";
    FD1S3AX d1_i33 (.D(d1_71__N_417[33]), .CK(osc_clk), .Q(d1[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i33.GSR = "ENABLED";
    FD1S3AX d1_i34 (.D(d1_71__N_417[34]), .CK(osc_clk), .Q(d1[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i34.GSR = "ENABLED";
    FD1S3AX d1_i35 (.D(d1_71__N_417[35]), .CK(osc_clk), .Q(d1[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i35.GSR = "ENABLED";
    FD1S3AX d1_i36 (.D(d1_71__N_417[36]), .CK(osc_clk), .Q(d1[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i36.GSR = "ENABLED";
    FD1S3AX d1_i37 (.D(d1_71__N_417[37]), .CK(osc_clk), .Q(d1[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i37.GSR = "ENABLED";
    FD1S3AX d1_i38 (.D(d1_71__N_417[38]), .CK(osc_clk), .Q(d1[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i38.GSR = "ENABLED";
    FD1S3AX d1_i39 (.D(d1_71__N_417[39]), .CK(osc_clk), .Q(d1[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i39.GSR = "ENABLED";
    FD1S3AX d1_i40 (.D(d1_71__N_417[40]), .CK(osc_clk), .Q(d1[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i40.GSR = "ENABLED";
    FD1S3AX d1_i41 (.D(d1_71__N_417[41]), .CK(osc_clk), .Q(d1[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i41.GSR = "ENABLED";
    FD1S3AX d1_i42 (.D(d1_71__N_417[42]), .CK(osc_clk), .Q(d1[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i42.GSR = "ENABLED";
    FD1S3AX d1_i43 (.D(d1_71__N_417[43]), .CK(osc_clk), .Q(d1[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i43.GSR = "ENABLED";
    FD1S3AX d1_i44 (.D(d1_71__N_417[44]), .CK(osc_clk), .Q(d1[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i44.GSR = "ENABLED";
    FD1S3AX d1_i45 (.D(d1_71__N_417[45]), .CK(osc_clk), .Q(d1[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i45.GSR = "ENABLED";
    FD1S3AX d1_i46 (.D(d1_71__N_417[46]), .CK(osc_clk), .Q(d1[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i46.GSR = "ENABLED";
    FD1S3AX d1_i47 (.D(d1_71__N_417[47]), .CK(osc_clk), .Q(d1[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i47.GSR = "ENABLED";
    FD1S3AX d1_i48 (.D(d1_71__N_417[48]), .CK(osc_clk), .Q(d1[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i48.GSR = "ENABLED";
    FD1S3AX d1_i49 (.D(d1_71__N_417[49]), .CK(osc_clk), .Q(d1[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i49.GSR = "ENABLED";
    FD1S3AX d1_i50 (.D(d1_71__N_417[50]), .CK(osc_clk), .Q(d1[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i50.GSR = "ENABLED";
    FD1S3AX d1_i51 (.D(d1_71__N_417[51]), .CK(osc_clk), .Q(d1[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i51.GSR = "ENABLED";
    FD1S3AX d1_i52 (.D(d1_71__N_417[52]), .CK(osc_clk), .Q(d1[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i52.GSR = "ENABLED";
    FD1S3AX d1_i53 (.D(d1_71__N_417[53]), .CK(osc_clk), .Q(d1[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i53.GSR = "ENABLED";
    FD1S3AX d1_i54 (.D(d1_71__N_417[54]), .CK(osc_clk), .Q(d1[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i54.GSR = "ENABLED";
    FD1S3AX d1_i55 (.D(d1_71__N_417[55]), .CK(osc_clk), .Q(d1[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i55.GSR = "ENABLED";
    FD1S3AX d1_i56 (.D(d1_71__N_417[56]), .CK(osc_clk), .Q(d1[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i56.GSR = "ENABLED";
    FD1S3AX d1_i57 (.D(d1_71__N_417[57]), .CK(osc_clk), .Q(d1[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i57.GSR = "ENABLED";
    FD1S3AX d1_i58 (.D(d1_71__N_417[58]), .CK(osc_clk), .Q(d1[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i58.GSR = "ENABLED";
    FD1S3AX d1_i59 (.D(d1_71__N_417[59]), .CK(osc_clk), .Q(d1[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i59.GSR = "ENABLED";
    FD1S3AX d1_i60 (.D(d1_71__N_417[60]), .CK(osc_clk), .Q(d1[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i60.GSR = "ENABLED";
    FD1S3AX d1_i61 (.D(d1_71__N_417[61]), .CK(osc_clk), .Q(d1[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i61.GSR = "ENABLED";
    FD1S3AX d1_i62 (.D(d1_71__N_417[62]), .CK(osc_clk), .Q(d1[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i62.GSR = "ENABLED";
    FD1S3AX d1_i63 (.D(d1_71__N_417[63]), .CK(osc_clk), .Q(d1[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i63.GSR = "ENABLED";
    FD1S3AX d1_i64 (.D(d1_71__N_417[64]), .CK(osc_clk), .Q(d1[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i64.GSR = "ENABLED";
    FD1S3AX d1_i65 (.D(d1_71__N_417[65]), .CK(osc_clk), .Q(d1[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i65.GSR = "ENABLED";
    FD1S3AX d1_i66 (.D(d1_71__N_417[66]), .CK(osc_clk), .Q(d1[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i66.GSR = "ENABLED";
    FD1S3AX d1_i67 (.D(d1_71__N_417[67]), .CK(osc_clk), .Q(d1[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i67.GSR = "ENABLED";
    FD1S3AX d1_i68 (.D(d1_71__N_417[68]), .CK(osc_clk), .Q(d1[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i68.GSR = "ENABLED";
    FD1S3AX d1_i69 (.D(d1_71__N_417[69]), .CK(osc_clk), .Q(d1[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i69.GSR = "ENABLED";
    FD1S3AX d1_i70 (.D(d1_71__N_417[70]), .CK(osc_clk), .Q(d1[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i70.GSR = "ENABLED";
    FD1S3AX d1_i71 (.D(d1_71__N_417[71]), .CK(osc_clk), .Q(d1[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam d1_i71.GSR = "ENABLED";
    LUT4 i5779_2_lut (.A(count[10]), .B(count[5]), .Z(n13228)) /* synthesis lut_function=(A (B)) */ ;
    defparam i5779_2_lut.init = 16'h8888;
    CCU2D add_1054_13 (.A0(d_d_tmp[46]), .B0(n6166), .C0(n6167[10]), .D0(d_tmp[46]), 
          .A1(d_d_tmp[47]), .B1(n6166), .C1(n6167[11]), .D1(d_tmp[47]), 
          .CIN(n11417), .COUT(n11418), .S0(d6_71__N_1458[46]), .S1(d6_71__N_1458[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1054_13.INIT0 = 16'hb874;
    defparam add_1054_13.INIT1 = 16'hb874;
    defparam add_1054_13.INJECT1_0 = "NO";
    defparam add_1054_13.INJECT1_1 = "NO";
    CCU2D add_1054_11 (.A0(d_d_tmp[44]), .B0(n6166), .C0(n6167[8]), .D0(d_tmp[44]), 
          .A1(d_d_tmp[45]), .B1(n6166), .C1(n6167[9]), .D1(d_tmp[45]), 
          .CIN(n11416), .COUT(n11417), .S0(d6_71__N_1458[44]), .S1(d6_71__N_1458[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1054_11.INIT0 = 16'hb874;
    defparam add_1054_11.INIT1 = 16'hb874;
    defparam add_1054_11.INJECT1_0 = "NO";
    defparam add_1054_11.INJECT1_1 = "NO";
    CCU2D add_1054_9 (.A0(d_d_tmp[42]), .B0(n6166), .C0(n6167[6]), .D0(d_tmp[42]), 
          .A1(d_d_tmp[43]), .B1(n6166), .C1(n6167[7]), .D1(d_tmp[43]), 
          .CIN(n11415), .COUT(n11416), .S0(d6_71__N_1458[42]), .S1(d6_71__N_1458[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1054_9.INIT0 = 16'hb874;
    defparam add_1054_9.INIT1 = 16'hb874;
    defparam add_1054_9.INJECT1_0 = "NO";
    defparam add_1054_9.INJECT1_1 = "NO";
    CCU2D add_1054_7 (.A0(d_d_tmp[40]), .B0(n6166), .C0(n6167[4]), .D0(d_tmp[40]), 
          .A1(d_d_tmp[41]), .B1(n6166), .C1(n6167[5]), .D1(d_tmp[41]), 
          .CIN(n11414), .COUT(n11415), .S0(d6_71__N_1458[40]), .S1(d6_71__N_1458[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1054_7.INIT0 = 16'hb874;
    defparam add_1054_7.INIT1 = 16'hb874;
    defparam add_1054_7.INJECT1_0 = "NO";
    defparam add_1054_7.INJECT1_1 = "NO";
    CCU2D add_1054_5 (.A0(d_d_tmp[38]), .B0(n6166), .C0(n6167[2]), .D0(d_tmp[38]), 
          .A1(d_d_tmp[39]), .B1(n6166), .C1(n6167[3]), .D1(d_tmp[39]), 
          .CIN(n11413), .COUT(n11414), .S0(d6_71__N_1458[38]), .S1(d6_71__N_1458[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1054_5.INIT0 = 16'hb874;
    defparam add_1054_5.INIT1 = 16'hb874;
    defparam add_1054_5.INJECT1_0 = "NO";
    defparam add_1054_5.INJECT1_1 = "NO";
    CCU2D add_1054_3 (.A0(d_d_tmp[36]), .B0(n6166), .C0(n6167[0]), .D0(d_tmp[36]), 
          .A1(d_d_tmp[37]), .B1(n6166), .C1(n6167[1]), .D1(d_tmp[37]), 
          .CIN(n11412), .COUT(n11413), .S0(d6_71__N_1458[36]), .S1(d6_71__N_1458[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1054_3.INIT0 = 16'hb874;
    defparam add_1054_3.INIT1 = 16'hb874;
    defparam add_1054_3.INJECT1_0 = "NO";
    defparam add_1054_3.INJECT1_1 = "NO";
    CCU2D add_1054_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n6166), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11412));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1054_1.INIT0 = 16'hF000;
    defparam add_1054_1.INIT1 = 16'h0555;
    defparam add_1054_1.INJECT1_0 = "NO";
    defparam add_1054_1.INJECT1_1 = "NO";
    LUT4 i4_4_lut (.A(n7), .B(count[15]), .C(count[11]), .D(count[14]), 
         .Z(n12867)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i4_4_lut.init = 16'hffef;
    CCU2D add_1014_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n4950), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11873));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1014_1.INIT0 = 16'hF000;
    defparam add_1014_1.INIT1 = 16'h0555;
    defparam add_1014_1.INJECT1_0 = "NO";
    defparam add_1014_1.INJECT1_1 = "NO";
    LUT4 shift_right_31_i61_3_lut (.A(\d10[60] ), .B(\d10[61] ), .C(\CICGain[0] ), 
         .Z(n61)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i61_3_lut.init = 16'hcaca;
    CCU2D add_1068_37 (.A0(d8[71]), .B0(d_d8[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11332), 
          .S0(n6623[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1068_37.INIT0 = 16'h5999;
    defparam add_1068_37.INIT1 = 16'h0000;
    defparam add_1068_37.INJECT1_0 = "NO";
    defparam add_1068_37.INJECT1_1 = "NO";
    CCU2D add_1068_35 (.A0(d8[69]), .B0(d_d8[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[70]), .B1(d_d8[70]), .C1(GND_net), .D1(GND_net), .CIN(n11331), 
          .COUT(n11332), .S0(n6623[33]), .S1(n6623[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1068_35.INIT0 = 16'h5999;
    defparam add_1068_35.INIT1 = 16'h5999;
    defparam add_1068_35.INJECT1_0 = "NO";
    defparam add_1068_35.INJECT1_1 = "NO";
    CCU2D add_1068_33 (.A0(d8[67]), .B0(d_d8[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[68]), .B1(d_d8[68]), .C1(GND_net), .D1(GND_net), .CIN(n11330), 
          .COUT(n11331), .S0(n6623[31]), .S1(n6623[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1068_33.INIT0 = 16'h5999;
    defparam add_1068_33.INIT1 = 16'h5999;
    defparam add_1068_33.INJECT1_0 = "NO";
    defparam add_1068_33.INJECT1_1 = "NO";
    CCU2D add_1068_31 (.A0(d8[65]), .B0(d_d8[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[66]), .B1(d_d8[66]), .C1(GND_net), .D1(GND_net), .CIN(n11329), 
          .COUT(n11330), .S0(n6623[29]), .S1(n6623[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1068_31.INIT0 = 16'h5999;
    defparam add_1068_31.INIT1 = 16'h5999;
    defparam add_1068_31.INJECT1_0 = "NO";
    defparam add_1068_31.INJECT1_1 = "NO";
    CCU2D add_1068_29 (.A0(d8[63]), .B0(d_d8[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[64]), .B1(d_d8[64]), .C1(GND_net), .D1(GND_net), .CIN(n11328), 
          .COUT(n11329), .S0(n6623[27]), .S1(n6623[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1068_29.INIT0 = 16'h5999;
    defparam add_1068_29.INIT1 = 16'h5999;
    defparam add_1068_29.INJECT1_0 = "NO";
    defparam add_1068_29.INJECT1_1 = "NO";
    CCU2D add_1068_27 (.A0(d8[61]), .B0(d_d8[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[62]), .B1(d_d8[62]), .C1(GND_net), .D1(GND_net), .CIN(n11327), 
          .COUT(n11328), .S0(n6623[25]), .S1(n6623[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1068_27.INIT0 = 16'h5999;
    defparam add_1068_27.INIT1 = 16'h5999;
    defparam add_1068_27.INJECT1_0 = "NO";
    defparam add_1068_27.INJECT1_1 = "NO";
    CCU2D add_1068_25 (.A0(d8[59]), .B0(d_d8[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[60]), .B1(d_d8[60]), .C1(GND_net), .D1(GND_net), .CIN(n11326), 
          .COUT(n11327), .S0(n6623[23]), .S1(n6623[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1068_25.INIT0 = 16'h5999;
    defparam add_1068_25.INIT1 = 16'h5999;
    defparam add_1068_25.INJECT1_0 = "NO";
    defparam add_1068_25.INJECT1_1 = "NO";
    CCU2D add_1068_23 (.A0(d8[57]), .B0(d_d8[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[58]), .B1(d_d8[58]), .C1(GND_net), .D1(GND_net), .CIN(n11325), 
          .COUT(n11326), .S0(n6623[21]), .S1(n6623[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1068_23.INIT0 = 16'h5999;
    defparam add_1068_23.INIT1 = 16'h5999;
    defparam add_1068_23.INJECT1_0 = "NO";
    defparam add_1068_23.INJECT1_1 = "NO";
    CCU2D add_1068_21 (.A0(d8[55]), .B0(d_d8[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[56]), .B1(d_d8[56]), .C1(GND_net), .D1(GND_net), .CIN(n11324), 
          .COUT(n11325), .S0(n6623[19]), .S1(n6623[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1068_21.INIT0 = 16'h5999;
    defparam add_1068_21.INIT1 = 16'h5999;
    defparam add_1068_21.INJECT1_0 = "NO";
    defparam add_1068_21.INJECT1_1 = "NO";
    CCU2D add_1068_19 (.A0(d8[53]), .B0(d_d8[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[54]), .B1(d_d8[54]), .C1(GND_net), .D1(GND_net), .CIN(n11323), 
          .COUT(n11324), .S0(n6623[17]), .S1(n6623[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1068_19.INIT0 = 16'h5999;
    defparam add_1068_19.INIT1 = 16'h5999;
    defparam add_1068_19.INJECT1_0 = "NO";
    defparam add_1068_19.INJECT1_1 = "NO";
    CCU2D add_1068_17 (.A0(d8[51]), .B0(d_d8[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[52]), .B1(d_d8[52]), .C1(GND_net), .D1(GND_net), .CIN(n11322), 
          .COUT(n11323), .S0(n6623[15]), .S1(n6623[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1068_17.INIT0 = 16'h5999;
    defparam add_1068_17.INIT1 = 16'h5999;
    defparam add_1068_17.INJECT1_0 = "NO";
    defparam add_1068_17.INJECT1_1 = "NO";
    CCU2D add_1068_15 (.A0(d8[49]), .B0(d_d8[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[50]), .B1(d_d8[50]), .C1(GND_net), .D1(GND_net), .CIN(n11321), 
          .COUT(n11322), .S0(n6623[13]), .S1(n6623[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1068_15.INIT0 = 16'h5999;
    defparam add_1068_15.INIT1 = 16'h5999;
    defparam add_1068_15.INJECT1_0 = "NO";
    defparam add_1068_15.INJECT1_1 = "NO";
    CCU2D add_1068_13 (.A0(d8[47]), .B0(d_d8[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[48]), .B1(d_d8[48]), .C1(GND_net), .D1(GND_net), .CIN(n11320), 
          .COUT(n11321), .S0(n6623[11]), .S1(n6623[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1068_13.INIT0 = 16'h5999;
    defparam add_1068_13.INIT1 = 16'h5999;
    defparam add_1068_13.INJECT1_0 = "NO";
    defparam add_1068_13.INJECT1_1 = "NO";
    CCU2D add_1068_11 (.A0(d8[45]), .B0(d_d8[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[46]), .B1(d_d8[46]), .C1(GND_net), .D1(GND_net), .CIN(n11319), 
          .COUT(n11320), .S0(n6623[9]), .S1(n6623[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1068_11.INIT0 = 16'h5999;
    defparam add_1068_11.INIT1 = 16'h5999;
    defparam add_1068_11.INJECT1_0 = "NO";
    defparam add_1068_11.INJECT1_1 = "NO";
    CCU2D add_1068_9 (.A0(d8[43]), .B0(d_d8[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[44]), .B1(d_d8[44]), .C1(GND_net), .D1(GND_net), .CIN(n11318), 
          .COUT(n11319), .S0(n6623[7]), .S1(n6623[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1068_9.INIT0 = 16'h5999;
    defparam add_1068_9.INIT1 = 16'h5999;
    defparam add_1068_9.INJECT1_0 = "NO";
    defparam add_1068_9.INJECT1_1 = "NO";
    CCU2D add_1068_7 (.A0(d8[41]), .B0(d_d8[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[42]), .B1(d_d8[42]), .C1(GND_net), .D1(GND_net), .CIN(n11317), 
          .COUT(n11318), .S0(n6623[5]), .S1(n6623[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1068_7.INIT0 = 16'h5999;
    defparam add_1068_7.INIT1 = 16'h5999;
    defparam add_1068_7.INJECT1_0 = "NO";
    defparam add_1068_7.INJECT1_1 = "NO";
    CCU2D add_1068_5 (.A0(d8[39]), .B0(d_d8[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[40]), .B1(d_d8[40]), .C1(GND_net), .D1(GND_net), .CIN(n11316), 
          .COUT(n11317), .S0(n6623[3]), .S1(n6623[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1068_5.INIT0 = 16'h5999;
    defparam add_1068_5.INIT1 = 16'h5999;
    defparam add_1068_5.INJECT1_0 = "NO";
    defparam add_1068_5.INJECT1_1 = "NO";
    CCU2D add_1068_3 (.A0(d8[37]), .B0(d_d8[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[38]), .B1(d_d8[38]), .C1(GND_net), .D1(GND_net), .CIN(n11315), 
          .COUT(n11316), .S0(n6623[1]), .S1(n6623[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1068_3.INIT0 = 16'h5999;
    defparam add_1068_3.INIT1 = 16'h5999;
    defparam add_1068_3.INJECT1_0 = "NO";
    defparam add_1068_3.INJECT1_1 = "NO";
    CCU2D add_1068_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d8[36]), .B1(d_d8[36]), .C1(GND_net), .D1(GND_net), .COUT(n11315), 
          .S1(n6623[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1068_1.INIT0 = 16'hF000;
    defparam add_1068_1.INIT1 = 16'h5999;
    defparam add_1068_1.INJECT1_0 = "NO";
    defparam add_1068_1.INJECT1_1 = "NO";
    CCU2D add_1069_37 (.A0(d_d8[70]), .B0(n6622), .C0(n6623[34]), .D0(d8[70]), 
          .A1(d_d8[71]), .B1(n6622), .C1(n6623[35]), .D1(d8[71]), .CIN(n11313), 
          .S0(d9_71__N_1674[70]), .S1(d9_71__N_1674[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1069_37.INIT0 = 16'hb874;
    defparam add_1069_37.INIT1 = 16'hb874;
    defparam add_1069_37.INJECT1_0 = "NO";
    defparam add_1069_37.INJECT1_1 = "NO";
    CCU2D add_1069_35 (.A0(d_d8[68]), .B0(n6622), .C0(n6623[32]), .D0(d8[68]), 
          .A1(d_d8[69]), .B1(n6622), .C1(n6623[33]), .D1(d8[69]), .CIN(n11312), 
          .COUT(n11313), .S0(d9_71__N_1674[68]), .S1(d9_71__N_1674[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1069_35.INIT0 = 16'hb874;
    defparam add_1069_35.INIT1 = 16'hb874;
    defparam add_1069_35.INJECT1_0 = "NO";
    defparam add_1069_35.INJECT1_1 = "NO";
    CCU2D add_1069_33 (.A0(d_d8[66]), .B0(n6622), .C0(n6623[30]), .D0(d8[66]), 
          .A1(d_d8[67]), .B1(n6622), .C1(n6623[31]), .D1(d8[67]), .CIN(n11311), 
          .COUT(n11312), .S0(d9_71__N_1674[66]), .S1(d9_71__N_1674[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1069_33.INIT0 = 16'hb874;
    defparam add_1069_33.INIT1 = 16'hb874;
    defparam add_1069_33.INJECT1_0 = "NO";
    defparam add_1069_33.INJECT1_1 = "NO";
    CCU2D add_1069_31 (.A0(d_d8[64]), .B0(n6622), .C0(n6623[28]), .D0(d8[64]), 
          .A1(d_d8[65]), .B1(n6622), .C1(n6623[29]), .D1(d8[65]), .CIN(n11310), 
          .COUT(n11311), .S0(d9_71__N_1674[64]), .S1(d9_71__N_1674[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1069_31.INIT0 = 16'hb874;
    defparam add_1069_31.INIT1 = 16'hb874;
    defparam add_1069_31.INJECT1_0 = "NO";
    defparam add_1069_31.INJECT1_1 = "NO";
    CCU2D add_1069_29 (.A0(d_d8[62]), .B0(n6622), .C0(n6623[26]), .D0(d8[62]), 
          .A1(d_d8[63]), .B1(n6622), .C1(n6623[27]), .D1(d8[63]), .CIN(n11309), 
          .COUT(n11310), .S0(d9_71__N_1674[62]), .S1(d9_71__N_1674[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1069_29.INIT0 = 16'hb874;
    defparam add_1069_29.INIT1 = 16'hb874;
    defparam add_1069_29.INJECT1_0 = "NO";
    defparam add_1069_29.INJECT1_1 = "NO";
    CCU2D add_1069_27 (.A0(d_d8[60]), .B0(n6622), .C0(n6623[24]), .D0(d8[60]), 
          .A1(d_d8[61]), .B1(n6622), .C1(n6623[25]), .D1(d8[61]), .CIN(n11308), 
          .COUT(n11309), .S0(d9_71__N_1674[60]), .S1(d9_71__N_1674[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1069_27.INIT0 = 16'hb874;
    defparam add_1069_27.INIT1 = 16'hb874;
    defparam add_1069_27.INJECT1_0 = "NO";
    defparam add_1069_27.INJECT1_1 = "NO";
    CCU2D add_1069_25 (.A0(d_d8[58]), .B0(n6622), .C0(n6623[22]), .D0(d8[58]), 
          .A1(d_d8[59]), .B1(n6622), .C1(n6623[23]), .D1(d8[59]), .CIN(n11307), 
          .COUT(n11308), .S0(d9_71__N_1674[58]), .S1(d9_71__N_1674[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1069_25.INIT0 = 16'hb874;
    defparam add_1069_25.INIT1 = 16'hb874;
    defparam add_1069_25.INJECT1_0 = "NO";
    defparam add_1069_25.INJECT1_1 = "NO";
    CCU2D add_1069_23 (.A0(d_d8[56]), .B0(n6622), .C0(n6623[20]), .D0(d8[56]), 
          .A1(d_d8[57]), .B1(n6622), .C1(n6623[21]), .D1(d8[57]), .CIN(n11306), 
          .COUT(n11307), .S0(d9_71__N_1674[56]), .S1(d9_71__N_1674[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1069_23.INIT0 = 16'hb874;
    defparam add_1069_23.INIT1 = 16'hb874;
    defparam add_1069_23.INJECT1_0 = "NO";
    defparam add_1069_23.INJECT1_1 = "NO";
    CCU2D add_1069_21 (.A0(d_d8[54]), .B0(n6622), .C0(n6623[18]), .D0(d8[54]), 
          .A1(d_d8[55]), .B1(n6622), .C1(n6623[19]), .D1(d8[55]), .CIN(n11305), 
          .COUT(n11306), .S0(d9_71__N_1674[54]), .S1(d9_71__N_1674[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1069_21.INIT0 = 16'hb874;
    defparam add_1069_21.INIT1 = 16'hb874;
    defparam add_1069_21.INJECT1_0 = "NO";
    defparam add_1069_21.INJECT1_1 = "NO";
    CCU2D add_1069_19 (.A0(d_d8[52]), .B0(n6622), .C0(n6623[16]), .D0(d8[52]), 
          .A1(d_d8[53]), .B1(n6622), .C1(n6623[17]), .D1(d8[53]), .CIN(n11304), 
          .COUT(n11305), .S0(d9_71__N_1674[52]), .S1(d9_71__N_1674[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1069_19.INIT0 = 16'hb874;
    defparam add_1069_19.INIT1 = 16'hb874;
    defparam add_1069_19.INJECT1_0 = "NO";
    defparam add_1069_19.INJECT1_1 = "NO";
    CCU2D add_1069_17 (.A0(d_d8[50]), .B0(n6622), .C0(n6623[14]), .D0(d8[50]), 
          .A1(d_d8[51]), .B1(n6622), .C1(n6623[15]), .D1(d8[51]), .CIN(n11303), 
          .COUT(n11304), .S0(d9_71__N_1674[50]), .S1(d9_71__N_1674[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1069_17.INIT0 = 16'hb874;
    defparam add_1069_17.INIT1 = 16'hb874;
    defparam add_1069_17.INJECT1_0 = "NO";
    defparam add_1069_17.INJECT1_1 = "NO";
    CCU2D add_1069_15 (.A0(d_d8[48]), .B0(n6622), .C0(n6623[12]), .D0(d8[48]), 
          .A1(d_d8[49]), .B1(n6622), .C1(n6623[13]), .D1(d8[49]), .CIN(n11302), 
          .COUT(n11303), .S0(d9_71__N_1674[48]), .S1(d9_71__N_1674[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1069_15.INIT0 = 16'hb874;
    defparam add_1069_15.INIT1 = 16'hb874;
    defparam add_1069_15.INJECT1_0 = "NO";
    defparam add_1069_15.INJECT1_1 = "NO";
    CCU2D add_1069_13 (.A0(d_d8[46]), .B0(n6622), .C0(n6623[10]), .D0(d8[46]), 
          .A1(d_d8[47]), .B1(n6622), .C1(n6623[11]), .D1(d8[47]), .CIN(n11301), 
          .COUT(n11302), .S0(d9_71__N_1674[46]), .S1(d9_71__N_1674[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1069_13.INIT0 = 16'hb874;
    defparam add_1069_13.INIT1 = 16'hb874;
    defparam add_1069_13.INJECT1_0 = "NO";
    defparam add_1069_13.INJECT1_1 = "NO";
    CCU2D add_1069_11 (.A0(d_d8[44]), .B0(n6622), .C0(n6623[8]), .D0(d8[44]), 
          .A1(d_d8[45]), .B1(n6622), .C1(n6623[9]), .D1(d8[45]), .CIN(n11300), 
          .COUT(n11301), .S0(d9_71__N_1674[44]), .S1(d9_71__N_1674[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1069_11.INIT0 = 16'hb874;
    defparam add_1069_11.INIT1 = 16'hb874;
    defparam add_1069_11.INJECT1_0 = "NO";
    defparam add_1069_11.INJECT1_1 = "NO";
    CCU2D add_1069_9 (.A0(d_d8[42]), .B0(n6622), .C0(n6623[6]), .D0(d8[42]), 
          .A1(d_d8[43]), .B1(n6622), .C1(n6623[7]), .D1(d8[43]), .CIN(n11299), 
          .COUT(n11300), .S0(d9_71__N_1674[42]), .S1(d9_71__N_1674[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1069_9.INIT0 = 16'hb874;
    defparam add_1069_9.INIT1 = 16'hb874;
    defparam add_1069_9.INJECT1_0 = "NO";
    defparam add_1069_9.INJECT1_1 = "NO";
    CCU2D add_1069_7 (.A0(d_d8[40]), .B0(n6622), .C0(n6623[4]), .D0(d8[40]), 
          .A1(d_d8[41]), .B1(n6622), .C1(n6623[5]), .D1(d8[41]), .CIN(n11298), 
          .COUT(n11299), .S0(d9_71__N_1674[40]), .S1(d9_71__N_1674[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1069_7.INIT0 = 16'hb874;
    defparam add_1069_7.INIT1 = 16'hb874;
    defparam add_1069_7.INJECT1_0 = "NO";
    defparam add_1069_7.INJECT1_1 = "NO";
    CCU2D add_1069_5 (.A0(d_d8[38]), .B0(n6622), .C0(n6623[2]), .D0(d8[38]), 
          .A1(d_d8[39]), .B1(n6622), .C1(n6623[3]), .D1(d8[39]), .CIN(n11297), 
          .COUT(n11298), .S0(d9_71__N_1674[38]), .S1(d9_71__N_1674[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1069_5.INIT0 = 16'hb874;
    defparam add_1069_5.INIT1 = 16'hb874;
    defparam add_1069_5.INJECT1_0 = "NO";
    defparam add_1069_5.INJECT1_1 = "NO";
    CCU2D add_1069_3 (.A0(d_d8[36]), .B0(n6622), .C0(n6623[0]), .D0(d8[36]), 
          .A1(d_d8[37]), .B1(n6622), .C1(n6623[1]), .D1(d8[37]), .CIN(n11296), 
          .COUT(n11297), .S0(d9_71__N_1674[36]), .S1(d9_71__N_1674[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1069_3.INIT0 = 16'hb874;
    defparam add_1069_3.INIT1 = 16'hb874;
    defparam add_1069_3.INJECT1_0 = "NO";
    defparam add_1069_3.INJECT1_1 = "NO";
    CCU2D add_1069_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n6622), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11296));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1069_1.INIT0 = 16'hF000;
    defparam add_1069_1.INIT1 = 16'h0555;
    defparam add_1069_1.INJECT1_0 = "NO";
    defparam add_1069_1.INJECT1_1 = "NO";
    CCU2D add_1073_37 (.A0(d9[71]), .B0(d_d9[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11292), 
          .S0(n6775[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1073_37.INIT0 = 16'h5999;
    defparam add_1073_37.INIT1 = 16'h0000;
    defparam add_1073_37.INJECT1_0 = "NO";
    defparam add_1073_37.INJECT1_1 = "NO";
    CCU2D add_1073_35 (.A0(d9[69]), .B0(d_d9[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[70]), .B1(d_d9[70]), .C1(GND_net), .D1(GND_net), .CIN(n11291), 
          .COUT(n11292), .S0(n6775[33]), .S1(n6775[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1073_35.INIT0 = 16'h5999;
    defparam add_1073_35.INIT1 = 16'h5999;
    defparam add_1073_35.INJECT1_0 = "NO";
    defparam add_1073_35.INJECT1_1 = "NO";
    CCU2D add_1073_33 (.A0(d9[67]), .B0(d_d9[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[68]), .B1(d_d9[68]), .C1(GND_net), .D1(GND_net), .CIN(n11290), 
          .COUT(n11291), .S0(n6775[31]), .S1(n6775[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1073_33.INIT0 = 16'h5999;
    defparam add_1073_33.INIT1 = 16'h5999;
    defparam add_1073_33.INJECT1_0 = "NO";
    defparam add_1073_33.INJECT1_1 = "NO";
    CCU2D add_1073_31 (.A0(d9[65]), .B0(d_d9[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[66]), .B1(d_d9[66]), .C1(GND_net), .D1(GND_net), .CIN(n11289), 
          .COUT(n11290), .S0(n6775[29]), .S1(n6775[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1073_31.INIT0 = 16'h5999;
    defparam add_1073_31.INIT1 = 16'h5999;
    defparam add_1073_31.INJECT1_0 = "NO";
    defparam add_1073_31.INJECT1_1 = "NO";
    CCU2D add_1073_29 (.A0(d9[63]), .B0(d_d9[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[64]), .B1(d_d9[64]), .C1(GND_net), .D1(GND_net), .CIN(n11288), 
          .COUT(n11289), .S0(n6775[27]), .S1(n6775[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1073_29.INIT0 = 16'h5999;
    defparam add_1073_29.INIT1 = 16'h5999;
    defparam add_1073_29.INJECT1_0 = "NO";
    defparam add_1073_29.INJECT1_1 = "NO";
    CCU2D add_1073_27 (.A0(d9[61]), .B0(d_d9[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[62]), .B1(d_d9[62]), .C1(GND_net), .D1(GND_net), .CIN(n11287), 
          .COUT(n11288), .S0(n6775[25]), .S1(n6775[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1073_27.INIT0 = 16'h5999;
    defparam add_1073_27.INIT1 = 16'h5999;
    defparam add_1073_27.INJECT1_0 = "NO";
    defparam add_1073_27.INJECT1_1 = "NO";
    CCU2D add_1073_25 (.A0(d9[59]), .B0(d_d9[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[60]), .B1(d_d9[60]), .C1(GND_net), .D1(GND_net), .CIN(n11286), 
          .COUT(n11287), .S0(n6775[23]), .S1(n6775[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1073_25.INIT0 = 16'h5999;
    defparam add_1073_25.INIT1 = 16'h5999;
    defparam add_1073_25.INJECT1_0 = "NO";
    defparam add_1073_25.INJECT1_1 = "NO";
    CCU2D add_1073_23 (.A0(d9[57]), .B0(d_d9[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[58]), .B1(d_d9[58]), .C1(GND_net), .D1(GND_net), .CIN(n11285), 
          .COUT(n11286), .S0(n6775[21]), .S1(n6775[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1073_23.INIT0 = 16'h5999;
    defparam add_1073_23.INIT1 = 16'h5999;
    defparam add_1073_23.INJECT1_0 = "NO";
    defparam add_1073_23.INJECT1_1 = "NO";
    CCU2D add_1073_21 (.A0(d9[55]), .B0(d_d9[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[56]), .B1(d_d9[56]), .C1(GND_net), .D1(GND_net), .CIN(n11284), 
          .COUT(n11285));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1073_21.INIT0 = 16'h5999;
    defparam add_1073_21.INIT1 = 16'h5999;
    defparam add_1073_21.INJECT1_0 = "NO";
    defparam add_1073_21.INJECT1_1 = "NO";
    CCU2D add_1073_19 (.A0(d9[53]), .B0(d_d9[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[54]), .B1(d_d9[54]), .C1(GND_net), .D1(GND_net), .CIN(n11283), 
          .COUT(n11284));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1073_19.INIT0 = 16'h5999;
    defparam add_1073_19.INIT1 = 16'h5999;
    defparam add_1073_19.INJECT1_0 = "NO";
    defparam add_1073_19.INJECT1_1 = "NO";
    CCU2D add_1073_17 (.A0(d9[51]), .B0(d_d9[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[52]), .B1(d_d9[52]), .C1(GND_net), .D1(GND_net), .CIN(n11282), 
          .COUT(n11283));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1073_17.INIT0 = 16'h5999;
    defparam add_1073_17.INIT1 = 16'h5999;
    defparam add_1073_17.INJECT1_0 = "NO";
    defparam add_1073_17.INJECT1_1 = "NO";
    CCU2D add_1073_15 (.A0(d9[49]), .B0(d_d9[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[50]), .B1(d_d9[50]), .C1(GND_net), .D1(GND_net), .CIN(n11281), 
          .COUT(n11282));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1073_15.INIT0 = 16'h5999;
    defparam add_1073_15.INIT1 = 16'h5999;
    defparam add_1073_15.INJECT1_0 = "NO";
    defparam add_1073_15.INJECT1_1 = "NO";
    CCU2D add_1073_13 (.A0(d9[47]), .B0(d_d9[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[48]), .B1(d_d9[48]), .C1(GND_net), .D1(GND_net), .CIN(n11280), 
          .COUT(n11281));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1073_13.INIT0 = 16'h5999;
    defparam add_1073_13.INIT1 = 16'h5999;
    defparam add_1073_13.INJECT1_0 = "NO";
    defparam add_1073_13.INJECT1_1 = "NO";
    CCU2D add_1073_11 (.A0(d9[45]), .B0(d_d9[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[46]), .B1(d_d9[46]), .C1(GND_net), .D1(GND_net), .CIN(n11279), 
          .COUT(n11280));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1073_11.INIT0 = 16'h5999;
    defparam add_1073_11.INIT1 = 16'h5999;
    defparam add_1073_11.INJECT1_0 = "NO";
    defparam add_1073_11.INJECT1_1 = "NO";
    CCU2D add_1073_9 (.A0(d9[43]), .B0(d_d9[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[44]), .B1(d_d9[44]), .C1(GND_net), .D1(GND_net), .CIN(n11278), 
          .COUT(n11279));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1073_9.INIT0 = 16'h5999;
    defparam add_1073_9.INIT1 = 16'h5999;
    defparam add_1073_9.INJECT1_0 = "NO";
    defparam add_1073_9.INJECT1_1 = "NO";
    CCU2D add_1073_7 (.A0(d9[41]), .B0(d_d9[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[42]), .B1(d_d9[42]), .C1(GND_net), .D1(GND_net), .CIN(n11277), 
          .COUT(n11278));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1073_7.INIT0 = 16'h5999;
    defparam add_1073_7.INIT1 = 16'h5999;
    defparam add_1073_7.INJECT1_0 = "NO";
    defparam add_1073_7.INJECT1_1 = "NO";
    CCU2D add_1073_5 (.A0(d9[39]), .B0(d_d9[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[40]), .B1(d_d9[40]), .C1(GND_net), .D1(GND_net), .CIN(n11276), 
          .COUT(n11277));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1073_5.INIT0 = 16'h5999;
    defparam add_1073_5.INIT1 = 16'h5999;
    defparam add_1073_5.INJECT1_0 = "NO";
    defparam add_1073_5.INJECT1_1 = "NO";
    CCU2D add_1073_3 (.A0(d9[37]), .B0(d_d9[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[38]), .B1(d_d9[38]), .C1(GND_net), .D1(GND_net), .CIN(n11275), 
          .COUT(n11276));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1073_3.INIT0 = 16'h5999;
    defparam add_1073_3.INIT1 = 16'h5999;
    defparam add_1073_3.INJECT1_0 = "NO";
    defparam add_1073_3.INJECT1_1 = "NO";
    CCU2D add_1073_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d9[36]), .B1(d_d9[36]), .C1(GND_net), .D1(GND_net), .COUT(n11275));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1073_1.INIT0 = 16'hF000;
    defparam add_1073_1.INIT1 = 16'h5999;
    defparam add_1073_1.INJECT1_0 = "NO";
    defparam add_1073_1.INJECT1_1 = "NO";
    CCU2D add_1074_37 (.A0(d9[71]), .B0(d_d9[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11274), 
          .S0(n6813[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1074_37.INIT0 = 16'h5999;
    defparam add_1074_37.INIT1 = 16'h0000;
    defparam add_1074_37.INJECT1_0 = "NO";
    defparam add_1074_37.INJECT1_1 = "NO";
    CCU2D add_1074_35 (.A0(d9[69]), .B0(d_d9[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[70]), .B1(d_d9[70]), .C1(GND_net), .D1(GND_net), .CIN(n11273), 
          .COUT(n11274), .S0(n6813[33]), .S1(n6813[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1074_35.INIT0 = 16'h5999;
    defparam add_1074_35.INIT1 = 16'h5999;
    defparam add_1074_35.INJECT1_0 = "NO";
    defparam add_1074_35.INJECT1_1 = "NO";
    CCU2D add_1074_33 (.A0(d9[67]), .B0(d_d9[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[68]), .B1(d_d9[68]), .C1(GND_net), .D1(GND_net), .CIN(n11272), 
          .COUT(n11273), .S0(n6813[31]), .S1(n6813[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1074_33.INIT0 = 16'h5999;
    defparam add_1074_33.INIT1 = 16'h5999;
    defparam add_1074_33.INJECT1_0 = "NO";
    defparam add_1074_33.INJECT1_1 = "NO";
    CCU2D add_1074_31 (.A0(d9[65]), .B0(d_d9[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[66]), .B1(d_d9[66]), .C1(GND_net), .D1(GND_net), .CIN(n11271), 
          .COUT(n11272), .S0(n6813[29]), .S1(n6813[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1074_31.INIT0 = 16'h5999;
    defparam add_1074_31.INIT1 = 16'h5999;
    defparam add_1074_31.INJECT1_0 = "NO";
    defparam add_1074_31.INJECT1_1 = "NO";
    CCU2D add_1074_29 (.A0(d9[63]), .B0(d_d9[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[64]), .B1(d_d9[64]), .C1(GND_net), .D1(GND_net), .CIN(n11270), 
          .COUT(n11271), .S0(n6813[27]), .S1(n6813[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1074_29.INIT0 = 16'h5999;
    defparam add_1074_29.INIT1 = 16'h5999;
    defparam add_1074_29.INJECT1_0 = "NO";
    defparam add_1074_29.INJECT1_1 = "NO";
    CCU2D add_1074_27 (.A0(d9[61]), .B0(d_d9[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[62]), .B1(d_d9[62]), .C1(GND_net), .D1(GND_net), .CIN(n11269), 
          .COUT(n11270), .S0(n6813[25]), .S1(n6813[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1074_27.INIT0 = 16'h5999;
    defparam add_1074_27.INIT1 = 16'h5999;
    defparam add_1074_27.INJECT1_0 = "NO";
    defparam add_1074_27.INJECT1_1 = "NO";
    CCU2D add_1074_25 (.A0(d9[59]), .B0(d_d9[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[60]), .B1(d_d9[60]), .C1(GND_net), .D1(GND_net), .CIN(n11268), 
          .COUT(n11269), .S0(n6813[23]), .S1(n6813[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1074_25.INIT0 = 16'h5999;
    defparam add_1074_25.INIT1 = 16'h5999;
    defparam add_1074_25.INJECT1_0 = "NO";
    defparam add_1074_25.INJECT1_1 = "NO";
    CCU2D add_1074_23 (.A0(d9[57]), .B0(d_d9[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[58]), .B1(d_d9[58]), .C1(GND_net), .D1(GND_net), .CIN(n11267), 
          .COUT(n11268), .S0(n6813[21]), .S1(n6813[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1074_23.INIT0 = 16'h5999;
    defparam add_1074_23.INIT1 = 16'h5999;
    defparam add_1074_23.INJECT1_0 = "NO";
    defparam add_1074_23.INJECT1_1 = "NO";
    CCU2D add_1074_21 (.A0(d9[55]), .B0(d_d9[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[56]), .B1(d_d9[56]), .C1(GND_net), .D1(GND_net), .CIN(n11266), 
          .COUT(n11267));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1074_21.INIT0 = 16'h5999;
    defparam add_1074_21.INIT1 = 16'h5999;
    defparam add_1074_21.INJECT1_0 = "NO";
    defparam add_1074_21.INJECT1_1 = "NO";
    CCU2D add_1074_19 (.A0(d9[53]), .B0(d_d9[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[54]), .B1(d_d9[54]), .C1(GND_net), .D1(GND_net), .CIN(n11265), 
          .COUT(n11266));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1074_19.INIT0 = 16'h5999;
    defparam add_1074_19.INIT1 = 16'h5999;
    defparam add_1074_19.INJECT1_0 = "NO";
    defparam add_1074_19.INJECT1_1 = "NO";
    CCU2D add_1074_17 (.A0(d9[51]), .B0(d_d9[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[52]), .B1(d_d9[52]), .C1(GND_net), .D1(GND_net), .CIN(n11264), 
          .COUT(n11265));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1074_17.INIT0 = 16'h5999;
    defparam add_1074_17.INIT1 = 16'h5999;
    defparam add_1074_17.INJECT1_0 = "NO";
    defparam add_1074_17.INJECT1_1 = "NO";
    CCU2D add_1074_15 (.A0(d9[49]), .B0(d_d9[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[50]), .B1(d_d9[50]), .C1(GND_net), .D1(GND_net), .CIN(n11263), 
          .COUT(n11264));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1074_15.INIT0 = 16'h5999;
    defparam add_1074_15.INIT1 = 16'h5999;
    defparam add_1074_15.INJECT1_0 = "NO";
    defparam add_1074_15.INJECT1_1 = "NO";
    CCU2D add_1074_13 (.A0(d9[47]), .B0(d_d9[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[48]), .B1(d_d9[48]), .C1(GND_net), .D1(GND_net), .CIN(n11262), 
          .COUT(n11263));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1074_13.INIT0 = 16'h5999;
    defparam add_1074_13.INIT1 = 16'h5999;
    defparam add_1074_13.INJECT1_0 = "NO";
    defparam add_1074_13.INJECT1_1 = "NO";
    CCU2D add_1074_11 (.A0(d9[45]), .B0(d_d9[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[46]), .B1(d_d9[46]), .C1(GND_net), .D1(GND_net), .CIN(n11261), 
          .COUT(n11262));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1074_11.INIT0 = 16'h5999;
    defparam add_1074_11.INIT1 = 16'h5999;
    defparam add_1074_11.INJECT1_0 = "NO";
    defparam add_1074_11.INJECT1_1 = "NO";
    CCU2D add_1074_9 (.A0(d9[43]), .B0(d_d9[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[44]), .B1(d_d9[44]), .C1(GND_net), .D1(GND_net), .CIN(n11260), 
          .COUT(n11261));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1074_9.INIT0 = 16'h5999;
    defparam add_1074_9.INIT1 = 16'h5999;
    defparam add_1074_9.INJECT1_0 = "NO";
    defparam add_1074_9.INJECT1_1 = "NO";
    CCU2D add_1074_7 (.A0(d9[41]), .B0(d_d9[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[42]), .B1(d_d9[42]), .C1(GND_net), .D1(GND_net), .CIN(n11259), 
          .COUT(n11260));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1074_7.INIT0 = 16'h5999;
    defparam add_1074_7.INIT1 = 16'h5999;
    defparam add_1074_7.INJECT1_0 = "NO";
    defparam add_1074_7.INJECT1_1 = "NO";
    CCU2D add_1074_5 (.A0(d9[39]), .B0(d_d9[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[40]), .B1(d_d9[40]), .C1(GND_net), .D1(GND_net), .CIN(n11258), 
          .COUT(n11259));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1074_5.INIT0 = 16'h5999;
    defparam add_1074_5.INIT1 = 16'h5999;
    defparam add_1074_5.INJECT1_0 = "NO";
    defparam add_1074_5.INJECT1_1 = "NO";
    CCU2D add_1074_3 (.A0(d9[37]), .B0(d_d9[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[38]), .B1(d_d9[38]), .C1(GND_net), .D1(GND_net), .CIN(n11257), 
          .COUT(n11258));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1074_3.INIT0 = 16'h5999;
    defparam add_1074_3.INIT1 = 16'h5999;
    defparam add_1074_3.INJECT1_0 = "NO";
    defparam add_1074_3.INJECT1_1 = "NO";
    CCU2D add_1074_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d9[36]), .B1(d_d9[36]), .C1(GND_net), .D1(GND_net), .COUT(n11257));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1074_1.INIT0 = 16'h0000;
    defparam add_1074_1.INIT1 = 16'h5999;
    defparam add_1074_1.INJECT1_0 = "NO";
    defparam add_1074_1.INJECT1_1 = "NO";
    CCU2D add_1013_18 (.A0(d1[52]), .B0(d2[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[53]), .B1(d2[53]), .C1(GND_net), .D1(GND_net), .CIN(n11900), 
          .COUT(n11901), .S0(n4951[16]), .S1(n4951[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1013_18.INIT0 = 16'h5666;
    defparam add_1013_18.INIT1 = 16'h5666;
    defparam add_1013_18.INJECT1_0 = "NO";
    defparam add_1013_18.INJECT1_1 = "NO";
    LUT4 i4803_2_lut (.A(MixerOutCos[11]), .B(d1[36]), .Z(n4799[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4803_2_lut.init = 16'h6666;
    LUT4 i2_2_lut (.A(count[13]), .B(count[12]), .Z(n7)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    CCU2D add_1043_37 (.A0(d7[71]), .B0(d_d7[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11666), 
          .S0(n5863[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1043_37.INIT0 = 16'h5999;
    defparam add_1043_37.INIT1 = 16'h0000;
    defparam add_1043_37.INJECT1_0 = "NO";
    defparam add_1043_37.INJECT1_1 = "NO";
    CCU2D add_1043_35 (.A0(d7[69]), .B0(d_d7[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[70]), .B1(d_d7[70]), .C1(GND_net), .D1(GND_net), .CIN(n11665), 
          .COUT(n11666), .S0(n5863[33]), .S1(n5863[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1043_35.INIT0 = 16'h5999;
    defparam add_1043_35.INIT1 = 16'h5999;
    defparam add_1043_35.INJECT1_0 = "NO";
    defparam add_1043_35.INJECT1_1 = "NO";
    LUT4 i5849_4_lut_rep_197 (.A(n13248), .B(n13), .C(n13250), .D(n13228), 
         .Z(n14125)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i5849_4_lut_rep_197.init = 16'h2000;
    CCU2D add_1043_33 (.A0(d7[67]), .B0(d_d7[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[68]), .B1(d_d7[68]), .C1(GND_net), .D1(GND_net), .CIN(n11664), 
          .COUT(n11665), .S0(n5863[31]), .S1(n5863[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1043_33.INIT0 = 16'h5999;
    defparam add_1043_33.INIT1 = 16'h5999;
    defparam add_1043_33.INJECT1_0 = "NO";
    defparam add_1043_33.INJECT1_1 = "NO";
    CCU2D add_1043_31 (.A0(d7[65]), .B0(d_d7[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[66]), .B1(d_d7[66]), .C1(GND_net), .D1(GND_net), .CIN(n11663), 
          .COUT(n11664), .S0(n5863[29]), .S1(n5863[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1043_31.INIT0 = 16'h5999;
    defparam add_1043_31.INIT1 = 16'h5999;
    defparam add_1043_31.INJECT1_0 = "NO";
    defparam add_1043_31.INJECT1_1 = "NO";
    CCU2D add_1043_29 (.A0(d7[63]), .B0(d_d7[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[64]), .B1(d_d7[64]), .C1(GND_net), .D1(GND_net), .CIN(n11662), 
          .COUT(n11663), .S0(n5863[27]), .S1(n5863[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1043_29.INIT0 = 16'h5999;
    defparam add_1043_29.INIT1 = 16'h5999;
    defparam add_1043_29.INJECT1_0 = "NO";
    defparam add_1043_29.INJECT1_1 = "NO";
    CCU2D add_1043_27 (.A0(d7[61]), .B0(d_d7[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[62]), .B1(d_d7[62]), .C1(GND_net), .D1(GND_net), .CIN(n11661), 
          .COUT(n11662), .S0(n5863[25]), .S1(n5863[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1043_27.INIT0 = 16'h5999;
    defparam add_1043_27.INIT1 = 16'h5999;
    defparam add_1043_27.INJECT1_0 = "NO";
    defparam add_1043_27.INJECT1_1 = "NO";
    CCU2D add_1043_25 (.A0(d7[59]), .B0(d_d7[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[60]), .B1(d_d7[60]), .C1(GND_net), .D1(GND_net), .CIN(n11660), 
          .COUT(n11661), .S0(n5863[23]), .S1(n5863[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1043_25.INIT0 = 16'h5999;
    defparam add_1043_25.INIT1 = 16'h5999;
    defparam add_1043_25.INJECT1_0 = "NO";
    defparam add_1043_25.INJECT1_1 = "NO";
    CCU2D add_1043_23 (.A0(d7[57]), .B0(d_d7[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[58]), .B1(d_d7[58]), .C1(GND_net), .D1(GND_net), .CIN(n11659), 
          .COUT(n11660), .S0(n5863[21]), .S1(n5863[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1043_23.INIT0 = 16'h5999;
    defparam add_1043_23.INIT1 = 16'h5999;
    defparam add_1043_23.INJECT1_0 = "NO";
    defparam add_1043_23.INJECT1_1 = "NO";
    CCU2D add_1043_21 (.A0(d7[55]), .B0(d_d7[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[56]), .B1(d_d7[56]), .C1(GND_net), .D1(GND_net), .CIN(n11658), 
          .COUT(n11659), .S0(n5863[19]), .S1(n5863[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1043_21.INIT0 = 16'h5999;
    defparam add_1043_21.INIT1 = 16'h5999;
    defparam add_1043_21.INJECT1_0 = "NO";
    defparam add_1043_21.INJECT1_1 = "NO";
    CCU2D add_1043_19 (.A0(d7[53]), .B0(d_d7[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[54]), .B1(d_d7[54]), .C1(GND_net), .D1(GND_net), .CIN(n11657), 
          .COUT(n11658), .S0(n5863[17]), .S1(n5863[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1043_19.INIT0 = 16'h5999;
    defparam add_1043_19.INIT1 = 16'h5999;
    defparam add_1043_19.INJECT1_0 = "NO";
    defparam add_1043_19.INJECT1_1 = "NO";
    CCU2D add_1043_17 (.A0(d7[51]), .B0(d_d7[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[52]), .B1(d_d7[52]), .C1(GND_net), .D1(GND_net), .CIN(n11656), 
          .COUT(n11657), .S0(n5863[15]), .S1(n5863[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1043_17.INIT0 = 16'h5999;
    defparam add_1043_17.INIT1 = 16'h5999;
    defparam add_1043_17.INJECT1_0 = "NO";
    defparam add_1043_17.INJECT1_1 = "NO";
    CCU2D add_1043_15 (.A0(d7[49]), .B0(d_d7[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[50]), .B1(d_d7[50]), .C1(GND_net), .D1(GND_net), .CIN(n11655), 
          .COUT(n11656), .S0(n5863[13]), .S1(n5863[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1043_15.INIT0 = 16'h5999;
    defparam add_1043_15.INIT1 = 16'h5999;
    defparam add_1043_15.INJECT1_0 = "NO";
    defparam add_1043_15.INJECT1_1 = "NO";
    CCU2D add_1043_13 (.A0(d7[47]), .B0(d_d7[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[48]), .B1(d_d7[48]), .C1(GND_net), .D1(GND_net), .CIN(n11654), 
          .COUT(n11655), .S0(n5863[11]), .S1(n5863[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1043_13.INIT0 = 16'h5999;
    defparam add_1043_13.INIT1 = 16'h5999;
    defparam add_1043_13.INJECT1_0 = "NO";
    defparam add_1043_13.INJECT1_1 = "NO";
    CCU2D add_1043_11 (.A0(d7[45]), .B0(d_d7[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[46]), .B1(d_d7[46]), .C1(GND_net), .D1(GND_net), .CIN(n11653), 
          .COUT(n11654), .S0(n5863[9]), .S1(n5863[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1043_11.INIT0 = 16'h5999;
    defparam add_1043_11.INIT1 = 16'h5999;
    defparam add_1043_11.INJECT1_0 = "NO";
    defparam add_1043_11.INJECT1_1 = "NO";
    CCU2D add_1043_9 (.A0(d7[43]), .B0(d_d7[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[44]), .B1(d_d7[44]), .C1(GND_net), .D1(GND_net), .CIN(n11652), 
          .COUT(n11653), .S0(n5863[7]), .S1(n5863[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1043_9.INIT0 = 16'h5999;
    defparam add_1043_9.INIT1 = 16'h5999;
    defparam add_1043_9.INJECT1_0 = "NO";
    defparam add_1043_9.INJECT1_1 = "NO";
    CCU2D add_1043_7 (.A0(d7[41]), .B0(d_d7[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[42]), .B1(d_d7[42]), .C1(GND_net), .D1(GND_net), .CIN(n11651), 
          .COUT(n11652), .S0(n5863[5]), .S1(n5863[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1043_7.INIT0 = 16'h5999;
    defparam add_1043_7.INIT1 = 16'h5999;
    defparam add_1043_7.INJECT1_0 = "NO";
    defparam add_1043_7.INJECT1_1 = "NO";
    CCU2D add_1043_5 (.A0(d7[39]), .B0(d_d7[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[40]), .B1(d_d7[40]), .C1(GND_net), .D1(GND_net), .CIN(n11650), 
          .COUT(n11651), .S0(n5863[3]), .S1(n5863[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1043_5.INIT0 = 16'h5999;
    defparam add_1043_5.INIT1 = 16'h5999;
    defparam add_1043_5.INJECT1_0 = "NO";
    defparam add_1043_5.INJECT1_1 = "NO";
    CCU2D add_1072_37 (.A0(d9[35]), .B0(d_d9[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11150), 
          .S1(n6774));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1072_37.INIT0 = 16'h5999;
    defparam add_1072_37.INIT1 = 16'h0000;
    defparam add_1072_37.INJECT1_0 = "NO";
    defparam add_1072_37.INJECT1_1 = "NO";
    CCU2D add_1072_35 (.A0(d9[33]), .B0(d_d9[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[34]), .B1(d_d9[34]), .C1(GND_net), .D1(GND_net), .CIN(n11149), 
          .COUT(n11150));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1072_35.INIT0 = 16'h5999;
    defparam add_1072_35.INIT1 = 16'h5999;
    defparam add_1072_35.INJECT1_0 = "NO";
    defparam add_1072_35.INJECT1_1 = "NO";
    CCU2D add_1072_33 (.A0(d9[31]), .B0(d_d9[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[32]), .B1(d_d9[32]), .C1(GND_net), .D1(GND_net), .CIN(n11148), 
          .COUT(n11149));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1072_33.INIT0 = 16'h5999;
    defparam add_1072_33.INIT1 = 16'h5999;
    defparam add_1072_33.INJECT1_0 = "NO";
    defparam add_1072_33.INJECT1_1 = "NO";
    CCU2D add_1072_31 (.A0(d9[29]), .B0(d_d9[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[30]), .B1(d_d9[30]), .C1(GND_net), .D1(GND_net), .CIN(n11147), 
          .COUT(n11148));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1072_31.INIT0 = 16'h5999;
    defparam add_1072_31.INIT1 = 16'h5999;
    defparam add_1072_31.INJECT1_0 = "NO";
    defparam add_1072_31.INJECT1_1 = "NO";
    CCU2D add_1072_29 (.A0(d9[27]), .B0(d_d9[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[28]), .B1(d_d9[28]), .C1(GND_net), .D1(GND_net), .CIN(n11146), 
          .COUT(n11147));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1072_29.INIT0 = 16'h5999;
    defparam add_1072_29.INIT1 = 16'h5999;
    defparam add_1072_29.INJECT1_0 = "NO";
    defparam add_1072_29.INJECT1_1 = "NO";
    CCU2D add_1072_27 (.A0(d9[25]), .B0(d_d9[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[26]), .B1(d_d9[26]), .C1(GND_net), .D1(GND_net), .CIN(n11145), 
          .COUT(n11146));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1072_27.INIT0 = 16'h5999;
    defparam add_1072_27.INIT1 = 16'h5999;
    defparam add_1072_27.INJECT1_0 = "NO";
    defparam add_1072_27.INJECT1_1 = "NO";
    CCU2D add_1072_25 (.A0(d9[23]), .B0(d_d9[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[24]), .B1(d_d9[24]), .C1(GND_net), .D1(GND_net), .CIN(n11144), 
          .COUT(n11145));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1072_25.INIT0 = 16'h5999;
    defparam add_1072_25.INIT1 = 16'h5999;
    defparam add_1072_25.INJECT1_0 = "NO";
    defparam add_1072_25.INJECT1_1 = "NO";
    CCU2D add_1072_23 (.A0(d9[21]), .B0(d_d9[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[22]), .B1(d_d9[22]), .C1(GND_net), .D1(GND_net), .CIN(n11143), 
          .COUT(n11144));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1072_23.INIT0 = 16'h5999;
    defparam add_1072_23.INIT1 = 16'h5999;
    defparam add_1072_23.INJECT1_0 = "NO";
    defparam add_1072_23.INJECT1_1 = "NO";
    CCU2D add_1072_21 (.A0(d9[19]), .B0(d_d9[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[20]), .B1(d_d9[20]), .C1(GND_net), .D1(GND_net), .CIN(n11142), 
          .COUT(n11143));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1072_21.INIT0 = 16'h5999;
    defparam add_1072_21.INIT1 = 16'h5999;
    defparam add_1072_21.INJECT1_0 = "NO";
    defparam add_1072_21.INJECT1_1 = "NO";
    CCU2D add_1072_19 (.A0(d9[17]), .B0(d_d9[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[18]), .B1(d_d9[18]), .C1(GND_net), .D1(GND_net), .CIN(n11141), 
          .COUT(n11142));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1072_19.INIT0 = 16'h5999;
    defparam add_1072_19.INIT1 = 16'h5999;
    defparam add_1072_19.INJECT1_0 = "NO";
    defparam add_1072_19.INJECT1_1 = "NO";
    CCU2D add_1072_17 (.A0(d9[15]), .B0(d_d9[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[16]), .B1(d_d9[16]), .C1(GND_net), .D1(GND_net), .CIN(n11140), 
          .COUT(n11141));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1072_17.INIT0 = 16'h5999;
    defparam add_1072_17.INIT1 = 16'h5999;
    defparam add_1072_17.INJECT1_0 = "NO";
    defparam add_1072_17.INJECT1_1 = "NO";
    CCU2D add_1072_15 (.A0(d9[13]), .B0(d_d9[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[14]), .B1(d_d9[14]), .C1(GND_net), .D1(GND_net), .CIN(n11139), 
          .COUT(n11140));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1072_15.INIT0 = 16'h5999;
    defparam add_1072_15.INIT1 = 16'h5999;
    defparam add_1072_15.INJECT1_0 = "NO";
    defparam add_1072_15.INJECT1_1 = "NO";
    CCU2D add_1072_13 (.A0(d9[11]), .B0(d_d9[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[12]), .B1(d_d9[12]), .C1(GND_net), .D1(GND_net), .CIN(n11138), 
          .COUT(n11139));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1072_13.INIT0 = 16'h5999;
    defparam add_1072_13.INIT1 = 16'h5999;
    defparam add_1072_13.INJECT1_0 = "NO";
    defparam add_1072_13.INJECT1_1 = "NO";
    CCU2D add_1072_11 (.A0(d9[9]), .B0(d_d9[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[10]), .B1(d_d9[10]), .C1(GND_net), .D1(GND_net), .CIN(n11137), 
          .COUT(n11138));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1072_11.INIT0 = 16'h5999;
    defparam add_1072_11.INIT1 = 16'h5999;
    defparam add_1072_11.INJECT1_0 = "NO";
    defparam add_1072_11.INJECT1_1 = "NO";
    CCU2D add_1072_9 (.A0(d9[7]), .B0(d_d9[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[8]), .B1(d_d9[8]), .C1(GND_net), .D1(GND_net), .CIN(n11136), 
          .COUT(n11137));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1072_9.INIT0 = 16'h5999;
    defparam add_1072_9.INIT1 = 16'h5999;
    defparam add_1072_9.INJECT1_0 = "NO";
    defparam add_1072_9.INJECT1_1 = "NO";
    CCU2D add_1072_7 (.A0(d9[5]), .B0(d_d9[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[6]), .B1(d_d9[6]), .C1(GND_net), .D1(GND_net), .CIN(n11135), 
          .COUT(n11136));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1072_7.INIT0 = 16'h5999;
    defparam add_1072_7.INIT1 = 16'h5999;
    defparam add_1072_7.INJECT1_0 = "NO";
    defparam add_1072_7.INJECT1_1 = "NO";
    CCU2D add_1072_5 (.A0(d9[3]), .B0(d_d9[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[4]), .B1(d_d9[4]), .C1(GND_net), .D1(GND_net), .CIN(n11134), 
          .COUT(n11135));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1072_5.INIT0 = 16'h5999;
    defparam add_1072_5.INIT1 = 16'h5999;
    defparam add_1072_5.INJECT1_0 = "NO";
    defparam add_1072_5.INJECT1_1 = "NO";
    CCU2D add_1072_3 (.A0(d9[1]), .B0(d_d9[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d9[2]), .B1(d_d9[2]), .C1(GND_net), .D1(GND_net), .CIN(n11133), 
          .COUT(n11134));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1072_3.INIT0 = 16'h5999;
    defparam add_1072_3.INIT1 = 16'h5999;
    defparam add_1072_3.INJECT1_0 = "NO";
    defparam add_1072_3.INJECT1_1 = "NO";
    CCU2D add_1072_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d9[0]), .B1(d_d9[0]), .C1(GND_net), .D1(GND_net), .COUT(n11133));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam add_1072_1.INIT0 = 16'h0000;
    defparam add_1072_1.INIT1 = 16'h5999;
    defparam add_1072_1.INJECT1_0 = "NO";
    defparam add_1072_1.INJECT1_1 = "NO";
    CCU2D add_1067_37 (.A0(d8[35]), .B0(d_d8[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11132), 
          .S0(d9_71__N_1674[35]), .S1(n6622));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1067_37.INIT0 = 16'h5999;
    defparam add_1067_37.INIT1 = 16'h0000;
    defparam add_1067_37.INJECT1_0 = "NO";
    defparam add_1067_37.INJECT1_1 = "NO";
    CCU2D add_1067_35 (.A0(d8[33]), .B0(d_d8[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[34]), .B1(d_d8[34]), .C1(GND_net), .D1(GND_net), .CIN(n11131), 
          .COUT(n11132), .S0(d9_71__N_1674[33]), .S1(d9_71__N_1674[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1067_35.INIT0 = 16'h5999;
    defparam add_1067_35.INIT1 = 16'h5999;
    defparam add_1067_35.INJECT1_0 = "NO";
    defparam add_1067_35.INJECT1_1 = "NO";
    CCU2D add_1067_33 (.A0(d8[31]), .B0(d_d8[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[32]), .B1(d_d8[32]), .C1(GND_net), .D1(GND_net), .CIN(n11130), 
          .COUT(n11131), .S0(d9_71__N_1674[31]), .S1(d9_71__N_1674[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1067_33.INIT0 = 16'h5999;
    defparam add_1067_33.INIT1 = 16'h5999;
    defparam add_1067_33.INJECT1_0 = "NO";
    defparam add_1067_33.INJECT1_1 = "NO";
    CCU2D add_1067_31 (.A0(d8[29]), .B0(d_d8[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[30]), .B1(d_d8[30]), .C1(GND_net), .D1(GND_net), .CIN(n11129), 
          .COUT(n11130), .S0(d9_71__N_1674[29]), .S1(d9_71__N_1674[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1067_31.INIT0 = 16'h5999;
    defparam add_1067_31.INIT1 = 16'h5999;
    defparam add_1067_31.INJECT1_0 = "NO";
    defparam add_1067_31.INJECT1_1 = "NO";
    CCU2D add_1067_29 (.A0(d8[27]), .B0(d_d8[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[28]), .B1(d_d8[28]), .C1(GND_net), .D1(GND_net), .CIN(n11128), 
          .COUT(n11129), .S0(d9_71__N_1674[27]), .S1(d9_71__N_1674[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1067_29.INIT0 = 16'h5999;
    defparam add_1067_29.INIT1 = 16'h5999;
    defparam add_1067_29.INJECT1_0 = "NO";
    defparam add_1067_29.INJECT1_1 = "NO";
    CCU2D add_1067_27 (.A0(d8[25]), .B0(d_d8[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[26]), .B1(d_d8[26]), .C1(GND_net), .D1(GND_net), .CIN(n11127), 
          .COUT(n11128), .S0(d9_71__N_1674[25]), .S1(d9_71__N_1674[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1067_27.INIT0 = 16'h5999;
    defparam add_1067_27.INIT1 = 16'h5999;
    defparam add_1067_27.INJECT1_0 = "NO";
    defparam add_1067_27.INJECT1_1 = "NO";
    CCU2D add_1067_25 (.A0(d8[23]), .B0(d_d8[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[24]), .B1(d_d8[24]), .C1(GND_net), .D1(GND_net), .CIN(n11126), 
          .COUT(n11127), .S0(d9_71__N_1674[23]), .S1(d9_71__N_1674[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1067_25.INIT0 = 16'h5999;
    defparam add_1067_25.INIT1 = 16'h5999;
    defparam add_1067_25.INJECT1_0 = "NO";
    defparam add_1067_25.INJECT1_1 = "NO";
    CCU2D add_1067_23 (.A0(d8[21]), .B0(d_d8[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[22]), .B1(d_d8[22]), .C1(GND_net), .D1(GND_net), .CIN(n11125), 
          .COUT(n11126), .S0(d9_71__N_1674[21]), .S1(d9_71__N_1674[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1067_23.INIT0 = 16'h5999;
    defparam add_1067_23.INIT1 = 16'h5999;
    defparam add_1067_23.INJECT1_0 = "NO";
    defparam add_1067_23.INJECT1_1 = "NO";
    CCU2D add_1067_21 (.A0(d8[19]), .B0(d_d8[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[20]), .B1(d_d8[20]), .C1(GND_net), .D1(GND_net), .CIN(n11124), 
          .COUT(n11125), .S0(d9_71__N_1674[19]), .S1(d9_71__N_1674[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1067_21.INIT0 = 16'h5999;
    defparam add_1067_21.INIT1 = 16'h5999;
    defparam add_1067_21.INJECT1_0 = "NO";
    defparam add_1067_21.INJECT1_1 = "NO";
    CCU2D add_1067_19 (.A0(d8[17]), .B0(d_d8[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[18]), .B1(d_d8[18]), .C1(GND_net), .D1(GND_net), .CIN(n11123), 
          .COUT(n11124), .S0(d9_71__N_1674[17]), .S1(d9_71__N_1674[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1067_19.INIT0 = 16'h5999;
    defparam add_1067_19.INIT1 = 16'h5999;
    defparam add_1067_19.INJECT1_0 = "NO";
    defparam add_1067_19.INJECT1_1 = "NO";
    CCU2D add_1067_17 (.A0(d8[15]), .B0(d_d8[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[16]), .B1(d_d8[16]), .C1(GND_net), .D1(GND_net), .CIN(n11122), 
          .COUT(n11123), .S0(d9_71__N_1674[15]), .S1(d9_71__N_1674[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1067_17.INIT0 = 16'h5999;
    defparam add_1067_17.INIT1 = 16'h5999;
    defparam add_1067_17.INJECT1_0 = "NO";
    defparam add_1067_17.INJECT1_1 = "NO";
    CCU2D add_1067_15 (.A0(d8[13]), .B0(d_d8[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[14]), .B1(d_d8[14]), .C1(GND_net), .D1(GND_net), .CIN(n11121), 
          .COUT(n11122), .S0(d9_71__N_1674[13]), .S1(d9_71__N_1674[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1067_15.INIT0 = 16'h5999;
    defparam add_1067_15.INIT1 = 16'h5999;
    defparam add_1067_15.INJECT1_0 = "NO";
    defparam add_1067_15.INJECT1_1 = "NO";
    CCU2D add_1067_13 (.A0(d8[11]), .B0(d_d8[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[12]), .B1(d_d8[12]), .C1(GND_net), .D1(GND_net), .CIN(n11120), 
          .COUT(n11121), .S0(d9_71__N_1674[11]), .S1(d9_71__N_1674[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1067_13.INIT0 = 16'h5999;
    defparam add_1067_13.INIT1 = 16'h5999;
    defparam add_1067_13.INJECT1_0 = "NO";
    defparam add_1067_13.INJECT1_1 = "NO";
    CCU2D add_1067_11 (.A0(d8[9]), .B0(d_d8[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[10]), .B1(d_d8[10]), .C1(GND_net), .D1(GND_net), .CIN(n11119), 
          .COUT(n11120), .S0(d9_71__N_1674[9]), .S1(d9_71__N_1674[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1067_11.INIT0 = 16'h5999;
    defparam add_1067_11.INIT1 = 16'h5999;
    defparam add_1067_11.INJECT1_0 = "NO";
    defparam add_1067_11.INJECT1_1 = "NO";
    CCU2D add_1067_9 (.A0(d8[7]), .B0(d_d8[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[8]), .B1(d_d8[8]), .C1(GND_net), .D1(GND_net), .CIN(n11118), 
          .COUT(n11119), .S0(d9_71__N_1674[7]), .S1(d9_71__N_1674[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1067_9.INIT0 = 16'h5999;
    defparam add_1067_9.INIT1 = 16'h5999;
    defparam add_1067_9.INJECT1_0 = "NO";
    defparam add_1067_9.INJECT1_1 = "NO";
    CCU2D add_1067_7 (.A0(d8[5]), .B0(d_d8[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[6]), .B1(d_d8[6]), .C1(GND_net), .D1(GND_net), .CIN(n11117), 
          .COUT(n11118), .S0(d9_71__N_1674[5]), .S1(d9_71__N_1674[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1067_7.INIT0 = 16'h5999;
    defparam add_1067_7.INIT1 = 16'h5999;
    defparam add_1067_7.INJECT1_0 = "NO";
    defparam add_1067_7.INJECT1_1 = "NO";
    CCU2D add_1067_5 (.A0(d8[3]), .B0(d_d8[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[4]), .B1(d_d8[4]), .C1(GND_net), .D1(GND_net), .CIN(n11116), 
          .COUT(n11117), .S0(d9_71__N_1674[3]), .S1(d9_71__N_1674[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1067_5.INIT0 = 16'h5999;
    defparam add_1067_5.INIT1 = 16'h5999;
    defparam add_1067_5.INJECT1_0 = "NO";
    defparam add_1067_5.INJECT1_1 = "NO";
    CCU2D add_1067_3 (.A0(d8[1]), .B0(d_d8[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d8[2]), .B1(d_d8[2]), .C1(GND_net), .D1(GND_net), .CIN(n11115), 
          .COUT(n11116), .S0(d9_71__N_1674[1]), .S1(d9_71__N_1674[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1067_3.INIT0 = 16'h5999;
    defparam add_1067_3.INIT1 = 16'h5999;
    defparam add_1067_3.INJECT1_0 = "NO";
    defparam add_1067_3.INJECT1_1 = "NO";
    CCU2D add_1067_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d8[0]), .B1(d_d8[0]), .C1(GND_net), .D1(GND_net), .COUT(n11115), 
          .S1(d9_71__N_1674[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(112[17:26])
    defparam add_1067_1.INIT0 = 16'h0000;
    defparam add_1067_1.INIT1 = 16'h5999;
    defparam add_1067_1.INJECT1_0 = "NO";
    defparam add_1067_1.INJECT1_1 = "NO";
    CCU2D add_1052_37 (.A0(d_tmp[35]), .B0(d_d_tmp[35]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11073), .S0(d6_71__N_1458[35]), .S1(n6166));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1052_37.INIT0 = 16'h5999;
    defparam add_1052_37.INIT1 = 16'h0000;
    defparam add_1052_37.INJECT1_0 = "NO";
    defparam add_1052_37.INJECT1_1 = "NO";
    CCU2D add_1052_35 (.A0(d_tmp[33]), .B0(d_d_tmp[33]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[34]), .B1(d_d_tmp[34]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11072), .COUT(n11073), .S0(d6_71__N_1458[33]), 
          .S1(d6_71__N_1458[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1052_35.INIT0 = 16'h5999;
    defparam add_1052_35.INIT1 = 16'h5999;
    defparam add_1052_35.INJECT1_0 = "NO";
    defparam add_1052_35.INJECT1_1 = "NO";
    CCU2D add_1052_33 (.A0(d_tmp[31]), .B0(d_d_tmp[31]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[32]), .B1(d_d_tmp[32]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11071), .COUT(n11072), .S0(d6_71__N_1458[31]), 
          .S1(d6_71__N_1458[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1052_33.INIT0 = 16'h5999;
    defparam add_1052_33.INIT1 = 16'h5999;
    defparam add_1052_33.INJECT1_0 = "NO";
    defparam add_1052_33.INJECT1_1 = "NO";
    CCU2D add_1052_31 (.A0(d_tmp[29]), .B0(d_d_tmp[29]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[30]), .B1(d_d_tmp[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11070), .COUT(n11071), .S0(d6_71__N_1458[29]), 
          .S1(d6_71__N_1458[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1052_31.INIT0 = 16'h5999;
    defparam add_1052_31.INIT1 = 16'h5999;
    defparam add_1052_31.INJECT1_0 = "NO";
    defparam add_1052_31.INJECT1_1 = "NO";
    CCU2D add_1052_29 (.A0(d_tmp[27]), .B0(d_d_tmp[27]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[28]), .B1(d_d_tmp[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11069), .COUT(n11070), .S0(d6_71__N_1458[27]), 
          .S1(d6_71__N_1458[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1052_29.INIT0 = 16'h5999;
    defparam add_1052_29.INIT1 = 16'h5999;
    defparam add_1052_29.INJECT1_0 = "NO";
    defparam add_1052_29.INJECT1_1 = "NO";
    CCU2D add_1052_27 (.A0(d_tmp[25]), .B0(d_d_tmp[25]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[26]), .B1(d_d_tmp[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11068), .COUT(n11069), .S0(d6_71__N_1458[25]), 
          .S1(d6_71__N_1458[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1052_27.INIT0 = 16'h5999;
    defparam add_1052_27.INIT1 = 16'h5999;
    defparam add_1052_27.INJECT1_0 = "NO";
    defparam add_1052_27.INJECT1_1 = "NO";
    CCU2D add_1052_25 (.A0(d_tmp[23]), .B0(d_d_tmp[23]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[24]), .B1(d_d_tmp[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11067), .COUT(n11068), .S0(d6_71__N_1458[23]), 
          .S1(d6_71__N_1458[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1052_25.INIT0 = 16'h5999;
    defparam add_1052_25.INIT1 = 16'h5999;
    defparam add_1052_25.INJECT1_0 = "NO";
    defparam add_1052_25.INJECT1_1 = "NO";
    CCU2D add_1052_23 (.A0(d_tmp[21]), .B0(d_d_tmp[21]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[22]), .B1(d_d_tmp[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11066), .COUT(n11067), .S0(d6_71__N_1458[21]), 
          .S1(d6_71__N_1458[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1052_23.INIT0 = 16'h5999;
    defparam add_1052_23.INIT1 = 16'h5999;
    defparam add_1052_23.INJECT1_0 = "NO";
    defparam add_1052_23.INJECT1_1 = "NO";
    CCU2D add_1052_21 (.A0(d_tmp[19]), .B0(d_d_tmp[19]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[20]), .B1(d_d_tmp[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11065), .COUT(n11066), .S0(d6_71__N_1458[19]), 
          .S1(d6_71__N_1458[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1052_21.INIT0 = 16'h5999;
    defparam add_1052_21.INIT1 = 16'h5999;
    defparam add_1052_21.INJECT1_0 = "NO";
    defparam add_1052_21.INJECT1_1 = "NO";
    CCU2D add_1052_19 (.A0(d_tmp[17]), .B0(d_d_tmp[17]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[18]), .B1(d_d_tmp[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11064), .COUT(n11065), .S0(d6_71__N_1458[17]), 
          .S1(d6_71__N_1458[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1052_19.INIT0 = 16'h5999;
    defparam add_1052_19.INIT1 = 16'h5999;
    defparam add_1052_19.INJECT1_0 = "NO";
    defparam add_1052_19.INJECT1_1 = "NO";
    CCU2D add_1052_17 (.A0(d_tmp[15]), .B0(d_d_tmp[15]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[16]), .B1(d_d_tmp[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11063), .COUT(n11064), .S0(d6_71__N_1458[15]), 
          .S1(d6_71__N_1458[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1052_17.INIT0 = 16'h5999;
    defparam add_1052_17.INIT1 = 16'h5999;
    defparam add_1052_17.INJECT1_0 = "NO";
    defparam add_1052_17.INJECT1_1 = "NO";
    CCU2D add_1052_15 (.A0(d_tmp[13]), .B0(d_d_tmp[13]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[14]), .B1(d_d_tmp[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11062), .COUT(n11063), .S0(d6_71__N_1458[13]), 
          .S1(d6_71__N_1458[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1052_15.INIT0 = 16'h5999;
    defparam add_1052_15.INIT1 = 16'h5999;
    defparam add_1052_15.INJECT1_0 = "NO";
    defparam add_1052_15.INJECT1_1 = "NO";
    CCU2D add_1052_13 (.A0(d_tmp[11]), .B0(d_d_tmp[11]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[12]), .B1(d_d_tmp[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11061), .COUT(n11062), .S0(d6_71__N_1458[11]), 
          .S1(d6_71__N_1458[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1052_13.INIT0 = 16'h5999;
    defparam add_1052_13.INIT1 = 16'h5999;
    defparam add_1052_13.INJECT1_0 = "NO";
    defparam add_1052_13.INJECT1_1 = "NO";
    CCU2D add_1052_11 (.A0(d_tmp[9]), .B0(d_d_tmp[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[10]), .B1(d_d_tmp[10]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11060), .COUT(n11061), .S0(d6_71__N_1458[9]), .S1(d6_71__N_1458[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1052_11.INIT0 = 16'h5999;
    defparam add_1052_11.INIT1 = 16'h5999;
    defparam add_1052_11.INJECT1_0 = "NO";
    defparam add_1052_11.INJECT1_1 = "NO";
    CCU2D add_1052_9 (.A0(d_tmp[7]), .B0(d_d_tmp[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[8]), .B1(d_d_tmp[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11059), .COUT(n11060), .S0(d6_71__N_1458[7]), .S1(d6_71__N_1458[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1052_9.INIT0 = 16'h5999;
    defparam add_1052_9.INIT1 = 16'h5999;
    defparam add_1052_9.INJECT1_0 = "NO";
    defparam add_1052_9.INJECT1_1 = "NO";
    CCU2D add_1052_7 (.A0(d_tmp[5]), .B0(d_d_tmp[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[6]), .B1(d_d_tmp[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11058), .COUT(n11059), .S0(d6_71__N_1458[5]), .S1(d6_71__N_1458[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1052_7.INIT0 = 16'h5999;
    defparam add_1052_7.INIT1 = 16'h5999;
    defparam add_1052_7.INJECT1_0 = "NO";
    defparam add_1052_7.INJECT1_1 = "NO";
    CCU2D add_1052_5 (.A0(d_tmp[3]), .B0(d_d_tmp[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[4]), .B1(d_d_tmp[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11057), .COUT(n11058), .S0(d6_71__N_1458[3]), .S1(d6_71__N_1458[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1052_5.INIT0 = 16'h5999;
    defparam add_1052_5.INIT1 = 16'h5999;
    defparam add_1052_5.INJECT1_0 = "NO";
    defparam add_1052_5.INJECT1_1 = "NO";
    CCU2D add_1052_3 (.A0(d_tmp[1]), .B0(d_d_tmp[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[2]), .B1(d_d_tmp[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n11056), .COUT(n11057), .S0(d6_71__N_1458[1]), .S1(d6_71__N_1458[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1052_3.INIT0 = 16'h5999;
    defparam add_1052_3.INIT1 = 16'h5999;
    defparam add_1052_3.INJECT1_0 = "NO";
    defparam add_1052_3.INJECT1_1 = "NO";
    CCU2D add_1052_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_tmp[0]), .B1(d_d_tmp[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n11056), .S1(d6_71__N_1458[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1052_1.INIT0 = 16'h0000;
    defparam add_1052_1.INIT1 = 16'h5999;
    defparam add_1052_1.INJECT1_0 = "NO";
    defparam add_1052_1.INJECT1_1 = "NO";
    CCU2D add_1047_37 (.A0(d6[35]), .B0(d_d6[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11055), 
          .S0(d7_71__N_1530[35]), .S1(n6014));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1047_37.INIT0 = 16'h5999;
    defparam add_1047_37.INIT1 = 16'h0000;
    defparam add_1047_37.INJECT1_0 = "NO";
    defparam add_1047_37.INJECT1_1 = "NO";
    CCU2D add_1047_35 (.A0(d6[33]), .B0(d_d6[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[34]), .B1(d_d6[34]), .C1(GND_net), .D1(GND_net), .CIN(n11054), 
          .COUT(n11055), .S0(d7_71__N_1530[33]), .S1(d7_71__N_1530[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1047_35.INIT0 = 16'h5999;
    defparam add_1047_35.INIT1 = 16'h5999;
    defparam add_1047_35.INJECT1_0 = "NO";
    defparam add_1047_35.INJECT1_1 = "NO";
    CCU2D add_1047_33 (.A0(d6[31]), .B0(d_d6[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[32]), .B1(d_d6[32]), .C1(GND_net), .D1(GND_net), .CIN(n11053), 
          .COUT(n11054), .S0(d7_71__N_1530[31]), .S1(d7_71__N_1530[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1047_33.INIT0 = 16'h5999;
    defparam add_1047_33.INIT1 = 16'h5999;
    defparam add_1047_33.INJECT1_0 = "NO";
    defparam add_1047_33.INJECT1_1 = "NO";
    CCU2D add_1047_31 (.A0(d6[29]), .B0(d_d6[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[30]), .B1(d_d6[30]), .C1(GND_net), .D1(GND_net), .CIN(n11052), 
          .COUT(n11053), .S0(d7_71__N_1530[29]), .S1(d7_71__N_1530[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1047_31.INIT0 = 16'h5999;
    defparam add_1047_31.INIT1 = 16'h5999;
    defparam add_1047_31.INJECT1_0 = "NO";
    defparam add_1047_31.INJECT1_1 = "NO";
    CCU2D add_1047_29 (.A0(d6[27]), .B0(d_d6[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[28]), .B1(d_d6[28]), .C1(GND_net), .D1(GND_net), .CIN(n11051), 
          .COUT(n11052), .S0(d7_71__N_1530[27]), .S1(d7_71__N_1530[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1047_29.INIT0 = 16'h5999;
    defparam add_1047_29.INIT1 = 16'h5999;
    defparam add_1047_29.INJECT1_0 = "NO";
    defparam add_1047_29.INJECT1_1 = "NO";
    CCU2D add_1047_27 (.A0(d6[25]), .B0(d_d6[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[26]), .B1(d_d6[26]), .C1(GND_net), .D1(GND_net), .CIN(n11050), 
          .COUT(n11051), .S0(d7_71__N_1530[25]), .S1(d7_71__N_1530[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1047_27.INIT0 = 16'h5999;
    defparam add_1047_27.INIT1 = 16'h5999;
    defparam add_1047_27.INJECT1_0 = "NO";
    defparam add_1047_27.INJECT1_1 = "NO";
    CCU2D add_1047_25 (.A0(d6[23]), .B0(d_d6[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[24]), .B1(d_d6[24]), .C1(GND_net), .D1(GND_net), .CIN(n11049), 
          .COUT(n11050), .S0(d7_71__N_1530[23]), .S1(d7_71__N_1530[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1047_25.INIT0 = 16'h5999;
    defparam add_1047_25.INIT1 = 16'h5999;
    defparam add_1047_25.INJECT1_0 = "NO";
    defparam add_1047_25.INJECT1_1 = "NO";
    CCU2D add_1047_23 (.A0(d6[21]), .B0(d_d6[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[22]), .B1(d_d6[22]), .C1(GND_net), .D1(GND_net), .CIN(n11048), 
          .COUT(n11049), .S0(d7_71__N_1530[21]), .S1(d7_71__N_1530[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1047_23.INIT0 = 16'h5999;
    defparam add_1047_23.INIT1 = 16'h5999;
    defparam add_1047_23.INJECT1_0 = "NO";
    defparam add_1047_23.INJECT1_1 = "NO";
    CCU2D add_1047_21 (.A0(d6[19]), .B0(d_d6[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[20]), .B1(d_d6[20]), .C1(GND_net), .D1(GND_net), .CIN(n11047), 
          .COUT(n11048), .S0(d7_71__N_1530[19]), .S1(d7_71__N_1530[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1047_21.INIT0 = 16'h5999;
    defparam add_1047_21.INIT1 = 16'h5999;
    defparam add_1047_21.INJECT1_0 = "NO";
    defparam add_1047_21.INJECT1_1 = "NO";
    CCU2D add_1047_19 (.A0(d6[17]), .B0(d_d6[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[18]), .B1(d_d6[18]), .C1(GND_net), .D1(GND_net), .CIN(n11046), 
          .COUT(n11047), .S0(d7_71__N_1530[17]), .S1(d7_71__N_1530[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1047_19.INIT0 = 16'h5999;
    defparam add_1047_19.INIT1 = 16'h5999;
    defparam add_1047_19.INJECT1_0 = "NO";
    defparam add_1047_19.INJECT1_1 = "NO";
    CCU2D add_1047_17 (.A0(d6[15]), .B0(d_d6[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[16]), .B1(d_d6[16]), .C1(GND_net), .D1(GND_net), .CIN(n11045), 
          .COUT(n11046), .S0(d7_71__N_1530[15]), .S1(d7_71__N_1530[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1047_17.INIT0 = 16'h5999;
    defparam add_1047_17.INIT1 = 16'h5999;
    defparam add_1047_17.INJECT1_0 = "NO";
    defparam add_1047_17.INJECT1_1 = "NO";
    CCU2D add_1047_15 (.A0(d6[13]), .B0(d_d6[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[14]), .B1(d_d6[14]), .C1(GND_net), .D1(GND_net), .CIN(n11044), 
          .COUT(n11045), .S0(d7_71__N_1530[13]), .S1(d7_71__N_1530[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1047_15.INIT0 = 16'h5999;
    defparam add_1047_15.INIT1 = 16'h5999;
    defparam add_1047_15.INJECT1_0 = "NO";
    defparam add_1047_15.INJECT1_1 = "NO";
    CCU2D add_1047_13 (.A0(d6[11]), .B0(d_d6[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[12]), .B1(d_d6[12]), .C1(GND_net), .D1(GND_net), .CIN(n11043), 
          .COUT(n11044), .S0(d7_71__N_1530[11]), .S1(d7_71__N_1530[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1047_13.INIT0 = 16'h5999;
    defparam add_1047_13.INIT1 = 16'h5999;
    defparam add_1047_13.INJECT1_0 = "NO";
    defparam add_1047_13.INJECT1_1 = "NO";
    CCU2D add_1047_11 (.A0(d6[9]), .B0(d_d6[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[10]), .B1(d_d6[10]), .C1(GND_net), .D1(GND_net), .CIN(n11042), 
          .COUT(n11043), .S0(d7_71__N_1530[9]), .S1(d7_71__N_1530[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1047_11.INIT0 = 16'h5999;
    defparam add_1047_11.INIT1 = 16'h5999;
    defparam add_1047_11.INJECT1_0 = "NO";
    defparam add_1047_11.INJECT1_1 = "NO";
    CCU2D add_1047_9 (.A0(d6[7]), .B0(d_d6[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[8]), .B1(d_d6[8]), .C1(GND_net), .D1(GND_net), .CIN(n11041), 
          .COUT(n11042), .S0(d7_71__N_1530[7]), .S1(d7_71__N_1530[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1047_9.INIT0 = 16'h5999;
    defparam add_1047_9.INIT1 = 16'h5999;
    defparam add_1047_9.INJECT1_0 = "NO";
    defparam add_1047_9.INJECT1_1 = "NO";
    CCU2D add_1047_7 (.A0(d6[5]), .B0(d_d6[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[6]), .B1(d_d6[6]), .C1(GND_net), .D1(GND_net), .CIN(n11040), 
          .COUT(n11041), .S0(d7_71__N_1530[5]), .S1(d7_71__N_1530[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1047_7.INIT0 = 16'h5999;
    defparam add_1047_7.INIT1 = 16'h5999;
    defparam add_1047_7.INJECT1_0 = "NO";
    defparam add_1047_7.INJECT1_1 = "NO";
    CCU2D add_1047_5 (.A0(d6[3]), .B0(d_d6[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[4]), .B1(d_d6[4]), .C1(GND_net), .D1(GND_net), .CIN(n11039), 
          .COUT(n11040), .S0(d7_71__N_1530[3]), .S1(d7_71__N_1530[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1047_5.INIT0 = 16'h5999;
    defparam add_1047_5.INIT1 = 16'h5999;
    defparam add_1047_5.INJECT1_0 = "NO";
    defparam add_1047_5.INJECT1_1 = "NO";
    CCU2D add_1047_3 (.A0(d6[1]), .B0(d_d6[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[2]), .B1(d_d6[2]), .C1(GND_net), .D1(GND_net), .CIN(n11038), 
          .COUT(n11039), .S0(d7_71__N_1530[1]), .S1(d7_71__N_1530[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1047_3.INIT0 = 16'h5999;
    defparam add_1047_3.INIT1 = 16'h5999;
    defparam add_1047_3.INJECT1_0 = "NO";
    defparam add_1047_3.INJECT1_1 = "NO";
    CCU2D add_1047_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d6[0]), .B1(d_d6[0]), .C1(GND_net), .D1(GND_net), .COUT(n11038), 
          .S1(d7_71__N_1530[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1047_1.INIT0 = 16'h0000;
    defparam add_1047_1.INIT1 = 16'h5999;
    defparam add_1047_1.INJECT1_0 = "NO";
    defparam add_1047_1.INJECT1_1 = "NO";
    CCU2D add_1042_37 (.A0(d7[35]), .B0(d_d7[35]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11037), 
          .S0(d8_71__N_1602[35]), .S1(n5862));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1042_37.INIT0 = 16'h5999;
    defparam add_1042_37.INIT1 = 16'h0000;
    defparam add_1042_37.INJECT1_0 = "NO";
    defparam add_1042_37.INJECT1_1 = "NO";
    CCU2D add_1042_35 (.A0(d7[33]), .B0(d_d7[33]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[34]), .B1(d_d7[34]), .C1(GND_net), .D1(GND_net), .CIN(n11036), 
          .COUT(n11037), .S0(d8_71__N_1602[33]), .S1(d8_71__N_1602[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1042_35.INIT0 = 16'h5999;
    defparam add_1042_35.INIT1 = 16'h5999;
    defparam add_1042_35.INJECT1_0 = "NO";
    defparam add_1042_35.INJECT1_1 = "NO";
    CCU2D add_1042_33 (.A0(d7[31]), .B0(d_d7[31]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[32]), .B1(d_d7[32]), .C1(GND_net), .D1(GND_net), .CIN(n11035), 
          .COUT(n11036), .S0(d8_71__N_1602[31]), .S1(d8_71__N_1602[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1042_33.INIT0 = 16'h5999;
    defparam add_1042_33.INIT1 = 16'h5999;
    defparam add_1042_33.INJECT1_0 = "NO";
    defparam add_1042_33.INJECT1_1 = "NO";
    CCU2D add_1042_31 (.A0(d7[29]), .B0(d_d7[29]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[30]), .B1(d_d7[30]), .C1(GND_net), .D1(GND_net), .CIN(n11034), 
          .COUT(n11035), .S0(d8_71__N_1602[29]), .S1(d8_71__N_1602[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1042_31.INIT0 = 16'h5999;
    defparam add_1042_31.INIT1 = 16'h5999;
    defparam add_1042_31.INJECT1_0 = "NO";
    defparam add_1042_31.INJECT1_1 = "NO";
    CCU2D add_1042_29 (.A0(d7[27]), .B0(d_d7[27]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[28]), .B1(d_d7[28]), .C1(GND_net), .D1(GND_net), .CIN(n11033), 
          .COUT(n11034), .S0(d8_71__N_1602[27]), .S1(d8_71__N_1602[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1042_29.INIT0 = 16'h5999;
    defparam add_1042_29.INIT1 = 16'h5999;
    defparam add_1042_29.INJECT1_0 = "NO";
    defparam add_1042_29.INJECT1_1 = "NO";
    CCU2D add_1042_27 (.A0(d7[25]), .B0(d_d7[25]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[26]), .B1(d_d7[26]), .C1(GND_net), .D1(GND_net), .CIN(n11032), 
          .COUT(n11033), .S0(d8_71__N_1602[25]), .S1(d8_71__N_1602[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1042_27.INIT0 = 16'h5999;
    defparam add_1042_27.INIT1 = 16'h5999;
    defparam add_1042_27.INJECT1_0 = "NO";
    defparam add_1042_27.INJECT1_1 = "NO";
    CCU2D add_1042_25 (.A0(d7[23]), .B0(d_d7[23]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[24]), .B1(d_d7[24]), .C1(GND_net), .D1(GND_net), .CIN(n11031), 
          .COUT(n11032), .S0(d8_71__N_1602[23]), .S1(d8_71__N_1602[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1042_25.INIT0 = 16'h5999;
    defparam add_1042_25.INIT1 = 16'h5999;
    defparam add_1042_25.INJECT1_0 = "NO";
    defparam add_1042_25.INJECT1_1 = "NO";
    CCU2D add_1042_23 (.A0(d7[21]), .B0(d_d7[21]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[22]), .B1(d_d7[22]), .C1(GND_net), .D1(GND_net), .CIN(n11030), 
          .COUT(n11031), .S0(d8_71__N_1602[21]), .S1(d8_71__N_1602[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1042_23.INIT0 = 16'h5999;
    defparam add_1042_23.INIT1 = 16'h5999;
    defparam add_1042_23.INJECT1_0 = "NO";
    defparam add_1042_23.INJECT1_1 = "NO";
    CCU2D add_1042_21 (.A0(d7[19]), .B0(d_d7[19]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[20]), .B1(d_d7[20]), .C1(GND_net), .D1(GND_net), .CIN(n11029), 
          .COUT(n11030), .S0(d8_71__N_1602[19]), .S1(d8_71__N_1602[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1042_21.INIT0 = 16'h5999;
    defparam add_1042_21.INIT1 = 16'h5999;
    defparam add_1042_21.INJECT1_0 = "NO";
    defparam add_1042_21.INJECT1_1 = "NO";
    CCU2D add_1042_19 (.A0(d7[17]), .B0(d_d7[17]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[18]), .B1(d_d7[18]), .C1(GND_net), .D1(GND_net), .CIN(n11028), 
          .COUT(n11029), .S0(d8_71__N_1602[17]), .S1(d8_71__N_1602[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1042_19.INIT0 = 16'h5999;
    defparam add_1042_19.INIT1 = 16'h5999;
    defparam add_1042_19.INJECT1_0 = "NO";
    defparam add_1042_19.INJECT1_1 = "NO";
    CCU2D add_1042_17 (.A0(d7[15]), .B0(d_d7[15]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[16]), .B1(d_d7[16]), .C1(GND_net), .D1(GND_net), .CIN(n11027), 
          .COUT(n11028), .S0(d8_71__N_1602[15]), .S1(d8_71__N_1602[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1042_17.INIT0 = 16'h5999;
    defparam add_1042_17.INIT1 = 16'h5999;
    defparam add_1042_17.INJECT1_0 = "NO";
    defparam add_1042_17.INJECT1_1 = "NO";
    CCU2D add_1042_15 (.A0(d7[13]), .B0(d_d7[13]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[14]), .B1(d_d7[14]), .C1(GND_net), .D1(GND_net), .CIN(n11026), 
          .COUT(n11027), .S0(d8_71__N_1602[13]), .S1(d8_71__N_1602[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1042_15.INIT0 = 16'h5999;
    defparam add_1042_15.INIT1 = 16'h5999;
    defparam add_1042_15.INJECT1_0 = "NO";
    defparam add_1042_15.INJECT1_1 = "NO";
    CCU2D add_1042_13 (.A0(d7[11]), .B0(d_d7[11]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[12]), .B1(d_d7[12]), .C1(GND_net), .D1(GND_net), .CIN(n11025), 
          .COUT(n11026), .S0(d8_71__N_1602[11]), .S1(d8_71__N_1602[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1042_13.INIT0 = 16'h5999;
    defparam add_1042_13.INIT1 = 16'h5999;
    defparam add_1042_13.INJECT1_0 = "NO";
    defparam add_1042_13.INJECT1_1 = "NO";
    CCU2D add_1042_11 (.A0(d7[9]), .B0(d_d7[9]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[10]), .B1(d_d7[10]), .C1(GND_net), .D1(GND_net), .CIN(n11024), 
          .COUT(n11025), .S0(d8_71__N_1602[9]), .S1(d8_71__N_1602[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1042_11.INIT0 = 16'h5999;
    defparam add_1042_11.INIT1 = 16'h5999;
    defparam add_1042_11.INJECT1_0 = "NO";
    defparam add_1042_11.INJECT1_1 = "NO";
    CCU2D add_1042_9 (.A0(d7[7]), .B0(d_d7[7]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[8]), .B1(d_d7[8]), .C1(GND_net), .D1(GND_net), .CIN(n11023), 
          .COUT(n11024), .S0(d8_71__N_1602[7]), .S1(d8_71__N_1602[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1042_9.INIT0 = 16'h5999;
    defparam add_1042_9.INIT1 = 16'h5999;
    defparam add_1042_9.INJECT1_0 = "NO";
    defparam add_1042_9.INJECT1_1 = "NO";
    CCU2D add_1042_7 (.A0(d7[5]), .B0(d_d7[5]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[6]), .B1(d_d7[6]), .C1(GND_net), .D1(GND_net), .CIN(n11022), 
          .COUT(n11023), .S0(d8_71__N_1602[5]), .S1(d8_71__N_1602[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1042_7.INIT0 = 16'h5999;
    defparam add_1042_7.INIT1 = 16'h5999;
    defparam add_1042_7.INJECT1_0 = "NO";
    defparam add_1042_7.INJECT1_1 = "NO";
    CCU2D add_1042_5 (.A0(d7[3]), .B0(d_d7[3]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[4]), .B1(d_d7[4]), .C1(GND_net), .D1(GND_net), .CIN(n11021), 
          .COUT(n11022), .S0(d8_71__N_1602[3]), .S1(d8_71__N_1602[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1042_5.INIT0 = 16'h5999;
    defparam add_1042_5.INIT1 = 16'h5999;
    defparam add_1042_5.INJECT1_0 = "NO";
    defparam add_1042_5.INJECT1_1 = "NO";
    CCU2D add_1042_3 (.A0(d7[1]), .B0(d_d7[1]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[2]), .B1(d_d7[2]), .C1(GND_net), .D1(GND_net), .CIN(n11020), 
          .COUT(n11021), .S0(d8_71__N_1602[1]), .S1(d8_71__N_1602[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1042_3.INIT0 = 16'h5999;
    defparam add_1042_3.INIT1 = 16'h5999;
    defparam add_1042_3.INJECT1_0 = "NO";
    defparam add_1042_3.INJECT1_1 = "NO";
    CCU2D add_1042_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d7[0]), .B1(d_d7[0]), .C1(GND_net), .D1(GND_net), .COUT(n11020), 
          .S1(d8_71__N_1602[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1042_1.INIT0 = 16'h0000;
    defparam add_1042_1.INIT1 = 16'h5999;
    defparam add_1042_1.INJECT1_0 = "NO";
    defparam add_1042_1.INJECT1_1 = "NO";
    CCU2D add_10_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10988), 
          .S0(n375[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_17.INIT0 = 16'h5aaa;
    defparam add_10_17.INIT1 = 16'h0000;
    defparam add_10_17.INJECT1_0 = "NO";
    defparam add_10_17.INJECT1_1 = "NO";
    CCU2D add_10_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n10987), .COUT(n10988), .S0(n375[13]), .S1(n375[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_15.INIT0 = 16'h5aaa;
    defparam add_10_15.INIT1 = 16'h5aaa;
    defparam add_10_15.INJECT1_0 = "NO";
    defparam add_10_15.INJECT1_1 = "NO";
    CCU2D add_10_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n10986), .COUT(n10987), .S0(n375[11]), .S1(n375[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_13.INIT0 = 16'h5aaa;
    defparam add_10_13.INIT1 = 16'h5aaa;
    defparam add_10_13.INJECT1_0 = "NO";
    defparam add_10_13.INJECT1_1 = "NO";
    CCU2D add_10_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n10985), .COUT(n10986), .S0(n375[9]), .S1(n375[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_11.INIT0 = 16'h5aaa;
    defparam add_10_11.INIT1 = 16'h5aaa;
    defparam add_10_11.INJECT1_0 = "NO";
    defparam add_10_11.INJECT1_1 = "NO";
    CCU2D add_10_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10984), 
          .COUT(n10985), .S0(n375[7]), .S1(n375[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_9.INIT0 = 16'h5aaa;
    defparam add_10_9.INIT1 = 16'h5aaa;
    defparam add_10_9.INJECT1_0 = "NO";
    defparam add_10_9.INJECT1_1 = "NO";
    CCU2D add_10_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10983), 
          .COUT(n10984), .S0(n375[5]), .S1(n375[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_7.INIT0 = 16'h5aaa;
    defparam add_10_7.INIT1 = 16'h5aaa;
    defparam add_10_7.INJECT1_0 = "NO";
    defparam add_10_7.INJECT1_1 = "NO";
    CCU2D add_10_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10982), 
          .COUT(n10983), .S0(n375[3]), .S1(n375[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_5.INIT0 = 16'h5aaa;
    defparam add_10_5.INIT1 = 16'h5aaa;
    defparam add_10_5.INJECT1_0 = "NO";
    defparam add_10_5.INJECT1_1 = "NO";
    CCU2D add_10_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10981), 
          .COUT(n10982), .S0(n375[1]), .S1(n375[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_3.INIT0 = 16'h5aaa;
    defparam add_10_3.INIT1 = 16'h5aaa;
    defparam add_10_3.INJECT1_0 = "NO";
    defparam add_10_3.INJECT1_1 = "NO";
    CCU2D add_10_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n10981), 
          .S1(n375[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(87[24:37])
    defparam add_10_1.INIT0 = 16'hF000;
    defparam add_10_1.INIT1 = 16'h5555;
    defparam add_10_1.INJECT1_0 = "NO";
    defparam add_10_1.INJECT1_1 = "NO";
    CCU2D add_1027_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10962), 
          .S0(n5406));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1027_cout.INIT0 = 16'h0000;
    defparam add_1027_cout.INIT1 = 16'h0000;
    defparam add_1027_cout.INJECT1_0 = "NO";
    defparam add_1027_cout.INJECT1_1 = "NO";
    CCU2D add_1027_36 (.A0(d4[34]), .B0(d5[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[35]), .B1(d5[35]), .C1(GND_net), .D1(GND_net), .CIN(n10961), 
          .COUT(n10962), .S0(d5_71__N_705[34]), .S1(d5_71__N_705[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1027_36.INIT0 = 16'h5666;
    defparam add_1027_36.INIT1 = 16'h5666;
    defparam add_1027_36.INJECT1_0 = "NO";
    defparam add_1027_36.INJECT1_1 = "NO";
    CCU2D add_1027_34 (.A0(d4[32]), .B0(d5[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[33]), .B1(d5[33]), .C1(GND_net), .D1(GND_net), .CIN(n10960), 
          .COUT(n10961), .S0(d5_71__N_705[32]), .S1(d5_71__N_705[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1027_34.INIT0 = 16'h5666;
    defparam add_1027_34.INIT1 = 16'h5666;
    defparam add_1027_34.INJECT1_0 = "NO";
    defparam add_1027_34.INJECT1_1 = "NO";
    CCU2D add_1027_32 (.A0(d4[30]), .B0(d5[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[31]), .B1(d5[31]), .C1(GND_net), .D1(GND_net), .CIN(n10959), 
          .COUT(n10960), .S0(d5_71__N_705[30]), .S1(d5_71__N_705[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1027_32.INIT0 = 16'h5666;
    defparam add_1027_32.INIT1 = 16'h5666;
    defparam add_1027_32.INJECT1_0 = "NO";
    defparam add_1027_32.INJECT1_1 = "NO";
    CCU2D add_1027_30 (.A0(d4[28]), .B0(d5[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[29]), .B1(d5[29]), .C1(GND_net), .D1(GND_net), .CIN(n10958), 
          .COUT(n10959), .S0(d5_71__N_705[28]), .S1(d5_71__N_705[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1027_30.INIT0 = 16'h5666;
    defparam add_1027_30.INIT1 = 16'h5666;
    defparam add_1027_30.INJECT1_0 = "NO";
    defparam add_1027_30.INJECT1_1 = "NO";
    CCU2D add_1027_28 (.A0(d4[26]), .B0(d5[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[27]), .B1(d5[27]), .C1(GND_net), .D1(GND_net), .CIN(n10957), 
          .COUT(n10958), .S0(d5_71__N_705[26]), .S1(d5_71__N_705[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1027_28.INIT0 = 16'h5666;
    defparam add_1027_28.INIT1 = 16'h5666;
    defparam add_1027_28.INJECT1_0 = "NO";
    defparam add_1027_28.INJECT1_1 = "NO";
    CCU2D add_1027_26 (.A0(d4[24]), .B0(d5[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[25]), .B1(d5[25]), .C1(GND_net), .D1(GND_net), .CIN(n10956), 
          .COUT(n10957), .S0(d5_71__N_705[24]), .S1(d5_71__N_705[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1027_26.INIT0 = 16'h5666;
    defparam add_1027_26.INIT1 = 16'h5666;
    defparam add_1027_26.INJECT1_0 = "NO";
    defparam add_1027_26.INJECT1_1 = "NO";
    CCU2D add_1027_24 (.A0(d4[22]), .B0(d5[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[23]), .B1(d5[23]), .C1(GND_net), .D1(GND_net), .CIN(n10955), 
          .COUT(n10956), .S0(d5_71__N_705[22]), .S1(d5_71__N_705[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1027_24.INIT0 = 16'h5666;
    defparam add_1027_24.INIT1 = 16'h5666;
    defparam add_1027_24.INJECT1_0 = "NO";
    defparam add_1027_24.INJECT1_1 = "NO";
    CCU2D add_1027_22 (.A0(d4[20]), .B0(d5[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[21]), .B1(d5[21]), .C1(GND_net), .D1(GND_net), .CIN(n10954), 
          .COUT(n10955), .S0(d5_71__N_705[20]), .S1(d5_71__N_705[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1027_22.INIT0 = 16'h5666;
    defparam add_1027_22.INIT1 = 16'h5666;
    defparam add_1027_22.INJECT1_0 = "NO";
    defparam add_1027_22.INJECT1_1 = "NO";
    CCU2D add_1027_20 (.A0(d4[18]), .B0(d5[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[19]), .B1(d5[19]), .C1(GND_net), .D1(GND_net), .CIN(n10953), 
          .COUT(n10954), .S0(d5_71__N_705[18]), .S1(d5_71__N_705[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1027_20.INIT0 = 16'h5666;
    defparam add_1027_20.INIT1 = 16'h5666;
    defparam add_1027_20.INJECT1_0 = "NO";
    defparam add_1027_20.INJECT1_1 = "NO";
    CCU2D add_1027_18 (.A0(d4[16]), .B0(d5[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[17]), .B1(d5[17]), .C1(GND_net), .D1(GND_net), .CIN(n10952), 
          .COUT(n10953), .S0(d5_71__N_705[16]), .S1(d5_71__N_705[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1027_18.INIT0 = 16'h5666;
    defparam add_1027_18.INIT1 = 16'h5666;
    defparam add_1027_18.INJECT1_0 = "NO";
    defparam add_1027_18.INJECT1_1 = "NO";
    CCU2D add_1027_16 (.A0(d4[14]), .B0(d5[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[15]), .B1(d5[15]), .C1(GND_net), .D1(GND_net), .CIN(n10951), 
          .COUT(n10952), .S0(d5_71__N_705[14]), .S1(d5_71__N_705[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1027_16.INIT0 = 16'h5666;
    defparam add_1027_16.INIT1 = 16'h5666;
    defparam add_1027_16.INJECT1_0 = "NO";
    defparam add_1027_16.INJECT1_1 = "NO";
    CCU2D add_1027_14 (.A0(d4[12]), .B0(d5[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[13]), .B1(d5[13]), .C1(GND_net), .D1(GND_net), .CIN(n10950), 
          .COUT(n10951), .S0(d5_71__N_705[12]), .S1(d5_71__N_705[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1027_14.INIT0 = 16'h5666;
    defparam add_1027_14.INIT1 = 16'h5666;
    defparam add_1027_14.INJECT1_0 = "NO";
    defparam add_1027_14.INJECT1_1 = "NO";
    CCU2D add_1027_12 (.A0(d4[10]), .B0(d5[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[11]), .B1(d5[11]), .C1(GND_net), .D1(GND_net), .CIN(n10949), 
          .COUT(n10950), .S0(d5_71__N_705[10]), .S1(d5_71__N_705[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1027_12.INIT0 = 16'h5666;
    defparam add_1027_12.INIT1 = 16'h5666;
    defparam add_1027_12.INJECT1_0 = "NO";
    defparam add_1027_12.INJECT1_1 = "NO";
    CCU2D add_1027_10 (.A0(d4[8]), .B0(d5[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[9]), .B1(d5[9]), .C1(GND_net), .D1(GND_net), .CIN(n10948), 
          .COUT(n10949), .S0(d5_71__N_705[8]), .S1(d5_71__N_705[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1027_10.INIT0 = 16'h5666;
    defparam add_1027_10.INIT1 = 16'h5666;
    defparam add_1027_10.INJECT1_0 = "NO";
    defparam add_1027_10.INJECT1_1 = "NO";
    CCU2D add_1027_8 (.A0(d4[6]), .B0(d5[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[7]), .B1(d5[7]), .C1(GND_net), .D1(GND_net), .CIN(n10947), 
          .COUT(n10948), .S0(d5_71__N_705[6]), .S1(d5_71__N_705[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1027_8.INIT0 = 16'h5666;
    defparam add_1027_8.INIT1 = 16'h5666;
    defparam add_1027_8.INJECT1_0 = "NO";
    defparam add_1027_8.INJECT1_1 = "NO";
    CCU2D add_1027_6 (.A0(d4[4]), .B0(d5[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[5]), .B1(d5[5]), .C1(GND_net), .D1(GND_net), .CIN(n10946), 
          .COUT(n10947), .S0(d5_71__N_705[4]), .S1(d5_71__N_705[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1027_6.INIT0 = 16'h5666;
    defparam add_1027_6.INIT1 = 16'h5666;
    defparam add_1027_6.INJECT1_0 = "NO";
    defparam add_1027_6.INJECT1_1 = "NO";
    CCU2D add_1027_4 (.A0(d4[2]), .B0(d5[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[3]), .B1(d5[3]), .C1(GND_net), .D1(GND_net), .CIN(n10945), 
          .COUT(n10946), .S0(d5_71__N_705[2]), .S1(d5_71__N_705[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1027_4.INIT0 = 16'h5666;
    defparam add_1027_4.INIT1 = 16'h5666;
    defparam add_1027_4.INJECT1_0 = "NO";
    defparam add_1027_4.INJECT1_1 = "NO";
    CCU2D add_1027_2 (.A0(d4[0]), .B0(d5[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d4[1]), .B1(d5[1]), .C1(GND_net), .D1(GND_net), .COUT(n10945), 
          .S1(d5_71__N_705[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(70[13:20])
    defparam add_1027_2.INIT0 = 16'h7000;
    defparam add_1027_2.INIT1 = 16'h5666;
    defparam add_1027_2.INJECT1_0 = "NO";
    defparam add_1027_2.INJECT1_1 = "NO";
    CCU2D add_1022_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10943), 
          .S0(n5254));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1022_cout.INIT0 = 16'h0000;
    defparam add_1022_cout.INIT1 = 16'h0000;
    defparam add_1022_cout.INJECT1_0 = "NO";
    defparam add_1022_cout.INJECT1_1 = "NO";
    CCU2D add_1022_36 (.A0(d3[34]), .B0(d4[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[35]), .B1(d4[35]), .C1(GND_net), .D1(GND_net), .CIN(n10942), 
          .COUT(n10943), .S0(d4_71__N_633[34]), .S1(d4_71__N_633[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1022_36.INIT0 = 16'h5666;
    defparam add_1022_36.INIT1 = 16'h5666;
    defparam add_1022_36.INJECT1_0 = "NO";
    defparam add_1022_36.INJECT1_1 = "NO";
    CCU2D add_1022_34 (.A0(d3[32]), .B0(d4[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[33]), .B1(d4[33]), .C1(GND_net), .D1(GND_net), .CIN(n10941), 
          .COUT(n10942), .S0(d4_71__N_633[32]), .S1(d4_71__N_633[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1022_34.INIT0 = 16'h5666;
    defparam add_1022_34.INIT1 = 16'h5666;
    defparam add_1022_34.INJECT1_0 = "NO";
    defparam add_1022_34.INJECT1_1 = "NO";
    CCU2D add_1022_32 (.A0(d3[30]), .B0(d4[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[31]), .B1(d4[31]), .C1(GND_net), .D1(GND_net), .CIN(n10940), 
          .COUT(n10941), .S0(d4_71__N_633[30]), .S1(d4_71__N_633[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1022_32.INIT0 = 16'h5666;
    defparam add_1022_32.INIT1 = 16'h5666;
    defparam add_1022_32.INJECT1_0 = "NO";
    defparam add_1022_32.INJECT1_1 = "NO";
    CCU2D add_1022_30 (.A0(d3[28]), .B0(d4[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[29]), .B1(d4[29]), .C1(GND_net), .D1(GND_net), .CIN(n10939), 
          .COUT(n10940), .S0(d4_71__N_633[28]), .S1(d4_71__N_633[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1022_30.INIT0 = 16'h5666;
    defparam add_1022_30.INIT1 = 16'h5666;
    defparam add_1022_30.INJECT1_0 = "NO";
    defparam add_1022_30.INJECT1_1 = "NO";
    CCU2D add_1022_28 (.A0(d3[26]), .B0(d4[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[27]), .B1(d4[27]), .C1(GND_net), .D1(GND_net), .CIN(n10938), 
          .COUT(n10939), .S0(d4_71__N_633[26]), .S1(d4_71__N_633[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1022_28.INIT0 = 16'h5666;
    defparam add_1022_28.INIT1 = 16'h5666;
    defparam add_1022_28.INJECT1_0 = "NO";
    defparam add_1022_28.INJECT1_1 = "NO";
    CCU2D add_1022_26 (.A0(d3[24]), .B0(d4[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[25]), .B1(d4[25]), .C1(GND_net), .D1(GND_net), .CIN(n10937), 
          .COUT(n10938), .S0(d4_71__N_633[24]), .S1(d4_71__N_633[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1022_26.INIT0 = 16'h5666;
    defparam add_1022_26.INIT1 = 16'h5666;
    defparam add_1022_26.INJECT1_0 = "NO";
    defparam add_1022_26.INJECT1_1 = "NO";
    CCU2D add_1022_24 (.A0(d3[22]), .B0(d4[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[23]), .B1(d4[23]), .C1(GND_net), .D1(GND_net), .CIN(n10936), 
          .COUT(n10937), .S0(d4_71__N_633[22]), .S1(d4_71__N_633[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1022_24.INIT0 = 16'h5666;
    defparam add_1022_24.INIT1 = 16'h5666;
    defparam add_1022_24.INJECT1_0 = "NO";
    defparam add_1022_24.INJECT1_1 = "NO";
    CCU2D add_1022_22 (.A0(d3[20]), .B0(d4[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[21]), .B1(d4[21]), .C1(GND_net), .D1(GND_net), .CIN(n10935), 
          .COUT(n10936), .S0(d4_71__N_633[20]), .S1(d4_71__N_633[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1022_22.INIT0 = 16'h5666;
    defparam add_1022_22.INIT1 = 16'h5666;
    defparam add_1022_22.INJECT1_0 = "NO";
    defparam add_1022_22.INJECT1_1 = "NO";
    CCU2D add_1022_20 (.A0(d3[18]), .B0(d4[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[19]), .B1(d4[19]), .C1(GND_net), .D1(GND_net), .CIN(n10934), 
          .COUT(n10935), .S0(d4_71__N_633[18]), .S1(d4_71__N_633[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1022_20.INIT0 = 16'h5666;
    defparam add_1022_20.INIT1 = 16'h5666;
    defparam add_1022_20.INJECT1_0 = "NO";
    defparam add_1022_20.INJECT1_1 = "NO";
    CCU2D add_1022_18 (.A0(d3[16]), .B0(d4[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[17]), .B1(d4[17]), .C1(GND_net), .D1(GND_net), .CIN(n10933), 
          .COUT(n10934), .S0(d4_71__N_633[16]), .S1(d4_71__N_633[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1022_18.INIT0 = 16'h5666;
    defparam add_1022_18.INIT1 = 16'h5666;
    defparam add_1022_18.INJECT1_0 = "NO";
    defparam add_1022_18.INJECT1_1 = "NO";
    CCU2D add_1022_16 (.A0(d3[14]), .B0(d4[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[15]), .B1(d4[15]), .C1(GND_net), .D1(GND_net), .CIN(n10932), 
          .COUT(n10933), .S0(d4_71__N_633[14]), .S1(d4_71__N_633[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1022_16.INIT0 = 16'h5666;
    defparam add_1022_16.INIT1 = 16'h5666;
    defparam add_1022_16.INJECT1_0 = "NO";
    defparam add_1022_16.INJECT1_1 = "NO";
    CCU2D add_1022_14 (.A0(d3[12]), .B0(d4[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[13]), .B1(d4[13]), .C1(GND_net), .D1(GND_net), .CIN(n10931), 
          .COUT(n10932), .S0(d4_71__N_633[12]), .S1(d4_71__N_633[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1022_14.INIT0 = 16'h5666;
    defparam add_1022_14.INIT1 = 16'h5666;
    defparam add_1022_14.INJECT1_0 = "NO";
    defparam add_1022_14.INJECT1_1 = "NO";
    CCU2D add_1022_12 (.A0(d3[10]), .B0(d4[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[11]), .B1(d4[11]), .C1(GND_net), .D1(GND_net), .CIN(n10930), 
          .COUT(n10931), .S0(d4_71__N_633[10]), .S1(d4_71__N_633[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1022_12.INIT0 = 16'h5666;
    defparam add_1022_12.INIT1 = 16'h5666;
    defparam add_1022_12.INJECT1_0 = "NO";
    defparam add_1022_12.INJECT1_1 = "NO";
    CCU2D add_1022_10 (.A0(d3[8]), .B0(d4[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[9]), .B1(d4[9]), .C1(GND_net), .D1(GND_net), .CIN(n10929), 
          .COUT(n10930), .S0(d4_71__N_633[8]), .S1(d4_71__N_633[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1022_10.INIT0 = 16'h5666;
    defparam add_1022_10.INIT1 = 16'h5666;
    defparam add_1022_10.INJECT1_0 = "NO";
    defparam add_1022_10.INJECT1_1 = "NO";
    CCU2D add_1022_8 (.A0(d3[6]), .B0(d4[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[7]), .B1(d4[7]), .C1(GND_net), .D1(GND_net), .CIN(n10928), 
          .COUT(n10929), .S0(d4_71__N_633[6]), .S1(d4_71__N_633[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1022_8.INIT0 = 16'h5666;
    defparam add_1022_8.INIT1 = 16'h5666;
    defparam add_1022_8.INJECT1_0 = "NO";
    defparam add_1022_8.INJECT1_1 = "NO";
    CCU2D add_1022_6 (.A0(d3[4]), .B0(d4[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[5]), .B1(d4[5]), .C1(GND_net), .D1(GND_net), .CIN(n10927), 
          .COUT(n10928), .S0(d4_71__N_633[4]), .S1(d4_71__N_633[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1022_6.INIT0 = 16'h5666;
    defparam add_1022_6.INIT1 = 16'h5666;
    defparam add_1022_6.INJECT1_0 = "NO";
    defparam add_1022_6.INJECT1_1 = "NO";
    CCU2D add_1022_4 (.A0(d3[2]), .B0(d4[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[3]), .B1(d4[3]), .C1(GND_net), .D1(GND_net), .CIN(n10926), 
          .COUT(n10927), .S0(d4_71__N_633[2]), .S1(d4_71__N_633[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1022_4.INIT0 = 16'h5666;
    defparam add_1022_4.INIT1 = 16'h5666;
    defparam add_1022_4.INJECT1_0 = "NO";
    defparam add_1022_4.INJECT1_1 = "NO";
    CCU2D add_1022_2 (.A0(d3[0]), .B0(d4[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d3[1]), .B1(d4[1]), .C1(GND_net), .D1(GND_net), .COUT(n10926), 
          .S1(d4_71__N_633[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(68[13:20])
    defparam add_1022_2.INIT0 = 16'h7000;
    defparam add_1022_2.INIT1 = 16'h5666;
    defparam add_1022_2.INJECT1_0 = "NO";
    defparam add_1022_2.INJECT1_1 = "NO";
    CCU2D add_1017_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10924), 
          .S0(n5102));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1017_cout.INIT0 = 16'h0000;
    defparam add_1017_cout.INIT1 = 16'h0000;
    defparam add_1017_cout.INJECT1_0 = "NO";
    defparam add_1017_cout.INJECT1_1 = "NO";
    CCU2D add_1017_36 (.A0(d2[34]), .B0(d3[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[35]), .B1(d3[35]), .C1(GND_net), .D1(GND_net), .CIN(n10923), 
          .COUT(n10924), .S0(d3_71__N_561[34]), .S1(d3_71__N_561[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1017_36.INIT0 = 16'h5666;
    defparam add_1017_36.INIT1 = 16'h5666;
    defparam add_1017_36.INJECT1_0 = "NO";
    defparam add_1017_36.INJECT1_1 = "NO";
    CCU2D add_1017_34 (.A0(d2[32]), .B0(d3[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[33]), .B1(d3[33]), .C1(GND_net), .D1(GND_net), .CIN(n10922), 
          .COUT(n10923), .S0(d3_71__N_561[32]), .S1(d3_71__N_561[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1017_34.INIT0 = 16'h5666;
    defparam add_1017_34.INIT1 = 16'h5666;
    defparam add_1017_34.INJECT1_0 = "NO";
    defparam add_1017_34.INJECT1_1 = "NO";
    CCU2D add_1017_32 (.A0(d2[30]), .B0(d3[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[31]), .B1(d3[31]), .C1(GND_net), .D1(GND_net), .CIN(n10921), 
          .COUT(n10922), .S0(d3_71__N_561[30]), .S1(d3_71__N_561[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1017_32.INIT0 = 16'h5666;
    defparam add_1017_32.INIT1 = 16'h5666;
    defparam add_1017_32.INJECT1_0 = "NO";
    defparam add_1017_32.INJECT1_1 = "NO";
    CCU2D add_1017_30 (.A0(d2[28]), .B0(d3[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[29]), .B1(d3[29]), .C1(GND_net), .D1(GND_net), .CIN(n10920), 
          .COUT(n10921), .S0(d3_71__N_561[28]), .S1(d3_71__N_561[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1017_30.INIT0 = 16'h5666;
    defparam add_1017_30.INIT1 = 16'h5666;
    defparam add_1017_30.INJECT1_0 = "NO";
    defparam add_1017_30.INJECT1_1 = "NO";
    CCU2D add_1017_28 (.A0(d2[26]), .B0(d3[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[27]), .B1(d3[27]), .C1(GND_net), .D1(GND_net), .CIN(n10919), 
          .COUT(n10920), .S0(d3_71__N_561[26]), .S1(d3_71__N_561[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1017_28.INIT0 = 16'h5666;
    defparam add_1017_28.INIT1 = 16'h5666;
    defparam add_1017_28.INJECT1_0 = "NO";
    defparam add_1017_28.INJECT1_1 = "NO";
    CCU2D add_1017_26 (.A0(d2[24]), .B0(d3[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[25]), .B1(d3[25]), .C1(GND_net), .D1(GND_net), .CIN(n10918), 
          .COUT(n10919), .S0(d3_71__N_561[24]), .S1(d3_71__N_561[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1017_26.INIT0 = 16'h5666;
    defparam add_1017_26.INIT1 = 16'h5666;
    defparam add_1017_26.INJECT1_0 = "NO";
    defparam add_1017_26.INJECT1_1 = "NO";
    CCU2D add_1017_24 (.A0(d2[22]), .B0(d3[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[23]), .B1(d3[23]), .C1(GND_net), .D1(GND_net), .CIN(n10917), 
          .COUT(n10918), .S0(d3_71__N_561[22]), .S1(d3_71__N_561[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1017_24.INIT0 = 16'h5666;
    defparam add_1017_24.INIT1 = 16'h5666;
    defparam add_1017_24.INJECT1_0 = "NO";
    defparam add_1017_24.INJECT1_1 = "NO";
    CCU2D add_1017_22 (.A0(d2[20]), .B0(d3[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[21]), .B1(d3[21]), .C1(GND_net), .D1(GND_net), .CIN(n10916), 
          .COUT(n10917), .S0(d3_71__N_561[20]), .S1(d3_71__N_561[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1017_22.INIT0 = 16'h5666;
    defparam add_1017_22.INIT1 = 16'h5666;
    defparam add_1017_22.INJECT1_0 = "NO";
    defparam add_1017_22.INJECT1_1 = "NO";
    CCU2D add_1017_20 (.A0(d2[18]), .B0(d3[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[19]), .B1(d3[19]), .C1(GND_net), .D1(GND_net), .CIN(n10915), 
          .COUT(n10916), .S0(d3_71__N_561[18]), .S1(d3_71__N_561[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1017_20.INIT0 = 16'h5666;
    defparam add_1017_20.INIT1 = 16'h5666;
    defparam add_1017_20.INJECT1_0 = "NO";
    defparam add_1017_20.INJECT1_1 = "NO";
    CCU2D add_1017_18 (.A0(d2[16]), .B0(d3[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[17]), .B1(d3[17]), .C1(GND_net), .D1(GND_net), .CIN(n10914), 
          .COUT(n10915), .S0(d3_71__N_561[16]), .S1(d3_71__N_561[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1017_18.INIT0 = 16'h5666;
    defparam add_1017_18.INIT1 = 16'h5666;
    defparam add_1017_18.INJECT1_0 = "NO";
    defparam add_1017_18.INJECT1_1 = "NO";
    CCU2D add_1017_16 (.A0(d2[14]), .B0(d3[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[15]), .B1(d3[15]), .C1(GND_net), .D1(GND_net), .CIN(n10913), 
          .COUT(n10914), .S0(d3_71__N_561[14]), .S1(d3_71__N_561[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1017_16.INIT0 = 16'h5666;
    defparam add_1017_16.INIT1 = 16'h5666;
    defparam add_1017_16.INJECT1_0 = "NO";
    defparam add_1017_16.INJECT1_1 = "NO";
    CCU2D add_1017_14 (.A0(d2[12]), .B0(d3[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[13]), .B1(d3[13]), .C1(GND_net), .D1(GND_net), .CIN(n10912), 
          .COUT(n10913), .S0(d3_71__N_561[12]), .S1(d3_71__N_561[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1017_14.INIT0 = 16'h5666;
    defparam add_1017_14.INIT1 = 16'h5666;
    defparam add_1017_14.INJECT1_0 = "NO";
    defparam add_1017_14.INJECT1_1 = "NO";
    CCU2D add_1017_12 (.A0(d2[10]), .B0(d3[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[11]), .B1(d3[11]), .C1(GND_net), .D1(GND_net), .CIN(n10911), 
          .COUT(n10912), .S0(d3_71__N_561[10]), .S1(d3_71__N_561[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1017_12.INIT0 = 16'h5666;
    defparam add_1017_12.INIT1 = 16'h5666;
    defparam add_1017_12.INJECT1_0 = "NO";
    defparam add_1017_12.INJECT1_1 = "NO";
    CCU2D add_1017_10 (.A0(d2[8]), .B0(d3[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[9]), .B1(d3[9]), .C1(GND_net), .D1(GND_net), .CIN(n10910), 
          .COUT(n10911), .S0(d3_71__N_561[8]), .S1(d3_71__N_561[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1017_10.INIT0 = 16'h5666;
    defparam add_1017_10.INIT1 = 16'h5666;
    defparam add_1017_10.INJECT1_0 = "NO";
    defparam add_1017_10.INJECT1_1 = "NO";
    CCU2D add_1017_8 (.A0(d2[6]), .B0(d3[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[7]), .B1(d3[7]), .C1(GND_net), .D1(GND_net), .CIN(n10909), 
          .COUT(n10910), .S0(d3_71__N_561[6]), .S1(d3_71__N_561[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1017_8.INIT0 = 16'h5666;
    defparam add_1017_8.INIT1 = 16'h5666;
    defparam add_1017_8.INJECT1_0 = "NO";
    defparam add_1017_8.INJECT1_1 = "NO";
    CCU2D add_1017_6 (.A0(d2[4]), .B0(d3[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[5]), .B1(d3[5]), .C1(GND_net), .D1(GND_net), .CIN(n10908), 
          .COUT(n10909), .S0(d3_71__N_561[4]), .S1(d3_71__N_561[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1017_6.INIT0 = 16'h5666;
    defparam add_1017_6.INIT1 = 16'h5666;
    defparam add_1017_6.INJECT1_0 = "NO";
    defparam add_1017_6.INJECT1_1 = "NO";
    CCU2D add_1017_4 (.A0(d2[2]), .B0(d3[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[3]), .B1(d3[3]), .C1(GND_net), .D1(GND_net), .CIN(n10907), 
          .COUT(n10908), .S0(d3_71__N_561[2]), .S1(d3_71__N_561[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1017_4.INIT0 = 16'h5666;
    defparam add_1017_4.INIT1 = 16'h5666;
    defparam add_1017_4.INJECT1_0 = "NO";
    defparam add_1017_4.INJECT1_1 = "NO";
    CCU2D add_1017_2 (.A0(d2[0]), .B0(d3[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[1]), .B1(d3[1]), .C1(GND_net), .D1(GND_net), .COUT(n10907), 
          .S1(d3_71__N_561[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1017_2.INIT0 = 16'h7000;
    defparam add_1017_2.INIT1 = 16'h5666;
    defparam add_1017_2.INJECT1_0 = "NO";
    defparam add_1017_2.INJECT1_1 = "NO";
    CCU2D add_1012_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10905), 
          .S0(n4950));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1012_cout.INIT0 = 16'h0000;
    defparam add_1012_cout.INIT1 = 16'h0000;
    defparam add_1012_cout.INJECT1_0 = "NO";
    defparam add_1012_cout.INJECT1_1 = "NO";
    CCU2D add_1012_36 (.A0(d1[34]), .B0(d2[34]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[35]), .B1(d2[35]), .C1(GND_net), .D1(GND_net), .CIN(n10904), 
          .COUT(n10905), .S0(d2_71__N_489[34]), .S1(d2_71__N_489[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1012_36.INIT0 = 16'h5666;
    defparam add_1012_36.INIT1 = 16'h5666;
    defparam add_1012_36.INJECT1_0 = "NO";
    defparam add_1012_36.INJECT1_1 = "NO";
    CCU2D add_1012_34 (.A0(d1[32]), .B0(d2[32]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[33]), .B1(d2[33]), .C1(GND_net), .D1(GND_net), .CIN(n10903), 
          .COUT(n10904), .S0(d2_71__N_489[32]), .S1(d2_71__N_489[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1012_34.INIT0 = 16'h5666;
    defparam add_1012_34.INIT1 = 16'h5666;
    defparam add_1012_34.INJECT1_0 = "NO";
    defparam add_1012_34.INJECT1_1 = "NO";
    CCU2D add_1012_32 (.A0(d1[30]), .B0(d2[30]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[31]), .B1(d2[31]), .C1(GND_net), .D1(GND_net), .CIN(n10902), 
          .COUT(n10903), .S0(d2_71__N_489[30]), .S1(d2_71__N_489[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1012_32.INIT0 = 16'h5666;
    defparam add_1012_32.INIT1 = 16'h5666;
    defparam add_1012_32.INJECT1_0 = "NO";
    defparam add_1012_32.INJECT1_1 = "NO";
    CCU2D add_1012_30 (.A0(d1[28]), .B0(d2[28]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[29]), .B1(d2[29]), .C1(GND_net), .D1(GND_net), .CIN(n10901), 
          .COUT(n10902), .S0(d2_71__N_489[28]), .S1(d2_71__N_489[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1012_30.INIT0 = 16'h5666;
    defparam add_1012_30.INIT1 = 16'h5666;
    defparam add_1012_30.INJECT1_0 = "NO";
    defparam add_1012_30.INJECT1_1 = "NO";
    CCU2D add_1012_28 (.A0(d1[26]), .B0(d2[26]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[27]), .B1(d2[27]), .C1(GND_net), .D1(GND_net), .CIN(n10900), 
          .COUT(n10901), .S0(d2_71__N_489[26]), .S1(d2_71__N_489[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1012_28.INIT0 = 16'h5666;
    defparam add_1012_28.INIT1 = 16'h5666;
    defparam add_1012_28.INJECT1_0 = "NO";
    defparam add_1012_28.INJECT1_1 = "NO";
    CCU2D add_1012_26 (.A0(d1[24]), .B0(d2[24]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[25]), .B1(d2[25]), .C1(GND_net), .D1(GND_net), .CIN(n10899), 
          .COUT(n10900), .S0(d2_71__N_489[24]), .S1(d2_71__N_489[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1012_26.INIT0 = 16'h5666;
    defparam add_1012_26.INIT1 = 16'h5666;
    defparam add_1012_26.INJECT1_0 = "NO";
    defparam add_1012_26.INJECT1_1 = "NO";
    CCU2D add_1012_24 (.A0(d1[22]), .B0(d2[22]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[23]), .B1(d2[23]), .C1(GND_net), .D1(GND_net), .CIN(n10898), 
          .COUT(n10899), .S0(d2_71__N_489[22]), .S1(d2_71__N_489[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1012_24.INIT0 = 16'h5666;
    defparam add_1012_24.INIT1 = 16'h5666;
    defparam add_1012_24.INJECT1_0 = "NO";
    defparam add_1012_24.INJECT1_1 = "NO";
    CCU2D add_1012_22 (.A0(d1[20]), .B0(d2[20]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[21]), .B1(d2[21]), .C1(GND_net), .D1(GND_net), .CIN(n10897), 
          .COUT(n10898), .S0(d2_71__N_489[20]), .S1(d2_71__N_489[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1012_22.INIT0 = 16'h5666;
    defparam add_1012_22.INIT1 = 16'h5666;
    defparam add_1012_22.INJECT1_0 = "NO";
    defparam add_1012_22.INJECT1_1 = "NO";
    CCU2D add_1012_20 (.A0(d1[18]), .B0(d2[18]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[19]), .B1(d2[19]), .C1(GND_net), .D1(GND_net), .CIN(n10896), 
          .COUT(n10897), .S0(d2_71__N_489[18]), .S1(d2_71__N_489[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1012_20.INIT0 = 16'h5666;
    defparam add_1012_20.INIT1 = 16'h5666;
    defparam add_1012_20.INJECT1_0 = "NO";
    defparam add_1012_20.INJECT1_1 = "NO";
    CCU2D add_1012_18 (.A0(d1[16]), .B0(d2[16]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[17]), .B1(d2[17]), .C1(GND_net), .D1(GND_net), .CIN(n10895), 
          .COUT(n10896), .S0(d2_71__N_489[16]), .S1(d2_71__N_489[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1012_18.INIT0 = 16'h5666;
    defparam add_1012_18.INIT1 = 16'h5666;
    defparam add_1012_18.INJECT1_0 = "NO";
    defparam add_1012_18.INJECT1_1 = "NO";
    CCU2D add_1012_16 (.A0(d1[14]), .B0(d2[14]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[15]), .B1(d2[15]), .C1(GND_net), .D1(GND_net), .CIN(n10894), 
          .COUT(n10895), .S0(d2_71__N_489[14]), .S1(d2_71__N_489[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1012_16.INIT0 = 16'h5666;
    defparam add_1012_16.INIT1 = 16'h5666;
    defparam add_1012_16.INJECT1_0 = "NO";
    defparam add_1012_16.INJECT1_1 = "NO";
    CCU2D add_1012_14 (.A0(d1[12]), .B0(d2[12]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[13]), .B1(d2[13]), .C1(GND_net), .D1(GND_net), .CIN(n10893), 
          .COUT(n10894), .S0(d2_71__N_489[12]), .S1(d2_71__N_489[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1012_14.INIT0 = 16'h5666;
    defparam add_1012_14.INIT1 = 16'h5666;
    defparam add_1012_14.INJECT1_0 = "NO";
    defparam add_1012_14.INJECT1_1 = "NO";
    CCU2D add_1012_12 (.A0(d1[10]), .B0(d2[10]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[11]), .B1(d2[11]), .C1(GND_net), .D1(GND_net), .CIN(n10892), 
          .COUT(n10893), .S0(d2_71__N_489[10]), .S1(d2_71__N_489[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1012_12.INIT0 = 16'h5666;
    defparam add_1012_12.INIT1 = 16'h5666;
    defparam add_1012_12.INJECT1_0 = "NO";
    defparam add_1012_12.INJECT1_1 = "NO";
    CCU2D add_1012_10 (.A0(d1[8]), .B0(d2[8]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[9]), .B1(d2[9]), .C1(GND_net), .D1(GND_net), .CIN(n10891), 
          .COUT(n10892), .S0(d2_71__N_489[8]), .S1(d2_71__N_489[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1012_10.INIT0 = 16'h5666;
    defparam add_1012_10.INIT1 = 16'h5666;
    defparam add_1012_10.INJECT1_0 = "NO";
    defparam add_1012_10.INJECT1_1 = "NO";
    CCU2D add_1012_8 (.A0(d1[6]), .B0(d2[6]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[7]), .B1(d2[7]), .C1(GND_net), .D1(GND_net), .CIN(n10890), 
          .COUT(n10891), .S0(d2_71__N_489[6]), .S1(d2_71__N_489[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1012_8.INIT0 = 16'h5666;
    defparam add_1012_8.INIT1 = 16'h5666;
    defparam add_1012_8.INJECT1_0 = "NO";
    defparam add_1012_8.INJECT1_1 = "NO";
    CCU2D add_1012_6 (.A0(d1[4]), .B0(d2[4]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[5]), .B1(d2[5]), .C1(GND_net), .D1(GND_net), .CIN(n10889), 
          .COUT(n10890), .S0(d2_71__N_489[4]), .S1(d2_71__N_489[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1012_6.INIT0 = 16'h5666;
    defparam add_1012_6.INIT1 = 16'h5666;
    defparam add_1012_6.INJECT1_0 = "NO";
    defparam add_1012_6.INJECT1_1 = "NO";
    CCU2D add_1012_4 (.A0(d1[2]), .B0(d2[2]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[3]), .B1(d2[3]), .C1(GND_net), .D1(GND_net), .CIN(n10888), 
          .COUT(n10889), .S0(d2_71__N_489[2]), .S1(d2_71__N_489[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1012_4.INIT0 = 16'h5666;
    defparam add_1012_4.INIT1 = 16'h5666;
    defparam add_1012_4.INJECT1_0 = "NO";
    defparam add_1012_4.INJECT1_1 = "NO";
    CCU2D add_1012_2 (.A0(d1[0]), .B0(d2[0]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[1]), .B1(d2[1]), .C1(GND_net), .D1(GND_net), .COUT(n10888), 
          .S1(d2_71__N_489[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1012_2.INIT0 = 16'h7000;
    defparam add_1012_2.INIT1 = 16'h5666;
    defparam add_1012_2.INJECT1_0 = "NO";
    defparam add_1012_2.INJECT1_1 = "NO";
    CCU2D add_1007_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10878), 
          .S0(n4798));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1007_cout.INIT0 = 16'h0000;
    defparam add_1007_cout.INIT1 = 16'h0000;
    defparam add_1007_cout.INJECT1_0 = "NO";
    defparam add_1007_cout.INJECT1_1 = "NO";
    CCU2D add_1007_36 (.A0(MixerOutCos[11]), .B0(d1[34]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[35]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10877), .COUT(n10878), .S0(d1_71__N_417[34]), 
          .S1(d1_71__N_417[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1007_36.INIT0 = 16'h5666;
    defparam add_1007_36.INIT1 = 16'h5666;
    defparam add_1007_36.INJECT1_0 = "NO";
    defparam add_1007_36.INJECT1_1 = "NO";
    CCU2D add_1007_34 (.A0(MixerOutCos[11]), .B0(d1[32]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[33]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10876), .COUT(n10877), .S0(d1_71__N_417[32]), 
          .S1(d1_71__N_417[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1007_34.INIT0 = 16'h5666;
    defparam add_1007_34.INIT1 = 16'h5666;
    defparam add_1007_34.INJECT1_0 = "NO";
    defparam add_1007_34.INJECT1_1 = "NO";
    CCU2D add_1007_32 (.A0(MixerOutCos[11]), .B0(d1[30]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10875), .COUT(n10876), .S0(d1_71__N_417[30]), 
          .S1(d1_71__N_417[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1007_32.INIT0 = 16'h5666;
    defparam add_1007_32.INIT1 = 16'h5666;
    defparam add_1007_32.INJECT1_0 = "NO";
    defparam add_1007_32.INJECT1_1 = "NO";
    CCU2D add_1007_30 (.A0(MixerOutCos[11]), .B0(d1[28]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10874), .COUT(n10875), .S0(d1_71__N_417[28]), 
          .S1(d1_71__N_417[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1007_30.INIT0 = 16'h5666;
    defparam add_1007_30.INIT1 = 16'h5666;
    defparam add_1007_30.INJECT1_0 = "NO";
    defparam add_1007_30.INJECT1_1 = "NO";
    CCU2D add_1007_28 (.A0(MixerOutCos[11]), .B0(d1[26]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10873), .COUT(n10874), .S0(d1_71__N_417[26]), 
          .S1(d1_71__N_417[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1007_28.INIT0 = 16'h5666;
    defparam add_1007_28.INIT1 = 16'h5666;
    defparam add_1007_28.INJECT1_0 = "NO";
    defparam add_1007_28.INJECT1_1 = "NO";
    CCU2D add_1007_26 (.A0(MixerOutCos[11]), .B0(d1[24]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10872), .COUT(n10873), .S0(d1_71__N_417[24]), 
          .S1(d1_71__N_417[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1007_26.INIT0 = 16'h5666;
    defparam add_1007_26.INIT1 = 16'h5666;
    defparam add_1007_26.INJECT1_0 = "NO";
    defparam add_1007_26.INJECT1_1 = "NO";
    CCU2D add_1007_24 (.A0(MixerOutCos[11]), .B0(d1[22]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10871), .COUT(n10872), .S0(d1_71__N_417[22]), 
          .S1(d1_71__N_417[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1007_24.INIT0 = 16'h5666;
    defparam add_1007_24.INIT1 = 16'h5666;
    defparam add_1007_24.INJECT1_0 = "NO";
    defparam add_1007_24.INJECT1_1 = "NO";
    CCU2D add_1007_22 (.A0(MixerOutCos[11]), .B0(d1[20]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10870), .COUT(n10871), .S0(d1_71__N_417[20]), 
          .S1(d1_71__N_417[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1007_22.INIT0 = 16'h5666;
    defparam add_1007_22.INIT1 = 16'h5666;
    defparam add_1007_22.INJECT1_0 = "NO";
    defparam add_1007_22.INJECT1_1 = "NO";
    CCU2D add_1007_20 (.A0(MixerOutCos[11]), .B0(d1[18]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10869), .COUT(n10870), .S0(d1_71__N_417[18]), 
          .S1(d1_71__N_417[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1007_20.INIT0 = 16'h5666;
    defparam add_1007_20.INIT1 = 16'h5666;
    defparam add_1007_20.INJECT1_0 = "NO";
    defparam add_1007_20.INJECT1_1 = "NO";
    CCU2D add_1007_18 (.A0(MixerOutCos[11]), .B0(d1[16]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10868), .COUT(n10869), .S0(d1_71__N_417[16]), 
          .S1(d1_71__N_417[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1007_18.INIT0 = 16'h5666;
    defparam add_1007_18.INIT1 = 16'h5666;
    defparam add_1007_18.INJECT1_0 = "NO";
    defparam add_1007_18.INJECT1_1 = "NO";
    CCU2D add_1007_16 (.A0(MixerOutCos[11]), .B0(d1[14]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10867), .COUT(n10868), .S0(d1_71__N_417[14]), 
          .S1(d1_71__N_417[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1007_16.INIT0 = 16'h5666;
    defparam add_1007_16.INIT1 = 16'h5666;
    defparam add_1007_16.INJECT1_0 = "NO";
    defparam add_1007_16.INJECT1_1 = "NO";
    CCU2D add_1007_14 (.A0(MixerOutCos[11]), .B0(d1[12]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10866), .COUT(n10867), .S0(d1_71__N_417[12]), 
          .S1(d1_71__N_417[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1007_14.INIT0 = 16'h5666;
    defparam add_1007_14.INIT1 = 16'h5666;
    defparam add_1007_14.INJECT1_0 = "NO";
    defparam add_1007_14.INJECT1_1 = "NO";
    CCU2D add_1007_12 (.A0(MixerOutCos[10]), .B0(d1[10]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10865), .COUT(n10866), .S0(d1_71__N_417[10]), 
          .S1(d1_71__N_417[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1007_12.INIT0 = 16'h5666;
    defparam add_1007_12.INIT1 = 16'h5666;
    defparam add_1007_12.INJECT1_0 = "NO";
    defparam add_1007_12.INJECT1_1 = "NO";
    CCU2D add_1007_10 (.A0(MixerOutCos[8]), .B0(d1[8]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[9]), .B1(d1[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10864), .COUT(n10865), .S0(d1_71__N_417[8]), 
          .S1(d1_71__N_417[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1007_10.INIT0 = 16'h5666;
    defparam add_1007_10.INIT1 = 16'h5666;
    defparam add_1007_10.INJECT1_0 = "NO";
    defparam add_1007_10.INJECT1_1 = "NO";
    CCU2D add_1007_8 (.A0(MixerOutCos[6]), .B0(d1[6]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutCos[7]), .B1(d1[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10863), .COUT(n10864), .S0(d1_71__N_417[6]), .S1(d1_71__N_417[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1007_8.INIT0 = 16'h5666;
    defparam add_1007_8.INIT1 = 16'h5666;
    defparam add_1007_8.INJECT1_0 = "NO";
    defparam add_1007_8.INJECT1_1 = "NO";
    CCU2D add_1007_6 (.A0(MixerOutCos[4]), .B0(d1[4]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutCos[5]), .B1(d1[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10862), .COUT(n10863), .S0(d1_71__N_417[4]), .S1(d1_71__N_417[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1007_6.INIT0 = 16'h5666;
    defparam add_1007_6.INIT1 = 16'h5666;
    defparam add_1007_6.INJECT1_0 = "NO";
    defparam add_1007_6.INJECT1_1 = "NO";
    CCU2D add_1007_4 (.A0(MixerOutCos[2]), .B0(d1[2]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutCos[3]), .B1(d1[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10861), .COUT(n10862), .S0(d1_71__N_417[2]), .S1(d1_71__N_417[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1007_4.INIT0 = 16'h5666;
    defparam add_1007_4.INIT1 = 16'h5666;
    defparam add_1007_4.INJECT1_0 = "NO";
    defparam add_1007_4.INJECT1_1 = "NO";
    CCU2D add_1007_2 (.A0(MixerOutCos[0]), .B0(d1[0]), .C0(GND_net), .D0(GND_net), 
          .A1(MixerOutCos[1]), .B1(d1[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n10861), .S1(d1_71__N_417[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1007_2.INIT0 = 16'h7000;
    defparam add_1007_2.INIT1 = 16'h5666;
    defparam add_1007_2.INJECT1_0 = "NO";
    defparam add_1007_2.INJECT1_1 = "NO";
    CCU2D add_1043_3 (.A0(d7[37]), .B0(d_d7[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d7[38]), .B1(d_d7[38]), .C1(GND_net), .D1(GND_net), .CIN(n11649), 
          .COUT(n11650), .S0(n5863[1]), .S1(n5863[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1043_3.INIT0 = 16'h5999;
    defparam add_1043_3.INIT1 = 16'h5999;
    defparam add_1043_3.INJECT1_0 = "NO";
    defparam add_1043_3.INJECT1_1 = "NO";
    CCU2D add_1043_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d7[36]), .B1(d_d7[36]), .C1(GND_net), .D1(GND_net), .COUT(n11649), 
          .S1(n5863[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1043_1.INIT0 = 16'hF000;
    defparam add_1043_1.INIT1 = 16'h5999;
    defparam add_1043_1.INJECT1_0 = "NO";
    defparam add_1043_1.INJECT1_1 = "NO";
    CCU2D add_1044_37 (.A0(d_d7[70]), .B0(n5862), .C0(n5863[34]), .D0(d7[70]), 
          .A1(d_d7[71]), .B1(n5862), .C1(n5863[35]), .D1(d7[71]), .CIN(n11647), 
          .S0(d8_71__N_1602[70]), .S1(d8_71__N_1602[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1044_37.INIT0 = 16'hb874;
    defparam add_1044_37.INIT1 = 16'hb874;
    defparam add_1044_37.INJECT1_0 = "NO";
    defparam add_1044_37.INJECT1_1 = "NO";
    CCU2D add_1044_35 (.A0(d_d7[68]), .B0(n5862), .C0(n5863[32]), .D0(d7[68]), 
          .A1(d_d7[69]), .B1(n5862), .C1(n5863[33]), .D1(d7[69]), .CIN(n11646), 
          .COUT(n11647), .S0(d8_71__N_1602[68]), .S1(d8_71__N_1602[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1044_35.INIT0 = 16'hb874;
    defparam add_1044_35.INIT1 = 16'hb874;
    defparam add_1044_35.INJECT1_0 = "NO";
    defparam add_1044_35.INJECT1_1 = "NO";
    CCU2D add_1044_33 (.A0(d_d7[66]), .B0(n5862), .C0(n5863[30]), .D0(d7[66]), 
          .A1(d_d7[67]), .B1(n5862), .C1(n5863[31]), .D1(d7[67]), .CIN(n11645), 
          .COUT(n11646), .S0(d8_71__N_1602[66]), .S1(d8_71__N_1602[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1044_33.INIT0 = 16'hb874;
    defparam add_1044_33.INIT1 = 16'hb874;
    defparam add_1044_33.INJECT1_0 = "NO";
    defparam add_1044_33.INJECT1_1 = "NO";
    CCU2D add_1044_31 (.A0(d_d7[64]), .B0(n5862), .C0(n5863[28]), .D0(d7[64]), 
          .A1(d_d7[65]), .B1(n5862), .C1(n5863[29]), .D1(d7[65]), .CIN(n11644), 
          .COUT(n11645), .S0(d8_71__N_1602[64]), .S1(d8_71__N_1602[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1044_31.INIT0 = 16'hb874;
    defparam add_1044_31.INIT1 = 16'hb874;
    defparam add_1044_31.INJECT1_0 = "NO";
    defparam add_1044_31.INJECT1_1 = "NO";
    CCU2D add_1044_29 (.A0(d_d7[62]), .B0(n5862), .C0(n5863[26]), .D0(d7[62]), 
          .A1(d_d7[63]), .B1(n5862), .C1(n5863[27]), .D1(d7[63]), .CIN(n11643), 
          .COUT(n11644), .S0(d8_71__N_1602[62]), .S1(d8_71__N_1602[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1044_29.INIT0 = 16'hb874;
    defparam add_1044_29.INIT1 = 16'hb874;
    defparam add_1044_29.INJECT1_0 = "NO";
    defparam add_1044_29.INJECT1_1 = "NO";
    CCU2D add_1044_27 (.A0(d_d7[60]), .B0(n5862), .C0(n5863[24]), .D0(d7[60]), 
          .A1(d_d7[61]), .B1(n5862), .C1(n5863[25]), .D1(d7[61]), .CIN(n11642), 
          .COUT(n11643), .S0(d8_71__N_1602[60]), .S1(d8_71__N_1602[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1044_27.INIT0 = 16'hb874;
    defparam add_1044_27.INIT1 = 16'hb874;
    defparam add_1044_27.INJECT1_0 = "NO";
    defparam add_1044_27.INJECT1_1 = "NO";
    CCU2D add_1044_25 (.A0(d_d7[58]), .B0(n5862), .C0(n5863[22]), .D0(d7[58]), 
          .A1(d_d7[59]), .B1(n5862), .C1(n5863[23]), .D1(d7[59]), .CIN(n11641), 
          .COUT(n11642), .S0(d8_71__N_1602[58]), .S1(d8_71__N_1602[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1044_25.INIT0 = 16'hb874;
    defparam add_1044_25.INIT1 = 16'hb874;
    defparam add_1044_25.INJECT1_0 = "NO";
    defparam add_1044_25.INJECT1_1 = "NO";
    CCU2D add_1044_23 (.A0(d_d7[56]), .B0(n5862), .C0(n5863[20]), .D0(d7[56]), 
          .A1(d_d7[57]), .B1(n5862), .C1(n5863[21]), .D1(d7[57]), .CIN(n11640), 
          .COUT(n11641), .S0(d8_71__N_1602[56]), .S1(d8_71__N_1602[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1044_23.INIT0 = 16'hb874;
    defparam add_1044_23.INIT1 = 16'hb874;
    defparam add_1044_23.INJECT1_0 = "NO";
    defparam add_1044_23.INJECT1_1 = "NO";
    CCU2D add_1044_21 (.A0(d_d7[54]), .B0(n5862), .C0(n5863[18]), .D0(d7[54]), 
          .A1(d_d7[55]), .B1(n5862), .C1(n5863[19]), .D1(d7[55]), .CIN(n11639), 
          .COUT(n11640), .S0(d8_71__N_1602[54]), .S1(d8_71__N_1602[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1044_21.INIT0 = 16'hb874;
    defparam add_1044_21.INIT1 = 16'hb874;
    defparam add_1044_21.INJECT1_0 = "NO";
    defparam add_1044_21.INJECT1_1 = "NO";
    CCU2D add_1044_19 (.A0(d_d7[52]), .B0(n5862), .C0(n5863[16]), .D0(d7[52]), 
          .A1(d_d7[53]), .B1(n5862), .C1(n5863[17]), .D1(d7[53]), .CIN(n11638), 
          .COUT(n11639), .S0(d8_71__N_1602[52]), .S1(d8_71__N_1602[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1044_19.INIT0 = 16'hb874;
    defparam add_1044_19.INIT1 = 16'hb874;
    defparam add_1044_19.INJECT1_0 = "NO";
    defparam add_1044_19.INJECT1_1 = "NO";
    CCU2D add_1044_17 (.A0(d_d7[50]), .B0(n5862), .C0(n5863[14]), .D0(d7[50]), 
          .A1(d_d7[51]), .B1(n5862), .C1(n5863[15]), .D1(d7[51]), .CIN(n11637), 
          .COUT(n11638), .S0(d8_71__N_1602[50]), .S1(d8_71__N_1602[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1044_17.INIT0 = 16'hb874;
    defparam add_1044_17.INIT1 = 16'hb874;
    defparam add_1044_17.INJECT1_0 = "NO";
    defparam add_1044_17.INJECT1_1 = "NO";
    CCU2D add_1044_15 (.A0(d_d7[48]), .B0(n5862), .C0(n5863[12]), .D0(d7[48]), 
          .A1(d_d7[49]), .B1(n5862), .C1(n5863[13]), .D1(d7[49]), .CIN(n11636), 
          .COUT(n11637), .S0(d8_71__N_1602[48]), .S1(d8_71__N_1602[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1044_15.INIT0 = 16'hb874;
    defparam add_1044_15.INIT1 = 16'hb874;
    defparam add_1044_15.INJECT1_0 = "NO";
    defparam add_1044_15.INJECT1_1 = "NO";
    CCU2D add_1044_13 (.A0(d_d7[46]), .B0(n5862), .C0(n5863[10]), .D0(d7[46]), 
          .A1(d_d7[47]), .B1(n5862), .C1(n5863[11]), .D1(d7[47]), .CIN(n11635), 
          .COUT(n11636), .S0(d8_71__N_1602[46]), .S1(d8_71__N_1602[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1044_13.INIT0 = 16'hb874;
    defparam add_1044_13.INIT1 = 16'hb874;
    defparam add_1044_13.INJECT1_0 = "NO";
    defparam add_1044_13.INJECT1_1 = "NO";
    CCU2D add_1044_11 (.A0(d_d7[44]), .B0(n5862), .C0(n5863[8]), .D0(d7[44]), 
          .A1(d_d7[45]), .B1(n5862), .C1(n5863[9]), .D1(d7[45]), .CIN(n11634), 
          .COUT(n11635), .S0(d8_71__N_1602[44]), .S1(d8_71__N_1602[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1044_11.INIT0 = 16'hb874;
    defparam add_1044_11.INIT1 = 16'hb874;
    defparam add_1044_11.INJECT1_0 = "NO";
    defparam add_1044_11.INJECT1_1 = "NO";
    CCU2D add_1044_9 (.A0(d_d7[42]), .B0(n5862), .C0(n5863[6]), .D0(d7[42]), 
          .A1(d_d7[43]), .B1(n5862), .C1(n5863[7]), .D1(d7[43]), .CIN(n11633), 
          .COUT(n11634), .S0(d8_71__N_1602[42]), .S1(d8_71__N_1602[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1044_9.INIT0 = 16'hb874;
    defparam add_1044_9.INIT1 = 16'hb874;
    defparam add_1044_9.INJECT1_0 = "NO";
    defparam add_1044_9.INJECT1_1 = "NO";
    CCU2D add_1044_7 (.A0(d_d7[40]), .B0(n5862), .C0(n5863[4]), .D0(d7[40]), 
          .A1(d_d7[41]), .B1(n5862), .C1(n5863[5]), .D1(d7[41]), .CIN(n11632), 
          .COUT(n11633), .S0(d8_71__N_1602[40]), .S1(d8_71__N_1602[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1044_7.INIT0 = 16'hb874;
    defparam add_1044_7.INIT1 = 16'hb874;
    defparam add_1044_7.INJECT1_0 = "NO";
    defparam add_1044_7.INJECT1_1 = "NO";
    CCU2D add_1044_5 (.A0(d_d7[38]), .B0(n5862), .C0(n5863[2]), .D0(d7[38]), 
          .A1(d_d7[39]), .B1(n5862), .C1(n5863[3]), .D1(d7[39]), .CIN(n11631), 
          .COUT(n11632), .S0(d8_71__N_1602[38]), .S1(d8_71__N_1602[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1044_5.INIT0 = 16'hb874;
    defparam add_1044_5.INIT1 = 16'hb874;
    defparam add_1044_5.INJECT1_0 = "NO";
    defparam add_1044_5.INJECT1_1 = "NO";
    CCU2D add_1044_3 (.A0(d_d7[36]), .B0(n5862), .C0(n5863[0]), .D0(d7[36]), 
          .A1(d_d7[37]), .B1(n5862), .C1(n5863[1]), .D1(d7[37]), .CIN(n11630), 
          .COUT(n11631), .S0(d8_71__N_1602[36]), .S1(d8_71__N_1602[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1044_3.INIT0 = 16'hb874;
    defparam add_1044_3.INIT1 = 16'hb874;
    defparam add_1044_3.INJECT1_0 = "NO";
    defparam add_1044_3.INJECT1_1 = "NO";
    CCU2D add_1044_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5862), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11630));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(109[17:26])
    defparam add_1044_1.INIT0 = 16'hF000;
    defparam add_1044_1.INIT1 = 16'h0555;
    defparam add_1044_1.INJECT1_0 = "NO";
    defparam add_1044_1.INJECT1_1 = "NO";
    CCU2D add_1048_37 (.A0(d6[71]), .B0(d_d6[71]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n11488), 
          .S0(n6015[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1048_37.INIT0 = 16'h5999;
    defparam add_1048_37.INIT1 = 16'h0000;
    defparam add_1048_37.INJECT1_0 = "NO";
    defparam add_1048_37.INJECT1_1 = "NO";
    CCU2D add_1048_35 (.A0(d6[69]), .B0(d_d6[69]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[70]), .B1(d_d6[70]), .C1(GND_net), .D1(GND_net), .CIN(n11487), 
          .COUT(n11488), .S0(n6015[33]), .S1(n6015[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1048_35.INIT0 = 16'h5999;
    defparam add_1048_35.INIT1 = 16'h5999;
    defparam add_1048_35.INJECT1_0 = "NO";
    defparam add_1048_35.INJECT1_1 = "NO";
    CCU2D add_1048_33 (.A0(d6[67]), .B0(d_d6[67]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[68]), .B1(d_d6[68]), .C1(GND_net), .D1(GND_net), .CIN(n11486), 
          .COUT(n11487), .S0(n6015[31]), .S1(n6015[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1048_33.INIT0 = 16'h5999;
    defparam add_1048_33.INIT1 = 16'h5999;
    defparam add_1048_33.INJECT1_0 = "NO";
    defparam add_1048_33.INJECT1_1 = "NO";
    CCU2D add_1048_31 (.A0(d6[65]), .B0(d_d6[65]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[66]), .B1(d_d6[66]), .C1(GND_net), .D1(GND_net), .CIN(n11485), 
          .COUT(n11486), .S0(n6015[29]), .S1(n6015[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1048_31.INIT0 = 16'h5999;
    defparam add_1048_31.INIT1 = 16'h5999;
    defparam add_1048_31.INJECT1_0 = "NO";
    defparam add_1048_31.INJECT1_1 = "NO";
    CCU2D add_1048_29 (.A0(d6[63]), .B0(d_d6[63]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[64]), .B1(d_d6[64]), .C1(GND_net), .D1(GND_net), .CIN(n11484), 
          .COUT(n11485), .S0(n6015[27]), .S1(n6015[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1048_29.INIT0 = 16'h5999;
    defparam add_1048_29.INIT1 = 16'h5999;
    defparam add_1048_29.INJECT1_0 = "NO";
    defparam add_1048_29.INJECT1_1 = "NO";
    CCU2D add_1048_27 (.A0(d6[61]), .B0(d_d6[61]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[62]), .B1(d_d6[62]), .C1(GND_net), .D1(GND_net), .CIN(n11483), 
          .COUT(n11484), .S0(n6015[25]), .S1(n6015[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1048_27.INIT0 = 16'h5999;
    defparam add_1048_27.INIT1 = 16'h5999;
    defparam add_1048_27.INJECT1_0 = "NO";
    defparam add_1048_27.INJECT1_1 = "NO";
    CCU2D add_1048_25 (.A0(d6[59]), .B0(d_d6[59]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[60]), .B1(d_d6[60]), .C1(GND_net), .D1(GND_net), .CIN(n11482), 
          .COUT(n11483), .S0(n6015[23]), .S1(n6015[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1048_25.INIT0 = 16'h5999;
    defparam add_1048_25.INIT1 = 16'h5999;
    defparam add_1048_25.INJECT1_0 = "NO";
    defparam add_1048_25.INJECT1_1 = "NO";
    CCU2D add_1048_23 (.A0(d6[57]), .B0(d_d6[57]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[58]), .B1(d_d6[58]), .C1(GND_net), .D1(GND_net), .CIN(n11481), 
          .COUT(n11482), .S0(n6015[21]), .S1(n6015[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1048_23.INIT0 = 16'h5999;
    defparam add_1048_23.INIT1 = 16'h5999;
    defparam add_1048_23.INJECT1_0 = "NO";
    defparam add_1048_23.INJECT1_1 = "NO";
    CCU2D add_1048_21 (.A0(d6[55]), .B0(d_d6[55]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[56]), .B1(d_d6[56]), .C1(GND_net), .D1(GND_net), .CIN(n11480), 
          .COUT(n11481), .S0(n6015[19]), .S1(n6015[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1048_21.INIT0 = 16'h5999;
    defparam add_1048_21.INIT1 = 16'h5999;
    defparam add_1048_21.INJECT1_0 = "NO";
    defparam add_1048_21.INJECT1_1 = "NO";
    CCU2D add_1048_19 (.A0(d6[53]), .B0(d_d6[53]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[54]), .B1(d_d6[54]), .C1(GND_net), .D1(GND_net), .CIN(n11479), 
          .COUT(n11480), .S0(n6015[17]), .S1(n6015[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1048_19.INIT0 = 16'h5999;
    defparam add_1048_19.INIT1 = 16'h5999;
    defparam add_1048_19.INJECT1_0 = "NO";
    defparam add_1048_19.INJECT1_1 = "NO";
    CCU2D add_1048_17 (.A0(d6[51]), .B0(d_d6[51]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[52]), .B1(d_d6[52]), .C1(GND_net), .D1(GND_net), .CIN(n11478), 
          .COUT(n11479), .S0(n6015[15]), .S1(n6015[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1048_17.INIT0 = 16'h5999;
    defparam add_1048_17.INIT1 = 16'h5999;
    defparam add_1048_17.INJECT1_0 = "NO";
    defparam add_1048_17.INJECT1_1 = "NO";
    CCU2D add_1048_15 (.A0(d6[49]), .B0(d_d6[49]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[50]), .B1(d_d6[50]), .C1(GND_net), .D1(GND_net), .CIN(n11477), 
          .COUT(n11478), .S0(n6015[13]), .S1(n6015[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1048_15.INIT0 = 16'h5999;
    defparam add_1048_15.INIT1 = 16'h5999;
    defparam add_1048_15.INJECT1_0 = "NO";
    defparam add_1048_15.INJECT1_1 = "NO";
    CCU2D add_1048_13 (.A0(d6[47]), .B0(d_d6[47]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[48]), .B1(d_d6[48]), .C1(GND_net), .D1(GND_net), .CIN(n11476), 
          .COUT(n11477), .S0(n6015[11]), .S1(n6015[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1048_13.INIT0 = 16'h5999;
    defparam add_1048_13.INIT1 = 16'h5999;
    defparam add_1048_13.INJECT1_0 = "NO";
    defparam add_1048_13.INJECT1_1 = "NO";
    CCU2D add_1048_11 (.A0(d6[45]), .B0(d_d6[45]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[46]), .B1(d_d6[46]), .C1(GND_net), .D1(GND_net), .CIN(n11475), 
          .COUT(n11476), .S0(n6015[9]), .S1(n6015[10]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1048_11.INIT0 = 16'h5999;
    defparam add_1048_11.INIT1 = 16'h5999;
    defparam add_1048_11.INJECT1_0 = "NO";
    defparam add_1048_11.INJECT1_1 = "NO";
    CCU2D add_1048_9 (.A0(d6[43]), .B0(d_d6[43]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[44]), .B1(d_d6[44]), .C1(GND_net), .D1(GND_net), .CIN(n11474), 
          .COUT(n11475), .S0(n6015[7]), .S1(n6015[8]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1048_9.INIT0 = 16'h5999;
    defparam add_1048_9.INIT1 = 16'h5999;
    defparam add_1048_9.INJECT1_0 = "NO";
    defparam add_1048_9.INJECT1_1 = "NO";
    CCU2D add_1048_7 (.A0(d6[41]), .B0(d_d6[41]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[42]), .B1(d_d6[42]), .C1(GND_net), .D1(GND_net), .CIN(n11473), 
          .COUT(n11474), .S0(n6015[5]), .S1(n6015[6]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1048_7.INIT0 = 16'h5999;
    defparam add_1048_7.INIT1 = 16'h5999;
    defparam add_1048_7.INJECT1_0 = "NO";
    defparam add_1048_7.INJECT1_1 = "NO";
    CCU2D add_1048_5 (.A0(d6[39]), .B0(d_d6[39]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[40]), .B1(d_d6[40]), .C1(GND_net), .D1(GND_net), .CIN(n11472), 
          .COUT(n11473), .S0(n6015[3]), .S1(n6015[4]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1048_5.INIT0 = 16'h5999;
    defparam add_1048_5.INIT1 = 16'h5999;
    defparam add_1048_5.INJECT1_0 = "NO";
    defparam add_1048_5.INJECT1_1 = "NO";
    CCU2D add_1048_3 (.A0(d6[37]), .B0(d_d6[37]), .C0(GND_net), .D0(GND_net), 
          .A1(d6[38]), .B1(d_d6[38]), .C1(GND_net), .D1(GND_net), .CIN(n11471), 
          .COUT(n11472), .S0(n6015[1]), .S1(n6015[2]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1048_3.INIT0 = 16'h5999;
    defparam add_1048_3.INIT1 = 16'h5999;
    defparam add_1048_3.INJECT1_0 = "NO";
    defparam add_1048_3.INJECT1_1 = "NO";
    CCU2D add_1048_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d6[36]), .B1(d_d6[36]), .C1(GND_net), .D1(GND_net), .COUT(n11471), 
          .S1(n6015[0]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1048_1.INIT0 = 16'hF000;
    defparam add_1048_1.INIT1 = 16'h5999;
    defparam add_1048_1.INJECT1_0 = "NO";
    defparam add_1048_1.INJECT1_1 = "NO";
    CCU2D add_1049_37 (.A0(d_d6[70]), .B0(n6014), .C0(n6015[34]), .D0(d6[70]), 
          .A1(d_d6[71]), .B1(n6014), .C1(n6015[35]), .D1(d6[71]), .CIN(n11469), 
          .S0(d7_71__N_1530[70]), .S1(d7_71__N_1530[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1049_37.INIT0 = 16'hb874;
    defparam add_1049_37.INIT1 = 16'hb874;
    defparam add_1049_37.INJECT1_0 = "NO";
    defparam add_1049_37.INJECT1_1 = "NO";
    CCU2D add_1049_35 (.A0(d_d6[68]), .B0(n6014), .C0(n6015[32]), .D0(d6[68]), 
          .A1(d_d6[69]), .B1(n6014), .C1(n6015[33]), .D1(d6[69]), .CIN(n11468), 
          .COUT(n11469), .S0(d7_71__N_1530[68]), .S1(d7_71__N_1530[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1049_35.INIT0 = 16'hb874;
    defparam add_1049_35.INIT1 = 16'hb874;
    defparam add_1049_35.INJECT1_0 = "NO";
    defparam add_1049_35.INJECT1_1 = "NO";
    CCU2D add_1049_33 (.A0(d_d6[66]), .B0(n6014), .C0(n6015[30]), .D0(d6[66]), 
          .A1(d_d6[67]), .B1(n6014), .C1(n6015[31]), .D1(d6[67]), .CIN(n11467), 
          .COUT(n11468), .S0(d7_71__N_1530[66]), .S1(d7_71__N_1530[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1049_33.INIT0 = 16'hb874;
    defparam add_1049_33.INIT1 = 16'hb874;
    defparam add_1049_33.INJECT1_0 = "NO";
    defparam add_1049_33.INJECT1_1 = "NO";
    CCU2D add_1049_31 (.A0(d_d6[64]), .B0(n6014), .C0(n6015[28]), .D0(d6[64]), 
          .A1(d_d6[65]), .B1(n6014), .C1(n6015[29]), .D1(d6[65]), .CIN(n11466), 
          .COUT(n11467), .S0(d7_71__N_1530[64]), .S1(d7_71__N_1530[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1049_31.INIT0 = 16'hb874;
    defparam add_1049_31.INIT1 = 16'hb874;
    defparam add_1049_31.INJECT1_0 = "NO";
    defparam add_1049_31.INJECT1_1 = "NO";
    CCU2D add_1049_29 (.A0(d_d6[62]), .B0(n6014), .C0(n6015[26]), .D0(d6[62]), 
          .A1(d_d6[63]), .B1(n6014), .C1(n6015[27]), .D1(d6[63]), .CIN(n11465), 
          .COUT(n11466), .S0(d7_71__N_1530[62]), .S1(d7_71__N_1530[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1049_29.INIT0 = 16'hb874;
    defparam add_1049_29.INIT1 = 16'hb874;
    defparam add_1049_29.INJECT1_0 = "NO";
    defparam add_1049_29.INJECT1_1 = "NO";
    CCU2D add_1049_27 (.A0(d_d6[60]), .B0(n6014), .C0(n6015[24]), .D0(d6[60]), 
          .A1(d_d6[61]), .B1(n6014), .C1(n6015[25]), .D1(d6[61]), .CIN(n11464), 
          .COUT(n11465), .S0(d7_71__N_1530[60]), .S1(d7_71__N_1530[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1049_27.INIT0 = 16'hb874;
    defparam add_1049_27.INIT1 = 16'hb874;
    defparam add_1049_27.INJECT1_0 = "NO";
    defparam add_1049_27.INJECT1_1 = "NO";
    CCU2D add_1049_25 (.A0(d_d6[58]), .B0(n6014), .C0(n6015[22]), .D0(d6[58]), 
          .A1(d_d6[59]), .B1(n6014), .C1(n6015[23]), .D1(d6[59]), .CIN(n11463), 
          .COUT(n11464), .S0(d7_71__N_1530[58]), .S1(d7_71__N_1530[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1049_25.INIT0 = 16'hb874;
    defparam add_1049_25.INIT1 = 16'hb874;
    defparam add_1049_25.INJECT1_0 = "NO";
    defparam add_1049_25.INJECT1_1 = "NO";
    CCU2D add_1049_23 (.A0(d_d6[56]), .B0(n6014), .C0(n6015[20]), .D0(d6[56]), 
          .A1(d_d6[57]), .B1(n6014), .C1(n6015[21]), .D1(d6[57]), .CIN(n11462), 
          .COUT(n11463), .S0(d7_71__N_1530[56]), .S1(d7_71__N_1530[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1049_23.INIT0 = 16'hb874;
    defparam add_1049_23.INIT1 = 16'hb874;
    defparam add_1049_23.INJECT1_0 = "NO";
    defparam add_1049_23.INJECT1_1 = "NO";
    CCU2D add_1049_21 (.A0(d_d6[54]), .B0(n6014), .C0(n6015[18]), .D0(d6[54]), 
          .A1(d_d6[55]), .B1(n6014), .C1(n6015[19]), .D1(d6[55]), .CIN(n11461), 
          .COUT(n11462), .S0(d7_71__N_1530[54]), .S1(d7_71__N_1530[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1049_21.INIT0 = 16'hb874;
    defparam add_1049_21.INIT1 = 16'hb874;
    defparam add_1049_21.INJECT1_0 = "NO";
    defparam add_1049_21.INJECT1_1 = "NO";
    CCU2D add_1049_19 (.A0(d_d6[52]), .B0(n6014), .C0(n6015[16]), .D0(d6[52]), 
          .A1(d_d6[53]), .B1(n6014), .C1(n6015[17]), .D1(d6[53]), .CIN(n11460), 
          .COUT(n11461), .S0(d7_71__N_1530[52]), .S1(d7_71__N_1530[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1049_19.INIT0 = 16'hb874;
    defparam add_1049_19.INIT1 = 16'hb874;
    defparam add_1049_19.INJECT1_0 = "NO";
    defparam add_1049_19.INJECT1_1 = "NO";
    CCU2D add_1049_17 (.A0(d_d6[50]), .B0(n6014), .C0(n6015[14]), .D0(d6[50]), 
          .A1(d_d6[51]), .B1(n6014), .C1(n6015[15]), .D1(d6[51]), .CIN(n11459), 
          .COUT(n11460), .S0(d7_71__N_1530[50]), .S1(d7_71__N_1530[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1049_17.INIT0 = 16'hb874;
    defparam add_1049_17.INIT1 = 16'hb874;
    defparam add_1049_17.INJECT1_0 = "NO";
    defparam add_1049_17.INJECT1_1 = "NO";
    CCU2D add_1049_15 (.A0(d_d6[48]), .B0(n6014), .C0(n6015[12]), .D0(d6[48]), 
          .A1(d_d6[49]), .B1(n6014), .C1(n6015[13]), .D1(d6[49]), .CIN(n11458), 
          .COUT(n11459), .S0(d7_71__N_1530[48]), .S1(d7_71__N_1530[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1049_15.INIT0 = 16'hb874;
    defparam add_1049_15.INIT1 = 16'hb874;
    defparam add_1049_15.INJECT1_0 = "NO";
    defparam add_1049_15.INJECT1_1 = "NO";
    CCU2D add_1049_13 (.A0(d_d6[46]), .B0(n6014), .C0(n6015[10]), .D0(d6[46]), 
          .A1(d_d6[47]), .B1(n6014), .C1(n6015[11]), .D1(d6[47]), .CIN(n11457), 
          .COUT(n11458), .S0(d7_71__N_1530[46]), .S1(d7_71__N_1530[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1049_13.INIT0 = 16'hb874;
    defparam add_1049_13.INIT1 = 16'hb874;
    defparam add_1049_13.INJECT1_0 = "NO";
    defparam add_1049_13.INJECT1_1 = "NO";
    CCU2D add_1049_11 (.A0(d_d6[44]), .B0(n6014), .C0(n6015[8]), .D0(d6[44]), 
          .A1(d_d6[45]), .B1(n6014), .C1(n6015[9]), .D1(d6[45]), .CIN(n11456), 
          .COUT(n11457), .S0(d7_71__N_1530[44]), .S1(d7_71__N_1530[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1049_11.INIT0 = 16'hb874;
    defparam add_1049_11.INIT1 = 16'hb874;
    defparam add_1049_11.INJECT1_0 = "NO";
    defparam add_1049_11.INJECT1_1 = "NO";
    CCU2D add_1049_9 (.A0(d_d6[42]), .B0(n6014), .C0(n6015[6]), .D0(d6[42]), 
          .A1(d_d6[43]), .B1(n6014), .C1(n6015[7]), .D1(d6[43]), .CIN(n11455), 
          .COUT(n11456), .S0(d7_71__N_1530[42]), .S1(d7_71__N_1530[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1049_9.INIT0 = 16'hb874;
    defparam add_1049_9.INIT1 = 16'hb874;
    defparam add_1049_9.INJECT1_0 = "NO";
    defparam add_1049_9.INJECT1_1 = "NO";
    CCU2D add_1049_7 (.A0(d_d6[40]), .B0(n6014), .C0(n6015[4]), .D0(d6[40]), 
          .A1(d_d6[41]), .B1(n6014), .C1(n6015[5]), .D1(d6[41]), .CIN(n11454), 
          .COUT(n11455), .S0(d7_71__N_1530[40]), .S1(d7_71__N_1530[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1049_7.INIT0 = 16'hb874;
    defparam add_1049_7.INIT1 = 16'hb874;
    defparam add_1049_7.INJECT1_0 = "NO";
    defparam add_1049_7.INJECT1_1 = "NO";
    CCU2D add_1049_5 (.A0(d_d6[38]), .B0(n6014), .C0(n6015[2]), .D0(d6[38]), 
          .A1(d_d6[39]), .B1(n6014), .C1(n6015[3]), .D1(d6[39]), .CIN(n11453), 
          .COUT(n11454), .S0(d7_71__N_1530[38]), .S1(d7_71__N_1530[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1049_5.INIT0 = 16'hb874;
    defparam add_1049_5.INIT1 = 16'hb874;
    defparam add_1049_5.INJECT1_0 = "NO";
    defparam add_1049_5.INJECT1_1 = "NO";
    CCU2D add_1049_3 (.A0(d_d6[36]), .B0(n6014), .C0(n6015[0]), .D0(d6[36]), 
          .A1(d_d6[37]), .B1(n6014), .C1(n6015[1]), .D1(d6[37]), .CIN(n11452), 
          .COUT(n11453), .S0(d7_71__N_1530[36]), .S1(d7_71__N_1530[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1049_3.INIT0 = 16'hb874;
    defparam add_1049_3.INIT1 = 16'hb874;
    defparam add_1049_3.INJECT1_0 = "NO";
    defparam add_1049_3.INJECT1_1 = "NO";
    CCU2D add_1049_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n6014), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11452));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(106[17:26])
    defparam add_1049_1.INIT0 = 16'hF000;
    defparam add_1049_1.INIT1 = 16'h0555;
    defparam add_1049_1.INJECT1_0 = "NO";
    defparam add_1049_1.INJECT1_1 = "NO";
    CCU2D add_1053_37 (.A0(d_tmp[71]), .B0(d_d_tmp[71]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n11448), .S0(n6167[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1053_37.INIT0 = 16'h5999;
    defparam add_1053_37.INIT1 = 16'h0000;
    defparam add_1053_37.INJECT1_0 = "NO";
    defparam add_1053_37.INJECT1_1 = "NO";
    CCU2D add_1053_35 (.A0(d_tmp[69]), .B0(d_d_tmp[69]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[70]), .B1(d_d_tmp[70]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11447), .COUT(n11448), .S0(n6167[33]), 
          .S1(n6167[34]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1053_35.INIT0 = 16'h5999;
    defparam add_1053_35.INIT1 = 16'h5999;
    defparam add_1053_35.INJECT1_0 = "NO";
    defparam add_1053_35.INJECT1_1 = "NO";
    CCU2D add_1053_33 (.A0(d_tmp[67]), .B0(d_d_tmp[67]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[68]), .B1(d_d_tmp[68]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11446), .COUT(n11447), .S0(n6167[31]), 
          .S1(n6167[32]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1053_33.INIT0 = 16'h5999;
    defparam add_1053_33.INIT1 = 16'h5999;
    defparam add_1053_33.INJECT1_0 = "NO";
    defparam add_1053_33.INJECT1_1 = "NO";
    CCU2D add_1053_31 (.A0(d_tmp[65]), .B0(d_d_tmp[65]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[66]), .B1(d_d_tmp[66]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11445), .COUT(n11446), .S0(n6167[29]), 
          .S1(n6167[30]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1053_31.INIT0 = 16'h5999;
    defparam add_1053_31.INIT1 = 16'h5999;
    defparam add_1053_31.INJECT1_0 = "NO";
    defparam add_1053_31.INJECT1_1 = "NO";
    CCU2D add_1053_29 (.A0(d_tmp[63]), .B0(d_d_tmp[63]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[64]), .B1(d_d_tmp[64]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11444), .COUT(n11445), .S0(n6167[27]), 
          .S1(n6167[28]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1053_29.INIT0 = 16'h5999;
    defparam add_1053_29.INIT1 = 16'h5999;
    defparam add_1053_29.INJECT1_0 = "NO";
    defparam add_1053_29.INJECT1_1 = "NO";
    CCU2D add_1053_27 (.A0(d_tmp[61]), .B0(d_d_tmp[61]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[62]), .B1(d_d_tmp[62]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11443), .COUT(n11444), .S0(n6167[25]), 
          .S1(n6167[26]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1053_27.INIT0 = 16'h5999;
    defparam add_1053_27.INIT1 = 16'h5999;
    defparam add_1053_27.INJECT1_0 = "NO";
    defparam add_1053_27.INJECT1_1 = "NO";
    CCU2D add_1053_25 (.A0(d_tmp[59]), .B0(d_d_tmp[59]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[60]), .B1(d_d_tmp[60]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11442), .COUT(n11443), .S0(n6167[23]), 
          .S1(n6167[24]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1053_25.INIT0 = 16'h5999;
    defparam add_1053_25.INIT1 = 16'h5999;
    defparam add_1053_25.INJECT1_0 = "NO";
    defparam add_1053_25.INJECT1_1 = "NO";
    CCU2D add_1053_23 (.A0(d_tmp[57]), .B0(d_d_tmp[57]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[58]), .B1(d_d_tmp[58]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11441), .COUT(n11442), .S0(n6167[21]), 
          .S1(n6167[22]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1053_23.INIT0 = 16'h5999;
    defparam add_1053_23.INIT1 = 16'h5999;
    defparam add_1053_23.INJECT1_0 = "NO";
    defparam add_1053_23.INJECT1_1 = "NO";
    CCU2D add_1053_21 (.A0(d_tmp[55]), .B0(d_d_tmp[55]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[56]), .B1(d_d_tmp[56]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11440), .COUT(n11441), .S0(n6167[19]), 
          .S1(n6167[20]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1053_21.INIT0 = 16'h5999;
    defparam add_1053_21.INIT1 = 16'h5999;
    defparam add_1053_21.INJECT1_0 = "NO";
    defparam add_1053_21.INJECT1_1 = "NO";
    CCU2D add_1053_19 (.A0(d_tmp[53]), .B0(d_d_tmp[53]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[54]), .B1(d_d_tmp[54]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11439), .COUT(n11440), .S0(n6167[17]), 
          .S1(n6167[18]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1053_19.INIT0 = 16'h5999;
    defparam add_1053_19.INIT1 = 16'h5999;
    defparam add_1053_19.INJECT1_0 = "NO";
    defparam add_1053_19.INJECT1_1 = "NO";
    CCU2D add_1053_17 (.A0(d_tmp[51]), .B0(d_d_tmp[51]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[52]), .B1(d_d_tmp[52]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11438), .COUT(n11439), .S0(n6167[15]), 
          .S1(n6167[16]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1053_17.INIT0 = 16'h5999;
    defparam add_1053_17.INIT1 = 16'h5999;
    defparam add_1053_17.INJECT1_0 = "NO";
    defparam add_1053_17.INJECT1_1 = "NO";
    CCU2D add_1053_15 (.A0(d_tmp[49]), .B0(d_d_tmp[49]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[50]), .B1(d_d_tmp[50]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11437), .COUT(n11438), .S0(n6167[13]), 
          .S1(n6167[14]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1053_15.INIT0 = 16'h5999;
    defparam add_1053_15.INIT1 = 16'h5999;
    defparam add_1053_15.INJECT1_0 = "NO";
    defparam add_1053_15.INJECT1_1 = "NO";
    CCU2D add_1053_13 (.A0(d_tmp[47]), .B0(d_d_tmp[47]), .C0(GND_net), 
          .D0(GND_net), .A1(d_tmp[48]), .B1(d_d_tmp[48]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11436), .COUT(n11437), .S0(n6167[11]), 
          .S1(n6167[12]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(103[17:32])
    defparam add_1053_13.INIT0 = 16'h5999;
    defparam add_1053_13.INIT1 = 16'h5999;
    defparam add_1053_13.INJECT1_0 = "NO";
    defparam add_1053_13.INJECT1_1 = "NO";
    FD1S3AX v_comb_66_rep_201 (.D(osc_clk_enable_743), .CK(osc_clk), .Q(osc_clk_enable_833)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_201.GSR = "ENABLED";
    LUT4 mux_1207_i2_3_lut (.A(n6775[21]), .B(n6813[21]), .C(n6774), .Z(d10_71__N_1746[57])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1207_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1207_i3_3_lut (.A(n6775[22]), .B(n6813[22]), .C(n6774), .Z(d10_71__N_1746[58])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1207_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1207_i4_3_lut (.A(n6775[23]), .B(n6813[23]), .C(n6774), .Z(d10_71__N_1746[59])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1207_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1207_i5_3_lut (.A(n6775[24]), .B(n6813[24]), .C(n6774), .Z(d10_71__N_1746[60])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1207_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1207_i6_3_lut (.A(n6775[25]), .B(n6813[25]), .C(n6774), .Z(d10_71__N_1746[61])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1207_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1207_i7_3_lut (.A(n6775[26]), .B(n6813[26]), .C(n6774), .Z(d10_71__N_1746[62])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1207_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1207_i8_3_lut (.A(n6775[27]), .B(n6813[27]), .C(n6774), .Z(d10_71__N_1746[63])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1207_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1207_i9_3_lut (.A(n6775[28]), .B(n6813[28]), .C(n6774), .Z(d10_71__N_1746[64])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1207_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1207_i10_3_lut (.A(n6775[29]), .B(n6813[29]), .C(n6774), 
         .Z(d10_71__N_1746[65])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1207_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1207_i11_3_lut (.A(n6775[30]), .B(n6813[30]), .C(n6774), 
         .Z(d10_71__N_1746[66])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1207_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1207_i12_3_lut (.A(n6775[31]), .B(n6813[31]), .C(n6774), 
         .Z(d10_71__N_1746[67])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1207_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1207_i13_3_lut (.A(n6775[32]), .B(n6813[32]), .C(n6774), 
         .Z(d10_71__N_1746[68])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1207_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1207_i14_3_lut (.A(n6775[33]), .B(n6813[33]), .C(n6774), 
         .Z(d10_71__N_1746[69])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1207_i14_3_lut.init = 16'hcaca;
    LUT4 i4800_2_lut (.A(d1[36]), .B(d2[36]), .Z(n4951[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4800_2_lut.init = 16'h6666;
    FD1S3AX v_comb_66_rep_200 (.D(osc_clk_enable_743), .CK(osc_clk), .Q(osc_clk_enable_783)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_200.GSR = "ENABLED";
    LUT4 mux_1207_i15_3_lut (.A(n6775[34]), .B(n6813[34]), .C(n6774), 
         .Z(d10_71__N_1746[70])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1207_i15_3_lut.init = 16'hcaca;
    LUT4 i4794_2_lut (.A(d3[36]), .B(d4[36]), .Z(n5255[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4794_2_lut.init = 16'h6666;
    LUT4 i4754_2_lut (.A(d1[0]), .B(d2[0]), .Z(d2_71__N_489[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4754_2_lut.init = 16'h6666;
    LUT4 mux_1207_i16_3_lut (.A(n6775[35]), .B(n6813[35]), .C(n6774), 
         .Z(d10_71__N_1746[71])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(115[18:27])
    defparam mux_1207_i16_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i62_3_lut (.A(\d10[61] ), .B(\d10[62] ), .C(\CICGain[0] ), 
         .Z(n62)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i62_3_lut.init = 16'hcaca;
    LUT4 i4755_2_lut (.A(d2[0]), .B(d3[0]), .Z(d3_71__N_561[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4755_2_lut.init = 16'h6666;
    LUT4 shift_right_31_i63_3_lut (.A(\d10[62] ), .B(\d10[63] ), .C(\CICGain[0] ), 
         .Z(n63)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i63_3_lut.init = 16'hcaca;
    LUT4 i4756_2_lut (.A(d3[0]), .B(d4[0]), .Z(d4_71__N_633[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4756_2_lut.init = 16'h6666;
    LUT4 shift_right_31_i64_3_lut (.A(\d10[63] ), .B(\d10[64] ), .C(\CICGain[0] ), 
         .Z(n64)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i64_3_lut.init = 16'hcaca;
    LUT4 i4757_2_lut (.A(d4[0]), .B(d5[0]), .Z(d5_71__N_705[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4757_2_lut.init = 16'h6666;
    PFUMX i6060 (.BLUT(n13828), .ALUT(n13829), .C0(\CICGain[0] ), .Z(d_out_11__N_1818[1]));
    LUT4 i5941_then_3_lut (.A(\CICGain[1] ), .B(\d10[59] ), .C(d10[57]), 
         .Z(n13826)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i5941_then_3_lut.init = 16'he4e4;
    LUT4 i5941_else_3_lut (.A(n61), .B(\CICGain[1] ), .C(d10[58]), .Z(n13825)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i5941_else_3_lut.init = 16'he2e2;
    LUT4 shift_right_31_i65_3_lut (.A(\d10[64] ), .B(\d10[65] ), .C(\CICGain[0] ), 
         .Z(n65)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i65_3_lut.init = 16'hcaca;
    LUT4 i4753_2_lut (.A(MixerOutCos[0]), .B(d1[0]), .Z(d1_71__N_417[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4753_2_lut.init = 16'h6666;
    PFUMX i6058 (.BLUT(n13825), .ALUT(n13826), .C0(\CICGain[0] ), .Z(d_out_11__N_1818[0]));
    LUT4 i5849_4_lut_rep_198 (.A(n13248), .B(n13), .C(n13250), .D(n13228), 
         .Z(osc_clk_enable_743)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i5849_4_lut_rep_198.init = 16'h2000;
    LUT4 shift_right_31_i66_3_lut (.A(\d10[65] ), .B(\d10[66] ), .C(\CICGain[0] ), 
         .Z(n66)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i66_3_lut.init = 16'hcaca;
    LUT4 i5997_then_3_lut (.A(\CICGain[1] ), .B(\d10[60] ), .C(d10[58]), 
         .Z(n13829)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i5997_then_3_lut.init = 16'he4e4;
    LUT4 i5997_else_3_lut (.A(n62), .B(\CICGain[1] ), .C(\d10[59] ), .Z(n13828)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i5997_else_3_lut.init = 16'he2e2;
    LUT4 i2670_2_lut (.A(n375[0]), .B(n31), .Z(count_15__N_1441[0])) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(86[13] 89[16])
    defparam i2670_2_lut.init = 16'hbbbb;
    LUT4 shift_right_31_i67_3_lut (.A(\d10[66] ), .B(\d10[67] ), .C(\CICGain[0] ), 
         .Z(n67)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i67_3_lut.init = 16'hcaca;
    LUT4 i11_4_lut (.A(n21), .B(n19), .C(n15), .D(n16), .Z(n31)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i9_4_lut (.A(count[9]), .B(count[3]), .C(count[4]), .D(count[0]), 
         .Z(n21)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 shift_right_31_i68_3_lut (.A(\d10[67] ), .B(\d10[68] ), .C(\CICGain[0] ), 
         .Z(n68)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i68_3_lut.init = 16'hcaca;
    LUT4 i7_4_lut (.A(count[10]), .B(count[1]), .C(count[5]), .D(count[6]), 
         .Z(n19)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 shift_right_31_i70_3_lut (.A(\d10[69] ), .B(\d10[70] ), .C(\CICGain[0] ), 
         .Z(n70)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(119[20:47])
    defparam shift_right_31_i70_3_lut.init = 16'hcaca;
    LUT4 i3_2_lut (.A(count[8]), .B(count[7]), .Z(n15)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(74[11:40])
    defparam i3_2_lut.init = 16'heeee;
    FD1S3AX v_comb_66_rep_212 (.D(osc_clk_enable_743), .CK(osc_clk), .Q(osc_clk_enable_1383)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_212.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_211 (.D(osc_clk_enable_743), .CK(osc_clk), .Q(osc_clk_enable_1333)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_211.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_210 (.D(osc_clk_enable_743), .CK(osc_clk), .Q(osc_clk_enable_1283)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_210.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_209 (.D(osc_clk_enable_743), .CK(osc_clk), .Q(osc_clk_enable_1233)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_209.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_208 (.D(osc_clk_enable_743), .CK(osc_clk), .Q(osc_clk_enable_1183)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_208.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_207 (.D(osc_clk_enable_743), .CK(osc_clk), .Q(osc_clk_enable_1133)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_207.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_206 (.D(osc_clk_enable_743), .CK(osc_clk), .Q(osc_clk_enable_1083)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_206.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_205 (.D(osc_clk_enable_743), .CK(osc_clk), .Q(osc_clk_enable_1033)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_205.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_204 (.D(osc_clk_enable_743), .CK(osc_clk), .Q(osc_clk_enable_983)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_204.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_203 (.D(osc_clk_enable_743), .CK(osc_clk), .Q(osc_clk_enable_933)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_203.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_202 (.D(osc_clk_enable_743), .CK(osc_clk), .Q(osc_clk_enable_883)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam v_comb_66_rep_202.GSR = "ENABLED";
    CCU2D add_1013_6 (.A0(d1[40]), .B0(d2[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[41]), .B1(d2[41]), .C1(GND_net), .D1(GND_net), .CIN(n11894), 
          .COUT(n11895), .S0(n4951[4]), .S1(n4951[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1013_6.INIT0 = 16'h5666;
    defparam add_1013_6.INIT1 = 16'h5666;
    defparam add_1013_6.INJECT1_0 = "NO";
    defparam add_1013_6.INJECT1_1 = "NO";
    CCU2D add_1013_16 (.A0(d1[50]), .B0(d2[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[51]), .B1(d2[51]), .C1(GND_net), .D1(GND_net), .CIN(n11899), 
          .COUT(n11900), .S0(n4951[14]), .S1(n4951[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1013_16.INIT0 = 16'h5666;
    defparam add_1013_16.INIT1 = 16'h5666;
    defparam add_1013_16.INJECT1_0 = "NO";
    defparam add_1013_16.INJECT1_1 = "NO";
    CCU2D add_1013_14 (.A0(d1[48]), .B0(d2[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[49]), .B1(d2[49]), .C1(GND_net), .D1(GND_net), .CIN(n11898), 
          .COUT(n11899), .S0(n4951[12]), .S1(n4951[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1013_14.INIT0 = 16'h5666;
    defparam add_1013_14.INIT1 = 16'h5666;
    defparam add_1013_14.INJECT1_0 = "NO";
    defparam add_1013_14.INJECT1_1 = "NO";
    FD1S3IX count__i2 (.D(n375[2]), .CK(osc_clk), .CD(n8412), .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n375[3]), .CK(osc_clk), .CD(n8412), .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n375[4]), .CK(osc_clk), .CD(n8412), .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n375[5]), .CK(osc_clk), .CD(n8412), .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n375[6]), .CK(osc_clk), .CD(n8412), .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n375[7]), .CK(osc_clk), .CD(n8412), .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n375[8]), .CK(osc_clk), .CD(n8412), .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n375[9]), .CK(osc_clk), .CD(n8412), .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n375[10]), .CK(osc_clk), .CD(n8412), .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_15__N_1441[11]), .CK(osc_clk), .CD(count_15__N_1457), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(n375[12]), .CK(osc_clk), .CD(n8412), .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(n375[13]), .CK(osc_clk), .CD(n8412), .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(n375[14]), .CK(osc_clk), .CD(n8412), .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(n375[15]), .CK(osc_clk), .CD(n8412), .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=2, LSE_LLINE=137, LSE_RLINE=143 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(57[10] 91[8])
    defparam count__i15.GSR = "ENABLED";
    CCU2D add_1019_31 (.A0(d3[64]), .B0(n5102), .C0(n5103[28]), .D0(d2[64]), 
          .A1(d3[65]), .B1(n5102), .C1(n5103[29]), .D1(d2[65]), .CIN(n11846), 
          .COUT(n11847), .S0(d3_71__N_561[64]), .S1(d3_71__N_561[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1019_31.INIT0 = 16'h74b8;
    defparam add_1019_31.INIT1 = 16'h74b8;
    defparam add_1019_31.INJECT1_0 = "NO";
    defparam add_1019_31.INJECT1_1 = "NO";
    CCU2D add_1019_35 (.A0(d3[68]), .B0(n5102), .C0(n5103[32]), .D0(d2[68]), 
          .A1(d3[69]), .B1(n5102), .C1(n5103[33]), .D1(d2[69]), .CIN(n11848), 
          .COUT(n11849), .S0(d3_71__N_561[68]), .S1(d3_71__N_561[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1019_35.INIT0 = 16'h74b8;
    defparam add_1019_35.INIT1 = 16'h74b8;
    defparam add_1019_35.INJECT1_0 = "NO";
    defparam add_1019_35.INJECT1_1 = "NO";
    CCU2D add_1018_2 (.A0(d2[36]), .B0(d3[36]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[37]), .B1(d3[37]), .C1(GND_net), .D1(GND_net), .COUT(n11852), 
          .S1(n5103[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1018_2.INIT0 = 16'h7000;
    defparam add_1018_2.INIT1 = 16'h5666;
    defparam add_1018_2.INJECT1_0 = "NO";
    defparam add_1018_2.INJECT1_1 = "NO";
    CCU2D add_1018_34 (.A0(d2[68]), .B0(d3[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[69]), .B1(d3[69]), .C1(GND_net), .D1(GND_net), .CIN(n11867), 
          .COUT(n11868), .S0(n5103[32]), .S1(n5103[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1018_34.INIT0 = 16'h5666;
    defparam add_1018_34.INIT1 = 16'h5666;
    defparam add_1018_34.INJECT1_0 = "NO";
    defparam add_1018_34.INJECT1_1 = "NO";
    CCU2D add_1018_36 (.A0(d2[70]), .B0(d3[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[71]), .B1(d3[71]), .C1(GND_net), .D1(GND_net), .CIN(n11868), 
          .S0(n5103[34]), .S1(n5103[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1018_36.INIT0 = 16'h5666;
    defparam add_1018_36.INIT1 = 16'h5666;
    defparam add_1018_36.INJECT1_0 = "NO";
    defparam add_1018_36.INJECT1_1 = "NO";
    CCU2D add_1018_30 (.A0(d2[64]), .B0(d3[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[65]), .B1(d3[65]), .C1(GND_net), .D1(GND_net), .CIN(n11865), 
          .COUT(n11866), .S0(n5103[28]), .S1(n5103[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1018_30.INIT0 = 16'h5666;
    defparam add_1018_30.INIT1 = 16'h5666;
    defparam add_1018_30.INJECT1_0 = "NO";
    defparam add_1018_30.INJECT1_1 = "NO";
    CCU2D add_1018_32 (.A0(d2[66]), .B0(d3[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[67]), .B1(d3[67]), .C1(GND_net), .D1(GND_net), .CIN(n11866), 
          .COUT(n11867), .S0(n5103[30]), .S1(n5103[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1018_32.INIT0 = 16'h5666;
    defparam add_1018_32.INIT1 = 16'h5666;
    defparam add_1018_32.INJECT1_0 = "NO";
    defparam add_1018_32.INJECT1_1 = "NO";
    CCU2D add_1018_26 (.A0(d2[60]), .B0(d3[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[61]), .B1(d3[61]), .C1(GND_net), .D1(GND_net), .CIN(n11863), 
          .COUT(n11864), .S0(n5103[24]), .S1(n5103[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1018_26.INIT0 = 16'h5666;
    defparam add_1018_26.INIT1 = 16'h5666;
    defparam add_1018_26.INJECT1_0 = "NO";
    defparam add_1018_26.INJECT1_1 = "NO";
    CCU2D add_1018_28 (.A0(d2[62]), .B0(d3[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[63]), .B1(d3[63]), .C1(GND_net), .D1(GND_net), .CIN(n11864), 
          .COUT(n11865), .S0(n5103[26]), .S1(n5103[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1018_28.INIT0 = 16'h5666;
    defparam add_1018_28.INIT1 = 16'h5666;
    defparam add_1018_28.INJECT1_0 = "NO";
    defparam add_1018_28.INJECT1_1 = "NO";
    CCU2D add_1018_22 (.A0(d2[56]), .B0(d3[56]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[57]), .B1(d3[57]), .C1(GND_net), .D1(GND_net), .CIN(n11861), 
          .COUT(n11862), .S0(n5103[20]), .S1(n5103[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1018_22.INIT0 = 16'h5666;
    defparam add_1018_22.INIT1 = 16'h5666;
    defparam add_1018_22.INJECT1_0 = "NO";
    defparam add_1018_22.INJECT1_1 = "NO";
    CCU2D add_1018_24 (.A0(d2[58]), .B0(d3[58]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[59]), .B1(d3[59]), .C1(GND_net), .D1(GND_net), .CIN(n11862), 
          .COUT(n11863), .S0(n5103[22]), .S1(n5103[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1018_24.INIT0 = 16'h5666;
    defparam add_1018_24.INIT1 = 16'h5666;
    defparam add_1018_24.INJECT1_0 = "NO";
    defparam add_1018_24.INJECT1_1 = "NO";
    CCU2D add_1018_18 (.A0(d2[52]), .B0(d3[52]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[53]), .B1(d3[53]), .C1(GND_net), .D1(GND_net), .CIN(n11859), 
          .COUT(n11860), .S0(n5103[16]), .S1(n5103[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1018_18.INIT0 = 16'h5666;
    defparam add_1018_18.INIT1 = 16'h5666;
    defparam add_1018_18.INJECT1_0 = "NO";
    defparam add_1018_18.INJECT1_1 = "NO";
    CCU2D add_1018_20 (.A0(d2[54]), .B0(d3[54]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[55]), .B1(d3[55]), .C1(GND_net), .D1(GND_net), .CIN(n11860), 
          .COUT(n11861), .S0(n5103[18]), .S1(n5103[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1018_20.INIT0 = 16'h5666;
    defparam add_1018_20.INIT1 = 16'h5666;
    defparam add_1018_20.INJECT1_0 = "NO";
    defparam add_1018_20.INJECT1_1 = "NO";
    CCU2D add_1018_14 (.A0(d2[48]), .B0(d3[48]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[49]), .B1(d3[49]), .C1(GND_net), .D1(GND_net), .CIN(n11857), 
          .COUT(n11858), .S0(n5103[12]), .S1(n5103[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1018_14.INIT0 = 16'h5666;
    defparam add_1018_14.INIT1 = 16'h5666;
    defparam add_1018_14.INJECT1_0 = "NO";
    defparam add_1018_14.INJECT1_1 = "NO";
    CCU2D add_1018_16 (.A0(d2[50]), .B0(d3[50]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[51]), .B1(d3[51]), .C1(GND_net), .D1(GND_net), .CIN(n11858), 
          .COUT(n11859), .S0(n5103[14]), .S1(n5103[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1018_16.INIT0 = 16'h5666;
    defparam add_1018_16.INIT1 = 16'h5666;
    defparam add_1018_16.INJECT1_0 = "NO";
    defparam add_1018_16.INJECT1_1 = "NO";
    CCU2D add_1018_10 (.A0(d2[44]), .B0(d3[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[45]), .B1(d3[45]), .C1(GND_net), .D1(GND_net), .CIN(n11855), 
          .COUT(n11856), .S0(n5103[8]), .S1(n5103[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1018_10.INIT0 = 16'h5666;
    defparam add_1018_10.INIT1 = 16'h5666;
    defparam add_1018_10.INJECT1_0 = "NO";
    defparam add_1018_10.INJECT1_1 = "NO";
    CCU2D add_1018_12 (.A0(d2[46]), .B0(d3[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[47]), .B1(d3[47]), .C1(GND_net), .D1(GND_net), .CIN(n11856), 
          .COUT(n11857), .S0(n5103[10]), .S1(n5103[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1018_12.INIT0 = 16'h5666;
    defparam add_1018_12.INIT1 = 16'h5666;
    defparam add_1018_12.INJECT1_0 = "NO";
    defparam add_1018_12.INJECT1_1 = "NO";
    CCU2D add_1018_8 (.A0(d2[42]), .B0(d3[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[43]), .B1(d3[43]), .C1(GND_net), .D1(GND_net), .CIN(n11854), 
          .COUT(n11855), .S0(n5103[6]), .S1(n5103[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1018_8.INIT0 = 16'h5666;
    defparam add_1018_8.INIT1 = 16'h5666;
    defparam add_1018_8.INJECT1_0 = "NO";
    defparam add_1018_8.INJECT1_1 = "NO";
    CCU2D add_1013_12 (.A0(d1[46]), .B0(d2[46]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[47]), .B1(d2[47]), .C1(GND_net), .D1(GND_net), .CIN(n11897), 
          .COUT(n11898), .S0(n4951[10]), .S1(n4951[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1013_12.INIT0 = 16'h5666;
    defparam add_1013_12.INIT1 = 16'h5666;
    defparam add_1013_12.INJECT1_0 = "NO";
    defparam add_1013_12.INJECT1_1 = "NO";
    CCU2D add_1009_9 (.A0(d1[42]), .B0(n4798), .C0(n4799[6]), .D0(MixerOutCos[11]), 
          .A1(d1[43]), .B1(n4798), .C1(n4799[7]), .D1(MixerOutCos[11]), 
          .CIN(n11917), .COUT(n11918), .S0(d1_71__N_417[42]), .S1(d1_71__N_417[43]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1009_9.INIT0 = 16'h74b8;
    defparam add_1009_9.INIT1 = 16'h74b8;
    defparam add_1009_9.INJECT1_0 = "NO";
    defparam add_1009_9.INJECT1_1 = "NO";
    CCU2D add_1008_36 (.A0(MixerOutCos[11]), .B0(d1[70]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[71]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11950), .S0(n4799[34]), .S1(n4799[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1008_36.INIT0 = 16'h5666;
    defparam add_1008_36.INIT1 = 16'h5666;
    defparam add_1008_36.INJECT1_0 = "NO";
    defparam add_1008_36.INJECT1_1 = "NO";
    CCU2D add_1008_34 (.A0(MixerOutCos[11]), .B0(d1[68]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[69]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11949), .COUT(n11950), .S0(n4799[32]), 
          .S1(n4799[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1008_34.INIT0 = 16'h5666;
    defparam add_1008_34.INIT1 = 16'h5666;
    defparam add_1008_34.INJECT1_0 = "NO";
    defparam add_1008_34.INJECT1_1 = "NO";
    LUT4 i4797_2_lut (.A(d2[36]), .B(d3[36]), .Z(n5103[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4797_2_lut.init = 16'h6666;
    CCU2D add_1008_32 (.A0(MixerOutCos[11]), .B0(d1[66]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[67]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11948), .COUT(n11949), .S0(n4799[30]), 
          .S1(n4799[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1008_32.INIT0 = 16'h5666;
    defparam add_1008_32.INIT1 = 16'h5666;
    defparam add_1008_32.INJECT1_0 = "NO";
    defparam add_1008_32.INJECT1_1 = "NO";
    CCU2D add_1008_30 (.A0(MixerOutCos[11]), .B0(d1[64]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[65]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11947), .COUT(n11948), .S0(n4799[28]), 
          .S1(n4799[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1008_30.INIT0 = 16'h5666;
    defparam add_1008_30.INIT1 = 16'h5666;
    defparam add_1008_30.INJECT1_0 = "NO";
    defparam add_1008_30.INJECT1_1 = "NO";
    CCU2D add_1009_7 (.A0(d1[40]), .B0(n4798), .C0(n4799[4]), .D0(MixerOutCos[11]), 
          .A1(d1[41]), .B1(n4798), .C1(n4799[5]), .D1(MixerOutCos[11]), 
          .CIN(n11916), .COUT(n11917), .S0(d1_71__N_417[40]), .S1(d1_71__N_417[41]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1009_7.INIT0 = 16'h74b8;
    defparam add_1009_7.INIT1 = 16'h74b8;
    defparam add_1009_7.INJECT1_0 = "NO";
    defparam add_1009_7.INJECT1_1 = "NO";
    CCU2D add_1008_28 (.A0(MixerOutCos[11]), .B0(d1[62]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[63]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11946), .COUT(n11947), .S0(n4799[26]), 
          .S1(n4799[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1008_28.INIT0 = 16'h5666;
    defparam add_1008_28.INIT1 = 16'h5666;
    defparam add_1008_28.INJECT1_0 = "NO";
    defparam add_1008_28.INJECT1_1 = "NO";
    CCU2D add_1009_5 (.A0(d1[38]), .B0(n4798), .C0(n4799[2]), .D0(MixerOutCos[11]), 
          .A1(d1[39]), .B1(n4798), .C1(n4799[3]), .D1(MixerOutCos[11]), 
          .CIN(n11915), .COUT(n11916), .S0(d1_71__N_417[38]), .S1(d1_71__N_417[39]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1009_5.INIT0 = 16'h74b8;
    defparam add_1009_5.INIT1 = 16'h74b8;
    defparam add_1009_5.INJECT1_0 = "NO";
    defparam add_1009_5.INJECT1_1 = "NO";
    CCU2D add_1008_26 (.A0(MixerOutCos[11]), .B0(d1[60]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[61]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11945), .COUT(n11946), .S0(n4799[24]), 
          .S1(n4799[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1008_26.INIT0 = 16'h5666;
    defparam add_1008_26.INIT1 = 16'h5666;
    defparam add_1008_26.INJECT1_0 = "NO";
    defparam add_1008_26.INJECT1_1 = "NO";
    CCU2D add_1008_24 (.A0(MixerOutCos[11]), .B0(d1[58]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[59]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11944), .COUT(n11945), .S0(n4799[22]), 
          .S1(n4799[23]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1008_24.INIT0 = 16'h5666;
    defparam add_1008_24.INIT1 = 16'h5666;
    defparam add_1008_24.INJECT1_0 = "NO";
    defparam add_1008_24.INJECT1_1 = "NO";
    CCU2D add_1008_22 (.A0(MixerOutCos[11]), .B0(d1[56]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[57]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11943), .COUT(n11944), .S0(n4799[20]), 
          .S1(n4799[21]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1008_22.INIT0 = 16'h5666;
    defparam add_1008_22.INIT1 = 16'h5666;
    defparam add_1008_22.INJECT1_0 = "NO";
    defparam add_1008_22.INJECT1_1 = "NO";
    CCU2D add_1009_3 (.A0(d1[36]), .B0(n4798), .C0(n4799[0]), .D0(MixerOutCos[11]), 
          .A1(d1[37]), .B1(n4798), .C1(n4799[1]), .D1(MixerOutCos[11]), 
          .CIN(n11914), .COUT(n11915), .S0(d1_71__N_417[36]), .S1(d1_71__N_417[37]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1009_3.INIT0 = 16'h74b8;
    defparam add_1009_3.INIT1 = 16'h74b8;
    defparam add_1009_3.INJECT1_0 = "NO";
    defparam add_1009_3.INJECT1_1 = "NO";
    CCU2D add_1008_20 (.A0(MixerOutCos[11]), .B0(d1[54]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[55]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11942), .COUT(n11943), .S0(n4799[18]), 
          .S1(n4799[19]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1008_20.INIT0 = 16'h5666;
    defparam add_1008_20.INIT1 = 16'h5666;
    defparam add_1008_20.INJECT1_0 = "NO";
    defparam add_1008_20.INJECT1_1 = "NO";
    CCU2D add_1008_18 (.A0(MixerOutCos[11]), .B0(d1[52]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[53]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11941), .COUT(n11942), .S0(n4799[16]), 
          .S1(n4799[17]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1008_18.INIT0 = 16'h5666;
    defparam add_1008_18.INIT1 = 16'h5666;
    defparam add_1008_18.INJECT1_0 = "NO";
    defparam add_1008_18.INJECT1_1 = "NO";
    CCU2D add_1008_16 (.A0(MixerOutCos[11]), .B0(d1[50]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[51]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11940), .COUT(n11941), .S0(n4799[14]), 
          .S1(n4799[15]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1008_16.INIT0 = 16'h5666;
    defparam add_1008_16.INIT1 = 16'h5666;
    defparam add_1008_16.INJECT1_0 = "NO";
    defparam add_1008_16.INJECT1_1 = "NO";
    CCU2D add_1008_14 (.A0(MixerOutCos[11]), .B0(d1[48]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[49]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11939), .COUT(n11940), .S0(n4799[12]), 
          .S1(n4799[13]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1008_14.INIT0 = 16'h5666;
    defparam add_1008_14.INIT1 = 16'h5666;
    defparam add_1008_14.INJECT1_0 = "NO";
    defparam add_1008_14.INJECT1_1 = "NO";
    CCU2D add_1008_12 (.A0(MixerOutCos[11]), .B0(d1[46]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[47]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11938), .COUT(n11939), .S0(n4799[10]), 
          .S1(n4799[11]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1008_12.INIT0 = 16'h5666;
    defparam add_1008_12.INIT1 = 16'h5666;
    defparam add_1008_12.INJECT1_0 = "NO";
    defparam add_1008_12.INJECT1_1 = "NO";
    CCU2D add_1008_10 (.A0(MixerOutCos[11]), .B0(d1[44]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[45]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11937), .COUT(n11938), .S0(n4799[8]), 
          .S1(n4799[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1008_10.INIT0 = 16'h5666;
    defparam add_1008_10.INIT1 = 16'h5666;
    defparam add_1008_10.INJECT1_0 = "NO";
    defparam add_1008_10.INJECT1_1 = "NO";
    CCU2D add_1008_8 (.A0(MixerOutCos[11]), .B0(d1[42]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[43]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11936), .COUT(n11937), .S0(n4799[6]), 
          .S1(n4799[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1008_8.INIT0 = 16'h5666;
    defparam add_1008_8.INIT1 = 16'h5666;
    defparam add_1008_8.INJECT1_0 = "NO";
    defparam add_1008_8.INJECT1_1 = "NO";
    CCU2D add_1008_6 (.A0(MixerOutCos[11]), .B0(d1[40]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[41]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11935), .COUT(n11936), .S0(n4799[4]), 
          .S1(n4799[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1008_6.INIT0 = 16'h5666;
    defparam add_1008_6.INIT1 = 16'h5666;
    defparam add_1008_6.INJECT1_0 = "NO";
    defparam add_1008_6.INJECT1_1 = "NO";
    CCU2D add_1008_4 (.A0(MixerOutCos[11]), .B0(d1[38]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[39]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11934), .COUT(n11935), .S0(n4799[2]), 
          .S1(n4799[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1008_4.INIT0 = 16'h5666;
    defparam add_1008_4.INIT1 = 16'h5666;
    defparam add_1008_4.INJECT1_0 = "NO";
    defparam add_1008_4.INJECT1_1 = "NO";
    CCU2D add_1013_10 (.A0(d1[44]), .B0(d2[44]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[45]), .B1(d2[45]), .C1(GND_net), .D1(GND_net), .CIN(n11896), 
          .COUT(n11897), .S0(n4951[8]), .S1(n4951[9]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1013_10.INIT0 = 16'h5666;
    defparam add_1013_10.INIT1 = 16'h5666;
    defparam add_1013_10.INJECT1_0 = "NO";
    defparam add_1013_10.INJECT1_1 = "NO";
    CCU2D add_1008_2 (.A0(MixerOutCos[11]), .B0(d1[36]), .C0(GND_net), 
          .D0(GND_net), .A1(MixerOutCos[11]), .B1(d1[37]), .C1(GND_net), 
          .D1(GND_net), .COUT(n11934), .S1(n4799[1]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1008_2.INIT0 = 16'h7000;
    defparam add_1008_2.INIT1 = 16'h5666;
    defparam add_1008_2.INJECT1_0 = "NO";
    defparam add_1008_2.INJECT1_1 = "NO";
    CCU2D add_1009_37 (.A0(d1[70]), .B0(n4798), .C0(n4799[34]), .D0(MixerOutCos[11]), 
          .A1(d1[71]), .B1(n4798), .C1(n4799[35]), .D1(MixerOutCos[11]), 
          .CIN(n11931), .S0(d1_71__N_417[70]), .S1(d1_71__N_417[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1009_37.INIT0 = 16'h74b8;
    defparam add_1009_37.INIT1 = 16'h74b8;
    defparam add_1009_37.INJECT1_0 = "NO";
    defparam add_1009_37.INJECT1_1 = "NO";
    CCU2D add_1013_8 (.A0(d1[42]), .B0(d2[42]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[43]), .B1(d2[43]), .C1(GND_net), .D1(GND_net), .CIN(n11895), 
          .COUT(n11896), .S0(n4951[6]), .S1(n4951[7]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1013_8.INIT0 = 16'h5666;
    defparam add_1013_8.INIT1 = 16'h5666;
    defparam add_1013_8.INJECT1_0 = "NO";
    defparam add_1013_8.INJECT1_1 = "NO";
    CCU2D add_1009_35 (.A0(d1[68]), .B0(n4798), .C0(n4799[32]), .D0(MixerOutCos[11]), 
          .A1(d1[69]), .B1(n4798), .C1(n4799[33]), .D1(MixerOutCos[11]), 
          .CIN(n11930), .COUT(n11931), .S0(d1_71__N_417[68]), .S1(d1_71__N_417[69]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1009_35.INIT0 = 16'h74b8;
    defparam add_1009_35.INIT1 = 16'h74b8;
    defparam add_1009_35.INJECT1_0 = "NO";
    defparam add_1009_35.INJECT1_1 = "NO";
    CCU2D add_1009_33 (.A0(d1[66]), .B0(n4798), .C0(n4799[30]), .D0(MixerOutCos[11]), 
          .A1(d1[67]), .B1(n4798), .C1(n4799[31]), .D1(MixerOutCos[11]), 
          .CIN(n11929), .COUT(n11930), .S0(d1_71__N_417[66]), .S1(d1_71__N_417[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1009_33.INIT0 = 16'h74b8;
    defparam add_1009_33.INIT1 = 16'h74b8;
    defparam add_1009_33.INJECT1_0 = "NO";
    defparam add_1009_33.INJECT1_1 = "NO";
    CCU2D add_1009_31 (.A0(d1[64]), .B0(n4798), .C0(n4799[28]), .D0(MixerOutCos[11]), 
          .A1(d1[65]), .B1(n4798), .C1(n4799[29]), .D1(MixerOutCos[11]), 
          .CIN(n11928), .COUT(n11929), .S0(d1_71__N_417[64]), .S1(d1_71__N_417[65]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1009_31.INIT0 = 16'h74b8;
    defparam add_1009_31.INIT1 = 16'h74b8;
    defparam add_1009_31.INJECT1_0 = "NO";
    defparam add_1009_31.INJECT1_1 = "NO";
    CCU2D add_1009_29 (.A0(d1[62]), .B0(n4798), .C0(n4799[26]), .D0(MixerOutCos[11]), 
          .A1(d1[63]), .B1(n4798), .C1(n4799[27]), .D1(MixerOutCos[11]), 
          .CIN(n11927), .COUT(n11928), .S0(d1_71__N_417[62]), .S1(d1_71__N_417[63]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1009_29.INIT0 = 16'h74b8;
    defparam add_1009_29.INIT1 = 16'h74b8;
    defparam add_1009_29.INJECT1_0 = "NO";
    defparam add_1009_29.INJECT1_1 = "NO";
    CCU2D add_1009_27 (.A0(d1[60]), .B0(n4798), .C0(n4799[24]), .D0(MixerOutCos[11]), 
          .A1(d1[61]), .B1(n4798), .C1(n4799[25]), .D1(MixerOutCos[11]), 
          .CIN(n11926), .COUT(n11927), .S0(d1_71__N_417[60]), .S1(d1_71__N_417[61]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1009_27.INIT0 = 16'h74b8;
    defparam add_1009_27.INIT1 = 16'h74b8;
    defparam add_1009_27.INJECT1_0 = "NO";
    defparam add_1009_27.INJECT1_1 = "NO";
    CCU2D add_1009_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n4798), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n11914));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1009_1.INIT0 = 16'hF000;
    defparam add_1009_1.INIT1 = 16'h0555;
    defparam add_1009_1.INJECT1_0 = "NO";
    defparam add_1009_1.INJECT1_1 = "NO";
    CCU2D add_1009_25 (.A0(d1[58]), .B0(n4798), .C0(n4799[22]), .D0(MixerOutCos[11]), 
          .A1(d1[59]), .B1(n4798), .C1(n4799[23]), .D1(MixerOutCos[11]), 
          .CIN(n11925), .COUT(n11926), .S0(d1_71__N_417[58]), .S1(d1_71__N_417[59]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1009_25.INIT0 = 16'h74b8;
    defparam add_1009_25.INIT1 = 16'h74b8;
    defparam add_1009_25.INJECT1_0 = "NO";
    defparam add_1009_25.INJECT1_1 = "NO";
    CCU2D add_1009_23 (.A0(d1[56]), .B0(n4798), .C0(n4799[20]), .D0(MixerOutCos[11]), 
          .A1(d1[57]), .B1(n4798), .C1(n4799[21]), .D1(MixerOutCos[11]), 
          .CIN(n11924), .COUT(n11925), .S0(d1_71__N_417[56]), .S1(d1_71__N_417[57]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1009_23.INIT0 = 16'h74b8;
    defparam add_1009_23.INIT1 = 16'h74b8;
    defparam add_1009_23.INJECT1_0 = "NO";
    defparam add_1009_23.INJECT1_1 = "NO";
    CCU2D add_1018_6 (.A0(d2[40]), .B0(d3[40]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[41]), .B1(d3[41]), .C1(GND_net), .D1(GND_net), .CIN(n11853), 
          .COUT(n11854), .S0(n5103[4]), .S1(n5103[5]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1018_6.INIT0 = 16'h5666;
    defparam add_1018_6.INIT1 = 16'h5666;
    defparam add_1018_6.INJECT1_0 = "NO";
    defparam add_1018_6.INJECT1_1 = "NO";
    CCU2D add_1013_36 (.A0(d1[70]), .B0(d2[70]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[71]), .B1(d2[71]), .C1(GND_net), .D1(GND_net), .CIN(n11909), 
          .S0(n4951[34]), .S1(n4951[35]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1013_36.INIT0 = 16'h5666;
    defparam add_1013_36.INIT1 = 16'h5666;
    defparam add_1013_36.INJECT1_0 = "NO";
    defparam add_1013_36.INJECT1_1 = "NO";
    CCU2D add_1009_21 (.A0(d1[54]), .B0(n4798), .C0(n4799[18]), .D0(MixerOutCos[11]), 
          .A1(d1[55]), .B1(n4798), .C1(n4799[19]), .D1(MixerOutCos[11]), 
          .CIN(n11923), .COUT(n11924), .S0(d1_71__N_417[54]), .S1(d1_71__N_417[55]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1009_21.INIT0 = 16'h74b8;
    defparam add_1009_21.INIT1 = 16'h74b8;
    defparam add_1009_21.INJECT1_0 = "NO";
    defparam add_1009_21.INJECT1_1 = "NO";
    CCU2D add_1013_34 (.A0(d1[68]), .B0(d2[68]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[69]), .B1(d2[69]), .C1(GND_net), .D1(GND_net), .CIN(n11908), 
          .COUT(n11909), .S0(n4951[32]), .S1(n4951[33]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1013_34.INIT0 = 16'h5666;
    defparam add_1013_34.INIT1 = 16'h5666;
    defparam add_1013_34.INJECT1_0 = "NO";
    defparam add_1013_34.INJECT1_1 = "NO";
    CCU2D add_1009_19 (.A0(d1[52]), .B0(n4798), .C0(n4799[16]), .D0(MixerOutCos[11]), 
          .A1(d1[53]), .B1(n4798), .C1(n4799[17]), .D1(MixerOutCos[11]), 
          .CIN(n11922), .COUT(n11923), .S0(d1_71__N_417[52]), .S1(d1_71__N_417[53]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1009_19.INIT0 = 16'h74b8;
    defparam add_1009_19.INIT1 = 16'h74b8;
    defparam add_1009_19.INJECT1_0 = "NO";
    defparam add_1009_19.INJECT1_1 = "NO";
    CCU2D add_1013_32 (.A0(d1[66]), .B0(d2[66]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[67]), .B1(d2[67]), .C1(GND_net), .D1(GND_net), .CIN(n11907), 
          .COUT(n11908), .S0(n4951[30]), .S1(n4951[31]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1013_32.INIT0 = 16'h5666;
    defparam add_1013_32.INIT1 = 16'h5666;
    defparam add_1013_32.INJECT1_0 = "NO";
    defparam add_1013_32.INJECT1_1 = "NO";
    CCU2D add_1009_17 (.A0(d1[50]), .B0(n4798), .C0(n4799[14]), .D0(MixerOutCos[11]), 
          .A1(d1[51]), .B1(n4798), .C1(n4799[15]), .D1(MixerOutCos[11]), 
          .CIN(n11921), .COUT(n11922), .S0(d1_71__N_417[50]), .S1(d1_71__N_417[51]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1009_17.INIT0 = 16'h74b8;
    defparam add_1009_17.INIT1 = 16'h74b8;
    defparam add_1009_17.INJECT1_0 = "NO";
    defparam add_1009_17.INJECT1_1 = "NO";
    CCU2D add_1013_30 (.A0(d1[64]), .B0(d2[64]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[65]), .B1(d2[65]), .C1(GND_net), .D1(GND_net), .CIN(n11906), 
          .COUT(n11907), .S0(n4951[28]), .S1(n4951[29]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1013_30.INIT0 = 16'h5666;
    defparam add_1013_30.INIT1 = 16'h5666;
    defparam add_1013_30.INJECT1_0 = "NO";
    defparam add_1013_30.INJECT1_1 = "NO";
    CCU2D add_1009_15 (.A0(d1[48]), .B0(n4798), .C0(n4799[12]), .D0(MixerOutCos[11]), 
          .A1(d1[49]), .B1(n4798), .C1(n4799[13]), .D1(MixerOutCos[11]), 
          .CIN(n11920), .COUT(n11921), .S0(d1_71__N_417[48]), .S1(d1_71__N_417[49]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1009_15.INIT0 = 16'h74b8;
    defparam add_1009_15.INIT1 = 16'h74b8;
    defparam add_1009_15.INJECT1_0 = "NO";
    defparam add_1009_15.INJECT1_1 = "NO";
    CCU2D add_1013_28 (.A0(d1[62]), .B0(d2[62]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[63]), .B1(d2[63]), .C1(GND_net), .D1(GND_net), .CIN(n11905), 
          .COUT(n11906), .S0(n4951[26]), .S1(n4951[27]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1013_28.INIT0 = 16'h5666;
    defparam add_1013_28.INIT1 = 16'h5666;
    defparam add_1013_28.INJECT1_0 = "NO";
    defparam add_1013_28.INJECT1_1 = "NO";
    CCU2D add_1009_13 (.A0(d1[46]), .B0(n4798), .C0(n4799[10]), .D0(MixerOutCos[11]), 
          .A1(d1[47]), .B1(n4798), .C1(n4799[11]), .D1(MixerOutCos[11]), 
          .CIN(n11919), .COUT(n11920), .S0(d1_71__N_417[46]), .S1(d1_71__N_417[47]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1009_13.INIT0 = 16'h74b8;
    defparam add_1009_13.INIT1 = 16'h74b8;
    defparam add_1009_13.INJECT1_0 = "NO";
    defparam add_1009_13.INJECT1_1 = "NO";
    CCU2D add_1013_26 (.A0(d1[60]), .B0(d2[60]), .C0(GND_net), .D0(GND_net), 
          .A1(d1[61]), .B1(d2[61]), .C1(GND_net), .D1(GND_net), .CIN(n11904), 
          .COUT(n11905), .S0(n4951[24]), .S1(n4951[25]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(64[13:20])
    defparam add_1013_26.INIT0 = 16'h5666;
    defparam add_1013_26.INIT1 = 16'h5666;
    defparam add_1013_26.INJECT1_0 = "NO";
    defparam add_1013_26.INJECT1_1 = "NO";
    CCU2D add_1009_11 (.A0(d1[44]), .B0(n4798), .C0(n4799[8]), .D0(MixerOutCos[11]), 
          .A1(d1[45]), .B1(n4798), .C1(n4799[9]), .D1(MixerOutCos[11]), 
          .CIN(n11918), .COUT(n11919), .S0(d1_71__N_417[44]), .S1(d1_71__N_417[45]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(62[13:22])
    defparam add_1009_11.INIT0 = 16'h74b8;
    defparam add_1009_11.INIT1 = 16'h74b8;
    defparam add_1009_11.INJECT1_0 = "NO";
    defparam add_1009_11.INJECT1_1 = "NO";
    CCU2D add_1018_4 (.A0(d2[38]), .B0(d3[38]), .C0(GND_net), .D0(GND_net), 
          .A1(d2[39]), .B1(d3[39]), .C1(GND_net), .D1(GND_net), .CIN(n11852), 
          .COUT(n11853), .S0(n5103[2]), .S1(n5103[3]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1018_4.INIT0 = 16'h5666;
    defparam add_1018_4.INIT1 = 16'h5666;
    defparam add_1018_4.INJECT1_0 = "NO";
    defparam add_1018_4.INJECT1_1 = "NO";
    CCU2D add_1019_37 (.A0(d3[70]), .B0(n5102), .C0(n5103[34]), .D0(d2[70]), 
          .A1(d3[71]), .B1(n5102), .C1(n5103[35]), .D1(d2[71]), .CIN(n11849), 
          .S0(d3_71__N_561[70]), .S1(d3_71__N_561[71]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1019_37.INIT0 = 16'h74b8;
    defparam add_1019_37.INIT1 = 16'h74b8;
    defparam add_1019_37.INJECT1_0 = "NO";
    defparam add_1019_37.INJECT1_1 = "NO";
    CCU2D add_1019_33 (.A0(d3[66]), .B0(n5102), .C0(n5103[30]), .D0(d2[66]), 
          .A1(d3[67]), .B1(n5102), .C1(n5103[31]), .D1(d2[67]), .CIN(n11847), 
          .COUT(n11848), .S0(d3_71__N_561[66]), .S1(d3_71__N_561[67]));   // c:/users/user/lattice/1bitadcfpgasdr/cic.v(66[13:20])
    defparam add_1019_33.INIT0 = 16'h74b8;
    defparam add_1019_33.INIT1 = 16'h74b8;
    defparam add_1019_33.INJECT1_0 = "NO";
    defparam add_1019_33.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \uart_rx(CLKS_PER_BIT=87) 
//

module \uart_rx(CLKS_PER_BIT=87)  (\UartClk[2] , osc_clk, i_Rx_Serial_c, 
            o_Rx_DV_c_0, o_Rx_Byte_c_0, n7319, o_Rx_Byte_c_2, o_Rx_Byte_c_3, 
            o_Rx_Byte_c_4, o_Rx_Byte_c_5, o_Rx_Byte_c_6, o_Rx_Byte_c_7, 
            GND_net) /* synthesis syn_module_defined=1 */ ;
    input \UartClk[2] ;
    input osc_clk;
    input i_Rx_Serial_c;
    output o_Rx_DV_c_0;
    output o_Rx_Byte_c_0;
    output n7319;
    output o_Rx_Byte_c_2;
    output o_Rx_Byte_c_3;
    output o_Rx_Byte_c_4;
    output o_Rx_Byte_c_5;
    output o_Rx_Byte_c_6;
    output o_Rx_Byte_c_7;
    input GND_net;
    
    wire \UartClk[2]  /* synthesis SET_AS_NETWORK=\uart_tx1/UartClk[2], is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uarttx.v(37[14:21])
    wire osc_clk /* synthesis SET_AS_NETWORK=osc_clk, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(55[8:15])
    wire [15:0]r_Clock_Count;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(39[18:31])
    
    wire UartClk_2_enable_56, n8362;
    wire [15:0]n69;
    wire [2:0]r_Bit_Index;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(40[17:28])
    
    wire n12914, n13769;
    wire [2:0]r_SM_Main;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(43[17:26])
    
    wire n13545, r_Rx_DV_last, r_Rx_DV, r_Rx_Data_R, r_Rx_Data, n12362, 
        n13756, n8365, r_Rx_DV_last_N_2482, r_Rx_DV_N_2483;
    wire [7:0]r_Rx_Byte;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(41[17:26])
    
    wire UartClk_2_enable_10, n13030, n13872, n13050, UartClk_2_enable_11, 
        n13750, UartClk_2_enable_22, UartClk_2_enable_52, UartClk_2_enable_13, 
        UartClk_2_enable_15, UartClk_2_enable_17, UartClk_2_enable_18;
    wire [2:0]r_SM_Main_2__N_2417;
    
    wire n13754, n13782, n13760, UartClk_2_enable_21, UartClk_2_enable_29, 
        n12904, n13870, n8940, n13543, n13781, n13780, n13179, 
        n24, n13544, n12870, n13187, n11624, n11623, n11622, n11621, 
        n11620, n11619, n11618, n11617, n8998, n13171, n13163, 
        n13161, n10;
    
    FD1P3IX r_Clock_Count_932__i1 (.D(n69[1]), .SP(UartClk_2_enable_56), 
            .CD(n8362), .CK(\UartClk[2] ), .Q(r_Clock_Count[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932__i1.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(r_Bit_Index[1]), .B(r_Bit_Index[0]), .Z(n12914)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(112[17:39])
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 i1_3_lut_rep_176 (.A(r_Clock_Count[3]), .B(r_Clock_Count[5]), .C(r_Clock_Count[0]), 
         .Z(n13769)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_rep_176.init = 16'h8080;
    FD1S3IX r_SM_Main_i0 (.D(n13545), .CK(\UartClk[2] ), .CD(r_SM_Main[2]), 
            .Q(r_SM_Main[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_SM_Main_i0.GSR = "ENABLED";
    FD1S3AX r_Rx_DV_last_60 (.D(r_Rx_DV), .CK(osc_clk), .Q(r_Rx_DV_last)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(47[11] 52[8])
    defparam r_Rx_DV_last_60.GSR = "ENABLED";
    FD1S3AY r_Rx_Data_R_61 (.D(i_Rx_Serial_c), .CK(\UartClk[2] ), .Q(r_Rx_Data_R)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(57[12] 61[8])
    defparam r_Rx_Data_R_61.GSR = "ENABLED";
    FD1S3AY r_Rx_Data_62 (.D(r_Rx_Data_R), .CK(\UartClk[2] ), .Q(r_Rx_Data)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(57[12] 61[8])
    defparam r_Rx_Data_62.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_163_4_lut (.A(r_Clock_Count[3]), .B(r_Clock_Count[5]), 
         .C(r_Clock_Count[0]), .D(n12362), .Z(n13756)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_2_lut_rep_163_4_lut.init = 16'hff7f;
    FD1S3IX o_Rx_DV_59 (.D(r_Rx_DV_last_N_2482), .CK(osc_clk), .CD(n8365), 
            .Q(o_Rx_DV_c_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(47[11] 52[8])
    defparam o_Rx_DV_59.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i1 (.D(r_Rx_Byte[0]), .SP(r_Rx_DV_N_2483), .CK(\UartClk[2] ), 
            .Q(o_Rx_Byte_c_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam o_Rx_Byte_i1.GSR = "ENABLED";
    FD1P3AX r_Bit_Index_i0 (.D(n13030), .SP(UartClk_2_enable_10), .CK(\UartClk[2] ), 
            .Q(r_Bit_Index[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Bit_Index_i0.GSR = "ENABLED";
    FD1P3AX r_Bit_Index_i2 (.D(n13872), .SP(UartClk_2_enable_10), .CK(\UartClk[2] ), 
            .Q(r_Bit_Index[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Bit_Index_i2.GSR = "ENABLED";
    FD1P3AX r_Bit_Index_i1 (.D(n13050), .SP(UartClk_2_enable_10), .CK(\UartClk[2] ), 
            .Q(r_Bit_Index[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Bit_Index_i1.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i7 (.D(r_Rx_Data), .SP(UartClk_2_enable_11), .CK(\UartClk[2] ), 
            .Q(r_Rx_Byte[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Rx_Byte_i7.GSR = "ENABLED";
    LUT4 i5875_2_lut_3_lut_4_lut (.A(r_Bit_Index[2]), .B(n13750), .C(r_Bit_Index[1]), 
         .D(r_Bit_Index[0]), .Z(UartClk_2_enable_22)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(112[17:39])
    defparam i5875_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i2362_1_lut (.A(r_Rx_DV), .Z(n8365)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam i2362_1_lut.init = 16'h5555;
    LUT4 r_Rx_DV_last_I_0_1_lut (.A(r_Rx_DV_last), .Z(r_Rx_DV_last_N_2482)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(50[30:43])
    defparam r_Rx_DV_last_I_0_1_lut.init = 16'h5555;
    LUT4 i5846_2_lut_3_lut_4_lut (.A(r_Bit_Index[2]), .B(n13750), .C(r_Bit_Index[1]), 
         .D(r_Bit_Index[0]), .Z(UartClk_2_enable_52)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(112[17:39])
    defparam i5846_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i5885_2_lut_3_lut_4_lut (.A(r_Bit_Index[2]), .B(n13750), .C(r_Bit_Index[1]), 
         .D(r_Bit_Index[0]), .Z(UartClk_2_enable_13)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(112[17:39])
    defparam i5885_2_lut_3_lut_4_lut.init = 16'h0020;
    FD1P3AX r_Rx_Byte_i6 (.D(r_Rx_Data), .SP(UartClk_2_enable_13), .CK(\UartClk[2] ), 
            .Q(r_Rx_Byte[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Rx_Byte_i6.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i5 (.D(r_Rx_Data), .SP(UartClk_2_enable_15), .CK(\UartClk[2] ), 
            .Q(r_Rx_Byte[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Rx_Byte_i5.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_932__i0 (.D(n69[0]), .SP(UartClk_2_enable_56), 
            .CD(n8362), .CK(\UartClk[2] ), .Q(r_Clock_Count[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932__i0.GSR = "ENABLED";
    FD1P3AX r_Rx_DV_64 (.D(r_Rx_DV_N_2483), .SP(UartClk_2_enable_17), .CK(\UartClk[2] ), 
            .Q(r_Rx_DV)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Rx_DV_64.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i4 (.D(r_Rx_Data), .SP(UartClk_2_enable_18), .CK(\UartClk[2] ), 
            .Q(r_Rx_Byte[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Rx_Byte_i4.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(r_SM_Main[0]), .B(r_SM_Main_2__N_2417[2]), .C(r_SM_Main[2]), 
         .D(r_SM_Main[1]), .Z(UartClk_2_enable_10)) /* synthesis lut_function=(!(A+(B (C)+!B (C+(D))))) */ ;
    defparam i1_4_lut.init = 16'h0405;
    LUT4 i5883_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n13754), .C(n12914), 
         .D(r_Bit_Index[2]), .Z(UartClk_2_enable_15)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(112[17:39])
    defparam i5883_2_lut_3_lut_4_lut.init = 16'h0100;
    FD1S3IX r_SM_Main_i1 (.D(n13782), .CK(\UartClk[2] ), .CD(r_SM_Main[2]), 
            .Q(r_SM_Main[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_SM_Main_i1.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i2 (.D(r_Rx_Byte[1]), .SP(r_Rx_DV_N_2483), .CK(\UartClk[2] ), 
            .Q(n7319)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam o_Rx_Byte_i2.GSR = "ENABLED";
    LUT4 i5887_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n13754), .C(n13760), 
         .D(r_Bit_Index[2]), .Z(UartClk_2_enable_11)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(112[17:39])
    defparam i5887_2_lut_3_lut_4_lut.init = 16'h1000;
    FD1P3AX r_Rx_Byte_i3 (.D(r_Rx_Data), .SP(UartClk_2_enable_21), .CK(\UartClk[2] ), 
            .Q(r_Rx_Byte[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Rx_Byte_i3.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i2 (.D(r_Rx_Data), .SP(UartClk_2_enable_22), .CK(\UartClk[2] ), 
            .Q(r_Rx_Byte[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Rx_Byte_i2.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i3 (.D(r_Rx_Byte[2]), .SP(r_Rx_DV_N_2483), .CK(\UartClk[2] ), 
            .Q(o_Rx_Byte_c_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam o_Rx_Byte_i3.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i4 (.D(r_Rx_Byte[3]), .SP(r_Rx_DV_N_2483), .CK(\UartClk[2] ), 
            .Q(o_Rx_Byte_c_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam o_Rx_Byte_i4.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i5 (.D(r_Rx_Byte[4]), .SP(r_Rx_DV_N_2483), .CK(\UartClk[2] ), 
            .Q(o_Rx_Byte_c_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam o_Rx_Byte_i5.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i6 (.D(r_Rx_Byte[5]), .SP(r_Rx_DV_N_2483), .CK(\UartClk[2] ), 
            .Q(o_Rx_Byte_c_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam o_Rx_Byte_i6.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i7 (.D(r_Rx_Byte[6]), .SP(r_Rx_DV_N_2483), .CK(\UartClk[2] ), 
            .Q(o_Rx_Byte_c_6)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam o_Rx_Byte_i7.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i8 (.D(r_Rx_Byte[7]), .SP(r_Rx_DV_N_2483), .CK(\UartClk[2] ), 
            .Q(o_Rx_Byte_c_7)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam o_Rx_Byte_i8.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i1 (.D(r_Rx_Data), .SP(UartClk_2_enable_29), .CK(\UartClk[2] ), 
            .Q(r_Rx_Byte[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Rx_Byte_i1.GSR = "ENABLED";
    FD1S3IX r_SM_Main_i2 (.D(r_SM_Main_2__N_2417[2]), .CK(\UartClk[2] ), 
            .CD(n12904), .Q(r_SM_Main[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_SM_Main_i2.GSR = "ENABLED";
    LUT4 i5873_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n13754), .C(n12914), 
         .D(r_Bit_Index[2]), .Z(UartClk_2_enable_29)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(112[17:39])
    defparam i5873_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i5877_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n13754), .C(n13760), 
         .D(r_Bit_Index[2]), .Z(UartClk_2_enable_21)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(112[17:39])
    defparam i5877_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 CIC_out_clkSin_c_bdd_2_lut_6085_3_lut (.A(n13870), .B(r_SM_Main[1]), 
         .C(r_SM_Main_2__N_2417[2]), .Z(n13872)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam CIC_out_clkSin_c_bdd_2_lut_6085_3_lut.init = 16'h8080;
    LUT4 r_SM_Main_2__N_2417_2__bdd_3_lut_5926 (.A(r_SM_Main_2__N_2417[2]), 
         .B(n8940), .C(r_SM_Main[0]), .Z(n13543)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(C))) */ ;
    defparam r_SM_Main_2__N_2417_2__bdd_3_lut_5926.init = 16'h5858;
    LUT4 i5860_3_lut_4_lut (.A(r_SM_Main_2__N_2417[2]), .B(r_SM_Main[0]), 
         .C(r_Bit_Index[0]), .D(r_SM_Main[1]), .Z(n13030)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(67[7] 159[14])
    defparam i5860_3_lut_4_lut.init = 16'h0200;
    LUT4 r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_then_4_lut (.A(r_SM_Main_2__N_2417[2]), 
         .B(r_SM_Main[1]), .C(n13756), .D(r_Rx_Data), .Z(n13781)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B+!(C+(D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(67[7] 159[14])
    defparam r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_then_4_lut.init = 16'h4447;
    LUT4 r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_else_4_lut (.A(r_SM_Main[1]), 
         .Z(n13780)) /* synthesis lut_function=(A) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(67[7] 159[14])
    defparam r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_else_4_lut.init = 16'haaaa;
    LUT4 i5904_4_lut (.A(r_SM_Main[2]), .B(r_SM_Main[1]), .C(n13756), 
         .D(n13179), .Z(UartClk_2_enable_56)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(67[7] 159[14])
    defparam i5904_4_lut.init = 16'h5455;
    LUT4 i1_2_lut_adj_25 (.A(r_Rx_Data), .B(r_SM_Main[0]), .Z(n13179)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_25.init = 16'h8888;
    LUT4 i1_4_lut_adj_26 (.A(r_SM_Main[2]), .B(n24), .C(r_SM_Main_2__N_2417[2]), 
         .D(r_SM_Main[1]), .Z(n8362)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;
    defparam i1_4_lut_adj_26.init = 16'h5044;
    LUT4 i1_4_lut_adj_27 (.A(r_Rx_Data), .B(r_SM_Main[0]), .C(n12362), 
         .D(n13769), .Z(n24)) /* synthesis lut_function=(!(A (B)+!A (B (C+!(D))))) */ ;
    defparam i1_4_lut_adj_27.init = 16'h3733;
    LUT4 i5880_2_lut_3_lut_4_lut (.A(r_Bit_Index[2]), .B(n13750), .C(r_Bit_Index[1]), 
         .D(r_Bit_Index[0]), .Z(UartClk_2_enable_18)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(112[17:39])
    defparam i5880_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 r_SM_Main_2__N_2417_2__bdd_3_lut_4_lut (.A(n13769), .B(n12362), 
         .C(r_SM_Main[0]), .D(r_Rx_Data), .Z(n13544)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D))) */ ;
    defparam r_SM_Main_2__N_2417_2__bdd_3_lut_4_lut.init = 16'hd0df;
    LUT4 i1_4_lut_adj_28 (.A(r_Clock_Count[1]), .B(n12870), .C(n13187), 
         .D(r_Clock_Count[6]), .Z(n12362)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(83[17:52])
    defparam i1_4_lut_adj_28.init = 16'hfffd;
    LUT4 i1_2_lut_adj_29 (.A(r_Clock_Count[2]), .B(r_Clock_Count[4]), .Z(n13187)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(83[17:52])
    defparam i1_2_lut_adj_29.init = 16'heeee;
    LUT4 i1103_2_lut_rep_167 (.A(r_Bit_Index[1]), .B(r_Bit_Index[0]), .Z(n13760)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(117[36:54])
    defparam i1103_2_lut_rep_167.init = 16'h8888;
    CCU2D r_Clock_Count_932_add_4_17 (.A0(r_Clock_Count[15]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11624), .S0(n69[15]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932_add_4_17.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_932_add_4_17.INIT1 = 16'h0000;
    defparam r_Clock_Count_932_add_4_17.INJECT1_0 = "NO";
    defparam r_Clock_Count_932_add_4_17.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_932_add_4_15 (.A0(r_Clock_Count[13]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[14]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n11623), .COUT(n11624), .S0(n69[13]), 
          .S1(n69[14]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932_add_4_15.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_932_add_4_15.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_932_add_4_15.INJECT1_0 = "NO";
    defparam r_Clock_Count_932_add_4_15.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_932_add_4_13 (.A0(r_Clock_Count[11]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[12]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n11622), .COUT(n11623), .S0(n69[11]), 
          .S1(n69[12]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932_add_4_13.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_932_add_4_13.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_932_add_4_13.INJECT1_0 = "NO";
    defparam r_Clock_Count_932_add_4_13.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_932_add_4_11 (.A0(r_Clock_Count[9]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[10]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n11621), .COUT(n11622), .S0(n69[9]), 
          .S1(n69[10]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932_add_4_11.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_932_add_4_11.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_932_add_4_11.INJECT1_0 = "NO";
    defparam r_Clock_Count_932_add_4_11.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_932_add_4_9 (.A0(r_Clock_Count[7]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[8]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n11620), .COUT(n11621), .S0(n69[7]), 
          .S1(n69[8]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932_add_4_9.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_932_add_4_9.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_932_add_4_9.INJECT1_0 = "NO";
    defparam r_Clock_Count_932_add_4_9.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_932_add_4_7 (.A0(r_Clock_Count[5]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[6]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n11619), .COUT(n11620), .S0(n69[5]), 
          .S1(n69[6]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932_add_4_7.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_932_add_4_7.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_932_add_4_7.INJECT1_0 = "NO";
    defparam r_Clock_Count_932_add_4_7.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_932_add_4_5 (.A0(r_Clock_Count[3]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[4]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n11618), .COUT(n11619), .S0(n69[3]), 
          .S1(n69[4]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932_add_4_5.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_932_add_4_5.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_932_add_4_5.INJECT1_0 = "NO";
    defparam r_Clock_Count_932_add_4_5.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_932_add_4_3 (.A0(r_Clock_Count[1]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(r_Clock_Count[2]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n11617), .COUT(n11618), .S0(n69[1]), 
          .S1(n69[2]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932_add_4_3.INIT0 = 16'hfaaa;
    defparam r_Clock_Count_932_add_4_3.INIT1 = 16'hfaaa;
    defparam r_Clock_Count_932_add_4_3.INJECT1_0 = "NO";
    defparam r_Clock_Count_932_add_4_3.INJECT1_1 = "NO";
    CCU2D r_Clock_Count_932_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(r_Clock_Count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n11617), .S1(n69[0]));   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932_add_4_1.INIT0 = 16'hF000;
    defparam r_Clock_Count_932_add_4_1.INIT1 = 16'h0555;
    defparam r_Clock_Count_932_add_4_1.INJECT1_0 = "NO";
    defparam r_Clock_Count_932_add_4_1.INJECT1_1 = "NO";
    LUT4 i14_4_lut_4_lut (.A(r_SM_Main[1]), .B(r_SM_Main[2]), .C(r_SM_Main[0]), 
         .D(r_SM_Main_2__N_2417[2]), .Z(UartClk_2_enable_17)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (C))) */ ;
    defparam i14_4_lut_4_lut.init = 16'h2505;
    LUT4 i5870_2_lut_3_lut (.A(r_SM_Main[1]), .B(r_SM_Main[2]), .C(r_SM_Main[0]), 
         .Z(n12904)) /* synthesis lut_function=((B+!(C))+!A) */ ;
    defparam i5870_2_lut_3_lut.init = 16'hdfdf;
    LUT4 i1_4_lut_adj_30 (.A(n8998), .B(n12870), .C(r_Clock_Count[6]), 
         .D(r_Clock_Count[5]), .Z(r_SM_Main_2__N_2417[2])) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(83[17:52])
    defparam i1_4_lut_adj_30.init = 16'hfcec;
    LUT4 i2995_4_lut (.A(r_Clock_Count[1]), .B(r_Clock_Count[4]), .C(r_Clock_Count[3]), 
         .D(r_Clock_Count[2]), .Z(n8998)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i2995_4_lut.init = 16'hc8c0;
    LUT4 i5852_2_lut_3_lut_4_lut (.A(r_SM_Main[2]), .B(r_SM_Main[1]), .C(r_SM_Main[0]), 
         .D(r_SM_Main_2__N_2417[2]), .Z(r_Rx_DV_N_2483)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i5852_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_rep_161_3_lut (.A(r_SM_Main[2]), .B(r_SM_Main[1]), .C(r_SM_Main_2__N_2417[2]), 
         .Z(n13754)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i1_2_lut_rep_161_3_lut.init = 16'hbfbf;
    LUT4 i1_4_lut_adj_31 (.A(n13171), .B(n13163), .C(n13161), .D(r_Clock_Count[11]), 
         .Z(n12870)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(83[17:52])
    defparam i1_4_lut_adj_31.init = 16'hfffe;
    LUT4 i3_4_lut (.A(r_SM_Main_2__N_2417[2]), .B(n10), .C(r_SM_Main[0]), 
         .D(r_SM_Main[1]), .Z(n13050)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i3_4_lut.init = 16'h0800;
    LUT4 i24_2_lut (.A(r_Bit_Index[0]), .B(r_Bit_Index[1]), .Z(n10)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i24_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_rep_157_3_lut_4_lut (.A(r_SM_Main[2]), .B(r_SM_Main[1]), 
         .C(r_SM_Main[0]), .D(r_SM_Main_2__N_2417[2]), .Z(n13750)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;
    defparam i1_2_lut_rep_157_3_lut_4_lut.init = 16'hfbff;
    LUT4 i2_3_lut (.A(r_Bit_Index[1]), .B(r_Bit_Index[2]), .C(r_Bit_Index[0]), 
         .Z(n8940)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i1_4_lut_adj_32 (.A(r_Clock_Count[9]), .B(r_Clock_Count[14]), .C(r_Clock_Count[7]), 
         .D(r_Clock_Count[15]), .Z(n13171)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(83[17:52])
    defparam i1_4_lut_adj_32.init = 16'hfffe;
    LUT4 i1_2_lut_adj_33 (.A(r_Clock_Count[12]), .B(r_Clock_Count[8]), .Z(n13163)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(83[17:52])
    defparam i1_2_lut_adj_33.init = 16'heeee;
    LUT4 i1_2_lut_adj_34 (.A(r_Clock_Count[13]), .B(r_Clock_Count[10]), 
         .Z(n13161)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(83[17:52])
    defparam i1_2_lut_adj_34.init = 16'heeee;
    LUT4 r_Bit_Index_1__bdd_4_lut_6136 (.A(r_Bit_Index[1]), .B(r_Bit_Index[0]), 
         .C(r_SM_Main[0]), .D(r_Bit_Index[2]), .Z(n13870)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C+!(D)))+!A (C+!(D)))) */ ;
    defparam r_Bit_Index_1__bdd_4_lut_6136.init = 16'h0708;
    FD1P3IX r_Clock_Count_932__i15 (.D(n69[15]), .SP(UartClk_2_enable_56), 
            .CD(n8362), .CK(\UartClk[2] ), .Q(r_Clock_Count[15])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932__i15.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_932__i14 (.D(n69[14]), .SP(UartClk_2_enable_56), 
            .CD(n8362), .CK(\UartClk[2] ), .Q(r_Clock_Count[14])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932__i14.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_932__i13 (.D(n69[13]), .SP(UartClk_2_enable_56), 
            .CD(n8362), .CK(\UartClk[2] ), .Q(r_Clock_Count[13])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932__i13.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_932__i12 (.D(n69[12]), .SP(UartClk_2_enable_56), 
            .CD(n8362), .CK(\UartClk[2] ), .Q(r_Clock_Count[12])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932__i12.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_932__i11 (.D(n69[11]), .SP(UartClk_2_enable_56), 
            .CD(n8362), .CK(\UartClk[2] ), .Q(r_Clock_Count[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932__i11.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_932__i10 (.D(n69[10]), .SP(UartClk_2_enable_56), 
            .CD(n8362), .CK(\UartClk[2] ), .Q(r_Clock_Count[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932__i10.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_932__i9 (.D(n69[9]), .SP(UartClk_2_enable_56), 
            .CD(n8362), .CK(\UartClk[2] ), .Q(r_Clock_Count[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932__i9.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_932__i8 (.D(n69[8]), .SP(UartClk_2_enable_56), 
            .CD(n8362), .CK(\UartClk[2] ), .Q(r_Clock_Count[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932__i8.GSR = "ENABLED";
    PFUMX i6028 (.BLUT(n13780), .ALUT(n13781), .C0(r_SM_Main[0]), .Z(n13782));
    FD1P3IX r_Clock_Count_932__i7 (.D(n69[7]), .SP(UartClk_2_enable_56), 
            .CD(n8362), .CK(\UartClk[2] ), .Q(r_Clock_Count[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932__i7.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_932__i6 (.D(n69[6]), .SP(UartClk_2_enable_56), 
            .CD(n8362), .CK(\UartClk[2] ), .Q(r_Clock_Count[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932__i6.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i0 (.D(r_Rx_Data), .SP(UartClk_2_enable_52), .CK(\UartClk[2] ), 
            .Q(r_Rx_Byte[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=32, LSE_RCOL=2, LSE_LLINE=176, LSE_RLINE=181 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(64[10] 160[8])
    defparam r_Rx_Byte_i0.GSR = "ENABLED";
    PFUMX i5927 (.BLUT(n13544), .ALUT(n13543), .C0(r_SM_Main[1]), .Z(n13545));
    FD1P3IX r_Clock_Count_932__i5 (.D(n69[5]), .SP(UartClk_2_enable_56), 
            .CD(n8362), .CK(\UartClk[2] ), .Q(r_Clock_Count[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932__i5.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_932__i4 (.D(n69[4]), .SP(UartClk_2_enable_56), 
            .CD(n8362), .CK(\UartClk[2] ), .Q(r_Clock_Count[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932__i4.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_932__i3 (.D(n69[3]), .SP(UartClk_2_enable_56), 
            .CD(n8362), .CK(\UartClk[2] ), .Q(r_Clock_Count[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932__i3.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_932__i2 (.D(n69[2]), .SP(UartClk_2_enable_56), 
            .CD(n8362), .CK(\UartClk[2] ), .Q(r_Clock_Count[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/uartrx.v(135[34:54])
    defparam r_Clock_Count_932__i2.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module AMDemodulator
//

module AMDemodulator (CIC1_out_clkSin, \CIC1_outSin[0] , CIC1_outCos, 
            \DataInReg_11__N_1855[0] , GND_net, \CIC1_outSin[1] , \CIC1_outSin[2] , 
            \CIC1_outSin[3] , \CIC1_outSin[4] , \CIC1_outSin[5] , MYLED_c_0, 
            MYLED_c_1, MYLED_c_2, MYLED_c_3, MYLED_c_4, MYLED_c_5, 
            \DataInReg_11__N_1855[1] , \DataInReg_11__N_1855[2] , \DataInReg_11__N_1855[3] , 
            \DataInReg_11__N_1855[4] , \DataInReg_11__N_1855[5] , \DataInReg_11__N_1855[6] , 
            \DataInReg_11__N_1855[7] , \DataInReg_11__N_1855[8] , \DemodOut[9] , 
            VCC_net) /* synthesis syn_module_defined=1 */ ;
    input CIC1_out_clkSin;
    input \CIC1_outSin[0] ;
    input [11:0]CIC1_outCos;
    output \DataInReg_11__N_1855[0] ;
    input GND_net;
    input \CIC1_outSin[1] ;
    input \CIC1_outSin[2] ;
    input \CIC1_outSin[3] ;
    input \CIC1_outSin[4] ;
    input \CIC1_outSin[5] ;
    input MYLED_c_0;
    input MYLED_c_1;
    input MYLED_c_2;
    input MYLED_c_3;
    input MYLED_c_4;
    input MYLED_c_5;
    output \DataInReg_11__N_1855[1] ;
    output \DataInReg_11__N_1855[2] ;
    output \DataInReg_11__N_1855[3] ;
    output \DataInReg_11__N_1855[4] ;
    output \DataInReg_11__N_1855[5] ;
    output \DataInReg_11__N_1855[6] ;
    output \DataInReg_11__N_1855[7] ;
    output \DataInReg_11__N_1855[8] ;
    output \DemodOut[9] ;
    input VCC_net;
    
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(67[6:21])
    wire [11:0]MultDataB;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(29[21:30])
    wire [11:0]MultDataC;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(33[21:30])
    wire [31:0]ISquare;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(24[14:21])
    wire [31:0]ISquare_31__N_1894;
    wire [15:0]d_out_d;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(20[21:28])
    wire [23:0]MultResult1;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(30[22:33])
    wire [23:0]MultResult2;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(35[22:33])
    wire [17:0]d_out_d_11__N_1873;
    
    wire d_out_d_11__N_1872;
    wire [17:0]d_out_d_11__N_1893;
    wire [17:0]d_out_d_11__N_1871;
    
    wire d_out_d_11__N_1870, n12271, n12275, n12274, n209, n12273, 
        n12269;
    wire [17:0]d_out_d_11__N_1891;
    wire [17:0]d_out_d_11__N_2352;
    
    wire n12268, n12267, n12266;
    wire [17:0]d_out_d_11__N_1875;
    
    wire n12265;
    wire [17:0]d_out_d_11__N_1879;
    wire [17:0]d_out_d_11__N_1877;
    
    wire n12264;
    wire [17:0]d_out_d_11__N_1883;
    wire [17:0]d_out_d_11__N_1881;
    
    wire n12263;
    wire [17:0]d_out_d_11__N_1887;
    wire [17:0]d_out_d_11__N_1885;
    
    wire n12262;
    wire [17:0]d_out_d_11__N_1889;
    
    wire n11209, n11208, n11207, n11206, n11205, n11204, n11203, 
        n11202, n11201, n12233, n12232, n12231, n12230, n12229, 
        n12228, n12227, n12226, n12225, d_out_d_11__N_1890, d_out_d_11__N_1888, 
        d_out_d_11__N_1886, d_out_d_11__N_1884, d_out_d_11__N_1882, d_out_d_11__N_1880, 
        d_out_d_11__N_1878, d_out_d_11__N_1876, d_out_d_11__N_1874, n11001, 
        n11000, n10999, n10998, n10997, n10996, n10995, n10994, 
        n10993, n10992, n10991, n10990, n12184;
    wire [17:0]d_out_d_11__N_2334;
    
    wire n12183, n12182, n12181, n12180, n11548, n11547, n11546, 
        n11545, n11544, n11543, n11542, n11536, n11535, n11534, 
        n11533, n11532, n11531, n11525, n11524, n11523, n11522, 
        n11521, n11515, n11514, n11513, n11512, n11511, n11510, 
        n11509, n11508, n11507, n11501, n11500, n11499, n11498, 
        n11497, n11496, n11495, n11494, n11493, n12179, n12178, 
        n12177, n12175, n12174, n12173, n12172, n12171, n12170, 
        n12169, n12168, n12162, n12161, n12160, n12159, n12158, 
        n12157, n12156, n12155, n12154, n12148, n12147, n12146, 
        n12145, n12144, n12143, n12142, n12141, n12140;
    
    FD1S3AX MultDataB_i0 (.D(\CIC1_outSin[0] ), .CK(CIC1_out_clkSin), .Q(MultDataB[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i0.GSR = "ENABLED";
    FD1S3AX MultDataC_i0 (.D(CIC1_outCos[0]), .CK(CIC1_out_clkSin), .Q(MultDataC[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i0.GSR = "ENABLED";
    FD1S3AX ISquare_i1 (.D(ISquare_31__N_1894[0]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i1.GSR = "ENABLED";
    FD1S3AX d_out_i1 (.D(d_out_d[0]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1855[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i1.GSR = "ENABLED";
    LUT4 i4758_2_lut (.A(MultResult1[0]), .B(MultResult2[0]), .Z(ISquare_31__N_1894[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4758_2_lut.init = 16'h6666;
    LUT4 d_out_d_11__I_1_1_lut (.A(d_out_d_11__N_1873[17]), .Z(d_out_d_11__N_1872)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_1_1_lut.init = 16'h5555;
    FD1S3AX d_out_d__0_i1 (.D(d_out_d_11__N_1893[17]), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i1.GSR = "ENABLED";
    LUT4 d_out_d_11__I_0_1_lut (.A(d_out_d_11__N_1871[17]), .Z(d_out_d_11__N_1870)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_0_1_lut.init = 16'h5555;
    LUT4 i4829_2_lut (.A(ISquare[23]), .B(ISquare[22]), .Z(n12271)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i4829_2_lut.init = 16'h9999;
    CCU2D add_3288_8 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n12275), 
          .S0(d_out_d_11__N_1871[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_3288_8.INIT0 = 16'h0fff;
    defparam add_3288_8.INIT1 = 16'h0000;
    defparam add_3288_8.INJECT1_0 = "NO";
    defparam add_3288_8.INJECT1_1 = "NO";
    CCU2D add_3288_6 (.A0(n209), .B0(ISquare[31]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n12274), 
          .COUT(n12275), .S0(d_out_d_11__N_1871[4]), .S1(d_out_d_11__N_1871[5]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_3288_6.INIT0 = 16'h5666;
    defparam add_3288_6.INIT1 = 16'h0fff;
    defparam add_3288_6.INJECT1_0 = "NO";
    defparam add_3288_6.INJECT1_1 = "NO";
    CCU2D add_3288_4 (.A0(n209), .B0(ISquare[31]), .C0(GND_net), .D0(GND_net), 
          .A1(ISquare[31]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n12273), .COUT(n12274), .S0(d_out_d_11__N_1871[2]), .S1(d_out_d_11__N_1871[3]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_3288_4.INIT0 = 16'h5666;
    defparam add_3288_4.INIT1 = 16'h0555;
    defparam add_3288_4.INJECT1_0 = "NO";
    defparam add_3288_4.INJECT1_1 = "NO";
    CCU2D add_3288_2 (.A0(ISquare[23]), .B0(ISquare[22]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n12273), .S1(d_out_d_11__N_1871[1]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_3288_2.INIT0 = 16'h1000;
    defparam add_3288_2.INIT1 = 16'h0fff;
    defparam add_3288_2.INJECT1_0 = "NO";
    defparam add_3288_2.INJECT1_1 = "NO";
    CCU2D add_148_17 (.A0(d_out_d_11__N_1891[14]), .B0(ISquare[31]), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1891[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12269), .S1(d_out_d_11__N_2352[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_148_17.INIT0 = 16'h5666;
    defparam add_148_17.INIT1 = 16'h5aaa;
    defparam add_148_17.INJECT1_0 = "NO";
    defparam add_148_17.INJECT1_1 = "NO";
    CCU2D add_148_15 (.A0(d_out_d_11__N_1891[12]), .B0(ISquare[31]), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1891[13]), .B1(ISquare[31]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12268), .COUT(n12269));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_148_15.INIT0 = 16'h5666;
    defparam add_148_15.INIT1 = 16'h5666;
    defparam add_148_15.INJECT1_0 = "NO";
    defparam add_148_15.INJECT1_1 = "NO";
    CCU2D add_148_13 (.A0(d_out_d_11__N_1891[10]), .B0(d_out_d_11__N_1871[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1891[11]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12267), .COUT(n12268));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_148_13.INIT0 = 16'h5999;
    defparam add_148_13.INIT1 = 16'h5aaa;
    defparam add_148_13.INJECT1_0 = "NO";
    defparam add_148_13.INJECT1_1 = "NO";
    CCU2D add_148_11 (.A0(d_out_d_11__N_1891[8]), .B0(d_out_d_11__N_1875[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1891[9]), .B1(d_out_d_11__N_1873[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12266), .COUT(n12267));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_148_11.INIT0 = 16'h5999;
    defparam add_148_11.INIT1 = 16'h5999;
    defparam add_148_11.INJECT1_0 = "NO";
    defparam add_148_11.INJECT1_1 = "NO";
    CCU2D add_148_9 (.A0(d_out_d_11__N_1891[6]), .B0(d_out_d_11__N_1879[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1891[7]), .B1(d_out_d_11__N_1877[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12265), .COUT(n12266));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_148_9.INIT0 = 16'h5999;
    defparam add_148_9.INIT1 = 16'h5999;
    defparam add_148_9.INJECT1_0 = "NO";
    defparam add_148_9.INJECT1_1 = "NO";
    CCU2D add_148_7 (.A0(d_out_d_11__N_1891[4]), .B0(d_out_d_11__N_1883[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1891[5]), .B1(d_out_d_11__N_1881[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12264), .COUT(n12265));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_148_7.INIT0 = 16'h5999;
    defparam add_148_7.INIT1 = 16'h5999;
    defparam add_148_7.INJECT1_0 = "NO";
    defparam add_148_7.INJECT1_1 = "NO";
    CCU2D add_148_5 (.A0(d_out_d_11__N_1891[2]), .B0(d_out_d_11__N_1887[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1891[3]), .B1(d_out_d_11__N_1885[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12263), .COUT(n12264));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_148_5.INIT0 = 16'h5999;
    defparam add_148_5.INIT1 = 16'h5999;
    defparam add_148_5.INJECT1_0 = "NO";
    defparam add_148_5.INJECT1_1 = "NO";
    CCU2D add_148_3 (.A0(d_out_d_11__N_1891[0]), .B0(d_out_d_11__N_1891[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1891[1]), .B1(d_out_d_11__N_1889[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12262), .COUT(n12263));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_148_3.INIT0 = 16'h5999;
    defparam add_148_3.INIT1 = 16'h5999;
    defparam add_148_3.INJECT1_0 = "NO";
    defparam add_148_3.INJECT1_1 = "NO";
    CCU2D add_148_1 (.A0(ISquare[0]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(ISquare[1]), .B1(d_out_d_11__N_1891[17]), .C1(GND_net), 
          .D1(GND_net), .COUT(n12262));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(58[15:27])
    defparam add_148_1.INIT0 = 16'h5000;
    defparam add_148_1.INIT1 = 16'h5666;
    defparam add_148_1.INJECT1_0 = "NO";
    defparam add_148_1.INJECT1_1 = "NO";
    FD1S3AX MultDataB_i1 (.D(\CIC1_outSin[1] ), .CK(CIC1_out_clkSin), .Q(MultDataB[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i1.GSR = "ENABLED";
    FD1S3AX MultDataB_i2 (.D(\CIC1_outSin[2] ), .CK(CIC1_out_clkSin), .Q(MultDataB[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i2.GSR = "ENABLED";
    FD1S3AX MultDataB_i3 (.D(\CIC1_outSin[3] ), .CK(CIC1_out_clkSin), .Q(MultDataB[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i3.GSR = "ENABLED";
    FD1S3AX MultDataB_i4 (.D(\CIC1_outSin[4] ), .CK(CIC1_out_clkSin), .Q(MultDataB[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i4.GSR = "ENABLED";
    FD1S3AX MultDataB_i5 (.D(\CIC1_outSin[5] ), .CK(CIC1_out_clkSin), .Q(MultDataB[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i5.GSR = "ENABLED";
    FD1S3AX MultDataB_i6 (.D(MYLED_c_0), .CK(CIC1_out_clkSin), .Q(MultDataB[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i6.GSR = "ENABLED";
    FD1S3AX MultDataB_i7 (.D(MYLED_c_1), .CK(CIC1_out_clkSin), .Q(MultDataB[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i7.GSR = "ENABLED";
    FD1S3AX MultDataB_i8 (.D(MYLED_c_2), .CK(CIC1_out_clkSin), .Q(MultDataB[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i8.GSR = "ENABLED";
    FD1S3AX MultDataB_i9 (.D(MYLED_c_3), .CK(CIC1_out_clkSin), .Q(MultDataB[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i9.GSR = "ENABLED";
    FD1S3AX MultDataB_i10 (.D(MYLED_c_4), .CK(CIC1_out_clkSin), .Q(MultDataB[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i10.GSR = "ENABLED";
    FD1S3AX MultDataB_i11 (.D(MYLED_c_5), .CK(CIC1_out_clkSin), .Q(MultDataB[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataB_i11.GSR = "ENABLED";
    FD1S3AX MultDataC_i1 (.D(CIC1_outCos[1]), .CK(CIC1_out_clkSin), .Q(MultDataC[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i1.GSR = "ENABLED";
    FD1S3AX MultDataC_i2 (.D(CIC1_outCos[2]), .CK(CIC1_out_clkSin), .Q(MultDataC[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i2.GSR = "ENABLED";
    FD1S3AX MultDataC_i3 (.D(CIC1_outCos[3]), .CK(CIC1_out_clkSin), .Q(MultDataC[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i3.GSR = "ENABLED";
    FD1S3AX MultDataC_i4 (.D(CIC1_outCos[4]), .CK(CIC1_out_clkSin), .Q(MultDataC[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i4.GSR = "ENABLED";
    FD1S3AX MultDataC_i5 (.D(CIC1_outCos[5]), .CK(CIC1_out_clkSin), .Q(MultDataC[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i5.GSR = "ENABLED";
    FD1S3AX MultDataC_i6 (.D(CIC1_outCos[6]), .CK(CIC1_out_clkSin), .Q(MultDataC[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i6.GSR = "ENABLED";
    FD1S3AX MultDataC_i7 (.D(CIC1_outCos[7]), .CK(CIC1_out_clkSin), .Q(MultDataC[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i7.GSR = "ENABLED";
    FD1S3AX MultDataC_i8 (.D(CIC1_outCos[8]), .CK(CIC1_out_clkSin), .Q(MultDataC[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i8.GSR = "ENABLED";
    FD1S3AX MultDataC_i9 (.D(CIC1_outCos[9]), .CK(CIC1_out_clkSin), .Q(MultDataC[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i9.GSR = "ENABLED";
    FD1S3AX MultDataC_i10 (.D(CIC1_outCos[10]), .CK(CIC1_out_clkSin), .Q(MultDataC[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i10.GSR = "ENABLED";
    FD1S3AX MultDataC_i11 (.D(CIC1_outCos[11]), .CK(CIC1_out_clkSin), .Q(MultDataC[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam MultDataC_i11.GSR = "ENABLED";
    FD1S3AX ISquare_i2 (.D(ISquare_31__N_1894[1]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i2.GSR = "ENABLED";
    FD1S3AX ISquare_i3 (.D(ISquare_31__N_1894[2]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i3.GSR = "ENABLED";
    FD1S3AX ISquare_i4 (.D(ISquare_31__N_1894[3]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i4.GSR = "ENABLED";
    FD1S3AX ISquare_i5 (.D(ISquare_31__N_1894[4]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i5.GSR = "ENABLED";
    FD1S3AX ISquare_i6 (.D(ISquare_31__N_1894[5]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i6.GSR = "ENABLED";
    FD1S3AX ISquare_i7 (.D(ISquare_31__N_1894[6]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i7.GSR = "ENABLED";
    FD1S3AX ISquare_i8 (.D(ISquare_31__N_1894[7]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i8.GSR = "ENABLED";
    FD1S3AX ISquare_i9 (.D(ISquare_31__N_1894[8]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i9.GSR = "ENABLED";
    FD1S3AX ISquare_i10 (.D(ISquare_31__N_1894[9]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i10.GSR = "ENABLED";
    FD1S3AX ISquare_i11 (.D(ISquare_31__N_1894[10]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i11.GSR = "ENABLED";
    FD1S3AX ISquare_i12 (.D(ISquare_31__N_1894[11]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i12.GSR = "ENABLED";
    FD1S3AX ISquare_i13 (.D(ISquare_31__N_1894[12]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i13.GSR = "ENABLED";
    FD1S3AX ISquare_i14 (.D(ISquare_31__N_1894[13]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i14.GSR = "ENABLED";
    FD1S3AX ISquare_i15 (.D(ISquare_31__N_1894[14]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i15.GSR = "ENABLED";
    FD1S3AX ISquare_i16 (.D(ISquare_31__N_1894[15]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i16.GSR = "ENABLED";
    FD1S3AX ISquare_i17 (.D(ISquare_31__N_1894[16]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i17.GSR = "ENABLED";
    FD1S3AX ISquare_i18 (.D(ISquare_31__N_1894[17]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i18.GSR = "ENABLED";
    FD1S3AX ISquare_i19 (.D(ISquare_31__N_1894[18]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i19.GSR = "ENABLED";
    FD1S3AX ISquare_i20 (.D(ISquare_31__N_1894[19]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i20.GSR = "ENABLED";
    FD1S3AX ISquare_i21 (.D(ISquare_31__N_1894[20]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i21.GSR = "ENABLED";
    FD1S3AX ISquare_i22 (.D(ISquare_31__N_1894[21]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i22.GSR = "ENABLED";
    FD1S3AX ISquare_i23 (.D(ISquare_31__N_1894[22]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i23.GSR = "ENABLED";
    FD1S3AX ISquare_i24 (.D(ISquare_31__N_1894[23]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i24.GSR = "ENABLED";
    FD1S3AX ISquare_i25 (.D(ISquare_31__N_1894[24]), .CK(CIC1_out_clkSin), 
            .Q(ISquare[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam ISquare_i25.GSR = "ENABLED";
    FD1S3AX d_out_i2 (.D(d_out_d[1]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1855[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i2.GSR = "ENABLED";
    FD1S3AX d_out_i3 (.D(d_out_d[2]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1855[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i3.GSR = "ENABLED";
    FD1S3AX d_out_i4 (.D(d_out_d[3]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1855[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i4.GSR = "ENABLED";
    FD1S3AX d_out_i5 (.D(d_out_d[4]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1855[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i5.GSR = "ENABLED";
    FD1S3AX d_out_i6 (.D(d_out_d[5]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1855[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i6.GSR = "ENABLED";
    FD1S3AX d_out_i7 (.D(d_out_d[6]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1855[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i7.GSR = "ENABLED";
    FD1S3AX d_out_i8 (.D(d_out_d[7]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1855[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i8.GSR = "ENABLED";
    FD1S3AX d_out_i9 (.D(d_out_d[8]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1855[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i9.GSR = "ENABLED";
    FD1S3AX d_out_i10 (.D(d_out_d[9]), .CK(CIC1_out_clkSin), .Q(\DemodOut[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=10, LSE_LLINE=168, LSE_RLINE=173 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_i10.GSR = "ENABLED";
    CCU2D add_437_19 (.A0(d_out_d_11__N_1887[14]), .B0(d_out_d_11__N_1887[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1887[15]), .B1(d_out_d_11__N_1887[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11209), .S0(d_out_d_11__N_1889[15]), 
          .S1(d_out_d_11__N_1889[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_437_19.INIT0 = 16'h5999;
    defparam add_437_19.INIT1 = 16'h5999;
    defparam add_437_19.INJECT1_0 = "NO";
    defparam add_437_19.INJECT1_1 = "NO";
    CCU2D add_437_17 (.A0(ISquare[31]), .B0(d_out_d_11__N_1887[17]), .C0(d_out_d_11__N_1887[12]), 
          .D0(GND_net), .A1(d_out_d_11__N_1887[13]), .B1(d_out_d_11__N_1887[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11208), .COUT(n11209), .S0(d_out_d_11__N_1889[13]), 
          .S1(d_out_d_11__N_1889[14]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_437_17.INIT0 = 16'h6969;
    defparam add_437_17.INIT1 = 16'h5999;
    defparam add_437_17.INJECT1_0 = "NO";
    defparam add_437_17.INJECT1_1 = "NO";
    CCU2D add_437_15 (.A0(ISquare[31]), .B0(d_out_d_11__N_1887[17]), .C0(d_out_d_11__N_1887[10]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1887[17]), 
          .C1(d_out_d_11__N_1887[11]), .D1(GND_net), .CIN(n11207), .COUT(n11208), 
          .S0(d_out_d_11__N_1889[11]), .S1(d_out_d_11__N_1889[12]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_437_15.INIT0 = 16'h6969;
    defparam add_437_15.INIT1 = 16'h6969;
    defparam add_437_15.INJECT1_0 = "NO";
    defparam add_437_15.INJECT1_1 = "NO";
    CCU2D add_437_13 (.A0(d_out_d_11__N_1871[17]), .B0(d_out_d_11__N_1887[17]), 
          .C0(d_out_d_11__N_1887[8]), .D0(GND_net), .A1(d_out_d_11__N_1887[9]), 
          .B1(d_out_d_11__N_1887[17]), .C1(GND_net), .D1(GND_net), .CIN(n11206), 
          .COUT(n11207), .S0(d_out_d_11__N_1889[9]), .S1(d_out_d_11__N_1889[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_437_13.INIT0 = 16'h9696;
    defparam add_437_13.INIT1 = 16'h5999;
    defparam add_437_13.INJECT1_0 = "NO";
    defparam add_437_13.INJECT1_1 = "NO";
    CCU2D add_437_11 (.A0(d_out_d_11__N_1875[17]), .B0(d_out_d_11__N_1887[17]), 
          .C0(d_out_d_11__N_1887[6]), .D0(GND_net), .A1(d_out_d_11__N_1873[17]), 
          .B1(d_out_d_11__N_1887[17]), .C1(d_out_d_11__N_1887[7]), .D1(GND_net), 
          .CIN(n11205), .COUT(n11206), .S0(d_out_d_11__N_1889[7]), .S1(d_out_d_11__N_1889[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_437_11.INIT0 = 16'h9696;
    defparam add_437_11.INIT1 = 16'h9696;
    defparam add_437_11.INJECT1_0 = "NO";
    defparam add_437_11.INJECT1_1 = "NO";
    CCU2D add_437_9 (.A0(d_out_d_11__N_1879[17]), .B0(d_out_d_11__N_1887[17]), 
          .C0(d_out_d_11__N_1887[4]), .D0(GND_net), .A1(d_out_d_11__N_1877[17]), 
          .B1(d_out_d_11__N_1887[17]), .C1(d_out_d_11__N_1887[5]), .D1(GND_net), 
          .CIN(n11204), .COUT(n11205), .S0(d_out_d_11__N_1889[5]), .S1(d_out_d_11__N_1889[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_437_9.INIT0 = 16'h9696;
    defparam add_437_9.INIT1 = 16'h9696;
    defparam add_437_9.INJECT1_0 = "NO";
    defparam add_437_9.INJECT1_1 = "NO";
    CCU2D add_437_7 (.A0(d_out_d_11__N_1883[17]), .B0(d_out_d_11__N_1887[17]), 
          .C0(d_out_d_11__N_1887[2]), .D0(GND_net), .A1(d_out_d_11__N_1881[17]), 
          .B1(d_out_d_11__N_1887[17]), .C1(d_out_d_11__N_1887[3]), .D1(GND_net), 
          .CIN(n11203), .COUT(n11204), .S0(d_out_d_11__N_1889[3]), .S1(d_out_d_11__N_1889[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_437_7.INIT0 = 16'h9696;
    defparam add_437_7.INIT1 = 16'h9696;
    defparam add_437_7.INJECT1_0 = "NO";
    defparam add_437_7.INJECT1_1 = "NO";
    CCU2D add_437_5 (.A0(d_out_d_11__N_1887[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1885[17]), .B1(d_out_d_11__N_1887[17]), 
          .C1(d_out_d_11__N_1887[1]), .D1(GND_net), .CIN(n11202), .COUT(n11203), 
          .S0(d_out_d_11__N_1889[1]), .S1(d_out_d_11__N_1889[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_437_5.INIT0 = 16'h5aaa;
    defparam add_437_5.INIT1 = 16'h9696;
    defparam add_437_5.INJECT1_0 = "NO";
    defparam add_437_5.INJECT1_1 = "NO";
    CCU2D add_437_3 (.A0(ISquare[4]), .B0(d_out_d_11__N_1887[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11201), .COUT(n11202), .S1(d_out_d_11__N_1889[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_437_3.INIT0 = 16'h5666;
    defparam add_437_3.INIT1 = 16'h5555;
    defparam add_437_3.INJECT1_0 = "NO";
    defparam add_437_3.INJECT1_1 = "NO";
    CCU2D add_437_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1887[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n11201));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_437_1.INIT0 = 16'hF000;
    defparam add_437_1.INIT1 = 16'h0aaa;
    defparam add_437_1.INJECT1_0 = "NO";
    defparam add_437_1.INJECT1_1 = "NO";
    CCU2D add_457_19 (.A0(d_out_d_11__N_1885[14]), .B0(d_out_d_11__N_1885[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1885[15]), .B1(d_out_d_11__N_1885[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12233), .S0(d_out_d_11__N_1887[15]), 
          .S1(d_out_d_11__N_1887[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_457_19.INIT0 = 16'h5999;
    defparam add_457_19.INIT1 = 16'h5999;
    defparam add_457_19.INJECT1_0 = "NO";
    defparam add_457_19.INJECT1_1 = "NO";
    CCU2D add_457_17 (.A0(d_out_d_11__N_1885[12]), .B0(d_out_d_11__N_1885[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1885[13]), .B1(d_out_d_11__N_1885[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12232), .COUT(n12233), .S0(d_out_d_11__N_1887[13]), 
          .S1(d_out_d_11__N_1887[14]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_457_17.INIT0 = 16'h5999;
    defparam add_457_17.INIT1 = 16'h5999;
    defparam add_457_17.INJECT1_0 = "NO";
    defparam add_457_17.INJECT1_1 = "NO";
    CCU2D add_457_15 (.A0(ISquare[31]), .B0(d_out_d_11__N_1885[17]), .C0(d_out_d_11__N_1885[10]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1885[17]), 
          .C1(d_out_d_11__N_1885[11]), .D1(GND_net), .CIN(n12231), .COUT(n12232), 
          .S0(d_out_d_11__N_1887[11]), .S1(d_out_d_11__N_1887[12]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_457_15.INIT0 = 16'h6969;
    defparam add_457_15.INIT1 = 16'h6969;
    defparam add_457_15.INJECT1_0 = "NO";
    defparam add_457_15.INJECT1_1 = "NO";
    CCU2D add_457_13 (.A0(d_out_d_11__N_1885[8]), .B0(d_out_d_11__N_1885[17]), 
          .C0(GND_net), .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1885[17]), 
          .C1(d_out_d_11__N_1885[9]), .D1(GND_net), .CIN(n12230), .COUT(n12231), 
          .S0(d_out_d_11__N_1887[9]), .S1(d_out_d_11__N_1887[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_457_13.INIT0 = 16'h5999;
    defparam add_457_13.INIT1 = 16'h6969;
    defparam add_457_13.INJECT1_0 = "NO";
    defparam add_457_13.INJECT1_1 = "NO";
    CCU2D add_457_11 (.A0(d_out_d_11__N_1873[17]), .B0(d_out_d_11__N_1885[17]), 
          .C0(d_out_d_11__N_1885[6]), .D0(GND_net), .A1(d_out_d_11__N_1871[17]), 
          .B1(d_out_d_11__N_1885[17]), .C1(d_out_d_11__N_1885[7]), .D1(GND_net), 
          .CIN(n12229), .COUT(n12230), .S0(d_out_d_11__N_1887[7]), .S1(d_out_d_11__N_1887[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_457_11.INIT0 = 16'h9696;
    defparam add_457_11.INIT1 = 16'h9696;
    defparam add_457_11.INJECT1_0 = "NO";
    defparam add_457_11.INJECT1_1 = "NO";
    CCU2D add_457_9 (.A0(d_out_d_11__N_1877[17]), .B0(d_out_d_11__N_1885[17]), 
          .C0(d_out_d_11__N_1885[4]), .D0(GND_net), .A1(d_out_d_11__N_1875[17]), 
          .B1(d_out_d_11__N_1885[17]), .C1(d_out_d_11__N_1885[5]), .D1(GND_net), 
          .CIN(n12228), .COUT(n12229), .S0(d_out_d_11__N_1887[5]), .S1(d_out_d_11__N_1887[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_457_9.INIT0 = 16'h9696;
    defparam add_457_9.INIT1 = 16'h9696;
    defparam add_457_9.INJECT1_0 = "NO";
    defparam add_457_9.INJECT1_1 = "NO";
    CCU2D add_457_7 (.A0(d_out_d_11__N_1881[17]), .B0(d_out_d_11__N_1885[17]), 
          .C0(d_out_d_11__N_1885[2]), .D0(GND_net), .A1(d_out_d_11__N_1879[17]), 
          .B1(d_out_d_11__N_1885[17]), .C1(d_out_d_11__N_1885[3]), .D1(GND_net), 
          .CIN(n12227), .COUT(n12228), .S0(d_out_d_11__N_1887[3]), .S1(d_out_d_11__N_1887[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_457_7.INIT0 = 16'h9696;
    defparam add_457_7.INIT1 = 16'h9696;
    defparam add_457_7.INJECT1_0 = "NO";
    defparam add_457_7.INJECT1_1 = "NO";
    CCU2D add_457_5 (.A0(d_out_d_11__N_1885[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1883[17]), .B1(d_out_d_11__N_1885[17]), 
          .C1(d_out_d_11__N_1885[1]), .D1(GND_net), .CIN(n12226), .COUT(n12227), 
          .S0(d_out_d_11__N_1887[1]), .S1(d_out_d_11__N_1887[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_457_5.INIT0 = 16'h5aaa;
    defparam add_457_5.INIT1 = 16'h9696;
    defparam add_457_5.INJECT1_0 = "NO";
    defparam add_457_5.INJECT1_1 = "NO";
    CCU2D add_457_3 (.A0(ISquare[6]), .B0(d_out_d_11__N_1885[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12225), .COUT(n12226), .S1(d_out_d_11__N_1887[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_457_3.INIT0 = 16'h5666;
    defparam add_457_3.INIT1 = 16'h5555;
    defparam add_457_3.INJECT1_0 = "NO";
    defparam add_457_3.INJECT1_1 = "NO";
    CCU2D add_457_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1885[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n12225));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_457_1.INIT0 = 16'hF000;
    defparam add_457_1.INIT1 = 16'h0aaa;
    defparam add_457_1.INJECT1_0 = "NO";
    defparam add_457_1.INJECT1_1 = "NO";
    LUT4 d_out_d_11__I_10_1_lut (.A(d_out_d_11__N_1891[17]), .Z(d_out_d_11__N_1890)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_10_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_9_1_lut (.A(d_out_d_11__N_1889[17]), .Z(d_out_d_11__N_1888)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_9_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_8_1_lut (.A(d_out_d_11__N_1887[17]), .Z(d_out_d_11__N_1886)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_8_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_7_1_lut (.A(d_out_d_11__N_1885[17]), .Z(d_out_d_11__N_1884)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_7_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_6_1_lut (.A(d_out_d_11__N_1883[17]), .Z(d_out_d_11__N_1882)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_6_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_5_1_lut (.A(d_out_d_11__N_1881[17]), .Z(d_out_d_11__N_1880)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_5_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_4_1_lut (.A(d_out_d_11__N_1879[17]), .Z(d_out_d_11__N_1878)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_4_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_3_1_lut (.A(d_out_d_11__N_1877[17]), .Z(d_out_d_11__N_1876)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_3_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_2_1_lut (.A(d_out_d_11__N_1875[17]), .Z(d_out_d_11__N_1874)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(61[22:28])
    defparam d_out_d_11__I_2_1_lut.init = 16'h5555;
    FD1S3AX d_out_d__0_i2 (.D(d_out_d_11__N_1890), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[1]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i2.GSR = "ENABLED";
    CCU2D MultResult1_23__I_0_26 (.A0(MultResult1[23]), .B0(MultResult2[23]), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11001), .S0(ISquare_31__N_1894[24]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_26.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_26.INIT1 = 16'h0000;
    defparam MultResult1_23__I_0_26.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_26.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_24 (.A0(MultResult1[22]), .B0(MultResult2[22]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[23]), .B1(MultResult2[23]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11000), .COUT(n11001), .S0(ISquare_31__N_1894[22]), 
          .S1(ISquare_31__N_1894[23]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_24.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_24.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_24.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_24.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_22 (.A0(MultResult1[20]), .B0(MultResult2[20]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[21]), .B1(MultResult2[21]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10999), .COUT(n11000), .S0(ISquare_31__N_1894[20]), 
          .S1(ISquare_31__N_1894[21]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_22.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_22.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_22.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_22.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_20 (.A0(MultResult1[18]), .B0(MultResult2[18]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[19]), .B1(MultResult2[19]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10998), .COUT(n10999), .S0(ISquare_31__N_1894[18]), 
          .S1(ISquare_31__N_1894[19]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_20.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_20.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_20.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_20.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_18 (.A0(MultResult1[16]), .B0(MultResult2[16]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[17]), .B1(MultResult2[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10997), .COUT(n10998), .S0(ISquare_31__N_1894[16]), 
          .S1(ISquare_31__N_1894[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_18.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_18.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_18.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_18.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_16 (.A0(MultResult1[14]), .B0(MultResult2[14]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[15]), .B1(MultResult2[15]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10996), .COUT(n10997), .S0(ISquare_31__N_1894[14]), 
          .S1(ISquare_31__N_1894[15]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_16.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_16.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_16.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_16.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_14 (.A0(MultResult1[12]), .B0(MultResult2[12]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[13]), .B1(MultResult2[13]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10995), .COUT(n10996), .S0(ISquare_31__N_1894[12]), 
          .S1(ISquare_31__N_1894[13]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_14.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_14.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_14.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_14.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_12 (.A0(MultResult1[10]), .B0(MultResult2[10]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[11]), .B1(MultResult2[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10994), .COUT(n10995), .S0(ISquare_31__N_1894[10]), 
          .S1(ISquare_31__N_1894[11]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_12.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_12.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_12.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_12.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_10 (.A0(MultResult1[8]), .B0(MultResult2[8]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[9]), .B1(MultResult2[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10993), .COUT(n10994), .S0(ISquare_31__N_1894[8]), 
          .S1(ISquare_31__N_1894[9]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_10.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_10.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_10.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_10.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_8 (.A0(MultResult1[6]), .B0(MultResult2[6]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[7]), .B1(MultResult2[7]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10992), .COUT(n10993), .S0(ISquare_31__N_1894[6]), 
          .S1(ISquare_31__N_1894[7]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_8.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_8.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_8.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_8.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_6 (.A0(MultResult1[4]), .B0(MultResult2[4]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[5]), .B1(MultResult2[5]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10991), .COUT(n10992), .S0(ISquare_31__N_1894[4]), 
          .S1(ISquare_31__N_1894[5]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_6.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_6.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_6.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_6.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_4 (.A0(MultResult1[2]), .B0(MultResult2[2]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[3]), .B1(MultResult2[3]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10990), .COUT(n10991), .S0(ISquare_31__N_1894[2]), 
          .S1(ISquare_31__N_1894[3]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_4.INIT0 = 16'h5666;
    defparam MultResult1_23__I_0_4.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_4.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_4.INJECT1_1 = "NO";
    CCU2D MultResult1_23__I_0_2 (.A0(MultResult1[0]), .B0(MultResult2[0]), 
          .C0(GND_net), .D0(GND_net), .A1(MultResult1[1]), .B1(MultResult2[1]), 
          .C1(GND_net), .D1(GND_net), .COUT(n10990), .S1(ISquare_31__N_1894[1]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(92[16:41])
    defparam MultResult1_23__I_0_2.INIT0 = 16'h7000;
    defparam MultResult1_23__I_0_2.INIT1 = 16'h5666;
    defparam MultResult1_23__I_0_2.INJECT1_0 = "NO";
    defparam MultResult1_23__I_0_2.INJECT1_1 = "NO";
    FD1S3AX d_out_d__0_i3 (.D(d_out_d_11__N_1888), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i3.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i4 (.D(d_out_d_11__N_1886), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[3]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i4.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i5 (.D(d_out_d_11__N_1884), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i5.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i6 (.D(d_out_d_11__N_1882), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[5]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i6.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i7 (.D(d_out_d_11__N_1880), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i7.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i8 (.D(d_out_d_11__N_1878), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[7]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i8.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i9 (.D(d_out_d_11__N_1876), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i9.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i10 (.D(d_out_d_11__N_1874), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[9]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(86[9] 95[6])
    defparam d_out_d__0_i10.GSR = "ENABLED";
    CCU2D sub_78_add_2_18 (.A0(d_out_d_11__N_1891[14]), .B0(ISquare[31]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1891[15]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12184), .S1(d_out_d_11__N_2334[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_18.INIT0 = 16'h5999;
    defparam sub_78_add_2_18.INIT1 = 16'h5555;
    defparam sub_78_add_2_18.INJECT1_0 = "NO";
    defparam sub_78_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_16 (.A0(d_out_d_11__N_1891[12]), .B0(ISquare[31]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1891[13]), .B1(ISquare[31]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12183), .COUT(n12184));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_16.INIT0 = 16'h5999;
    defparam sub_78_add_2_16.INIT1 = 16'h5999;
    defparam sub_78_add_2_16.INJECT1_0 = "NO";
    defparam sub_78_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_14 (.A0(d_out_d_11__N_1891[10]), .B0(d_out_d_11__N_1871[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1891[11]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n12182), .COUT(n12183));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_14.INIT0 = 16'h5666;
    defparam sub_78_add_2_14.INIT1 = 16'h5555;
    defparam sub_78_add_2_14.INJECT1_0 = "NO";
    defparam sub_78_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_12 (.A0(d_out_d_11__N_1891[8]), .B0(d_out_d_11__N_1875[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1891[9]), .B1(d_out_d_11__N_1873[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12181), .COUT(n12182));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_12.INIT0 = 16'h5666;
    defparam sub_78_add_2_12.INIT1 = 16'h5666;
    defparam sub_78_add_2_12.INJECT1_0 = "NO";
    defparam sub_78_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_10 (.A0(d_out_d_11__N_1891[6]), .B0(d_out_d_11__N_1879[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1891[7]), .B1(d_out_d_11__N_1877[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12180), .COUT(n12181));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_10.INIT0 = 16'h5666;
    defparam sub_78_add_2_10.INIT1 = 16'h5666;
    defparam sub_78_add_2_10.INJECT1_0 = "NO";
    defparam sub_78_add_2_10.INJECT1_1 = "NO";
    CCU2D add_577_15 (.A0(d_out_d_11__N_1875[17]), .B0(d_out_d_11__N_1874), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1875[17]), .B1(d_out_d_11__N_1874), 
          .C1(GND_net), .D1(GND_net), .CIN(n11548), .S0(d_out_d_11__N_1877[11]), 
          .S1(d_out_d_11__N_1877[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_577_15.INIT0 = 16'h5666;
    defparam add_577_15.INIT1 = 16'h5666;
    defparam add_577_15.INJECT1_0 = "NO";
    defparam add_577_15.INJECT1_1 = "NO";
    CCU2D add_577_13 (.A0(d_out_d_11__N_1875[8]), .B0(d_out_d_11__N_1875[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1875[9]), .B1(d_out_d_11__N_1875[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11547), .COUT(n11548), .S0(d_out_d_11__N_1877[9]), 
          .S1(d_out_d_11__N_1877[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_577_13.INIT0 = 16'h5999;
    defparam add_577_13.INIT1 = 16'h5999;
    defparam add_577_13.INJECT1_0 = "NO";
    defparam add_577_13.INJECT1_1 = "NO";
    CCU2D add_577_11 (.A0(ISquare[31]), .B0(d_out_d_11__N_1875[17]), .C0(d_out_d_11__N_1875[6]), 
          .D0(GND_net), .A1(d_out_d_11__N_1875[7]), .B1(d_out_d_11__N_1875[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11546), .COUT(n11547), .S0(d_out_d_11__N_1877[7]), 
          .S1(d_out_d_11__N_1877[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_577_11.INIT0 = 16'h6969;
    defparam add_577_11.INIT1 = 16'h5999;
    defparam add_577_11.INJECT1_0 = "NO";
    defparam add_577_11.INJECT1_1 = "NO";
    CCU2D add_577_9 (.A0(ISquare[31]), .B0(d_out_d_11__N_1875[17]), .C0(d_out_d_11__N_1875[4]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1875[17]), 
          .C1(d_out_d_11__N_1875[5]), .D1(GND_net), .CIN(n11545), .COUT(n11546), 
          .S0(d_out_d_11__N_1877[5]), .S1(d_out_d_11__N_1877[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_577_9.INIT0 = 16'h6969;
    defparam add_577_9.INIT1 = 16'h6969;
    defparam add_577_9.INJECT1_0 = "NO";
    defparam add_577_9.INJECT1_1 = "NO";
    CCU2D add_577_7 (.A0(d_out_d_11__N_1871[17]), .B0(d_out_d_11__N_1875[17]), 
          .C0(d_out_d_11__N_1875[2]), .D0(GND_net), .A1(d_out_d_11__N_1875[3]), 
          .B1(d_out_d_11__N_1875[17]), .C1(GND_net), .D1(GND_net), .CIN(n11544), 
          .COUT(n11545), .S0(d_out_d_11__N_1877[3]), .S1(d_out_d_11__N_1877[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_577_7.INIT0 = 16'h9696;
    defparam add_577_7.INIT1 = 16'h5999;
    defparam add_577_7.INJECT1_0 = "NO";
    defparam add_577_7.INJECT1_1 = "NO";
    CCU2D add_577_5 (.A0(d_out_d_11__N_1875[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1873[17]), .B1(d_out_d_11__N_1875[17]), 
          .C1(d_out_d_11__N_1875[1]), .D1(GND_net), .CIN(n11543), .COUT(n11544), 
          .S0(d_out_d_11__N_1877[1]), .S1(d_out_d_11__N_1877[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_577_5.INIT0 = 16'h5aaa;
    defparam add_577_5.INIT1 = 16'h9696;
    defparam add_577_5.INJECT1_0 = "NO";
    defparam add_577_5.INJECT1_1 = "NO";
    CCU2D add_577_3 (.A0(ISquare[16]), .B0(d_out_d_11__N_1875[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11542), .COUT(n11543), .S1(d_out_d_11__N_1877[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_577_3.INIT0 = 16'h5666;
    defparam add_577_3.INIT1 = 16'h5555;
    defparam add_577_3.INJECT1_0 = "NO";
    defparam add_577_3.INJECT1_1 = "NO";
    CCU2D add_577_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1875[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n11542));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_577_1.INIT0 = 16'hF000;
    defparam add_577_1.INIT1 = 16'h0aaa;
    defparam add_577_1.INJECT1_0 = "NO";
    defparam add_577_1.INJECT1_1 = "NO";
    CCU2D add_597_13 (.A0(d_out_d_11__N_1873[17]), .B0(d_out_d_11__N_1872), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1873[17]), .B1(d_out_d_11__N_1872), 
          .C1(GND_net), .D1(GND_net), .CIN(n11536), .S0(d_out_d_11__N_1875[9]), 
          .S1(d_out_d_11__N_1875[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_597_13.INIT0 = 16'h5666;
    defparam add_597_13.INIT1 = 16'h5666;
    defparam add_597_13.INJECT1_0 = "NO";
    defparam add_597_13.INJECT1_1 = "NO";
    CCU2D add_597_11 (.A0(d_out_d_11__N_1873[6]), .B0(d_out_d_11__N_1873[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1873[7]), .B1(d_out_d_11__N_1873[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11535), .COUT(n11536), .S0(d_out_d_11__N_1875[7]), 
          .S1(d_out_d_11__N_1875[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_597_11.INIT0 = 16'h5999;
    defparam add_597_11.INIT1 = 16'h5999;
    defparam add_597_11.INJECT1_0 = "NO";
    defparam add_597_11.INJECT1_1 = "NO";
    CCU2D add_597_9 (.A0(ISquare[31]), .B0(d_out_d_11__N_1873[17]), .C0(d_out_d_11__N_1873[4]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1873[17]), 
          .C1(d_out_d_11__N_1873[5]), .D1(GND_net), .CIN(n11534), .COUT(n11535), 
          .S0(d_out_d_11__N_1875[5]), .S1(d_out_d_11__N_1875[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_597_9.INIT0 = 16'h6969;
    defparam add_597_9.INIT1 = 16'h6969;
    defparam add_597_9.INJECT1_0 = "NO";
    defparam add_597_9.INJECT1_1 = "NO";
    CCU2D add_597_7 (.A0(d_out_d_11__N_1873[2]), .B0(d_out_d_11__N_1873[17]), 
          .C0(GND_net), .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1873[17]), 
          .C1(d_out_d_11__N_1873[3]), .D1(GND_net), .CIN(n11533), .COUT(n11534), 
          .S0(d_out_d_11__N_1875[3]), .S1(d_out_d_11__N_1875[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_597_7.INIT0 = 16'h5999;
    defparam add_597_7.INIT1 = 16'h6969;
    defparam add_597_7.INJECT1_0 = "NO";
    defparam add_597_7.INJECT1_1 = "NO";
    CCU2D add_597_5 (.A0(d_out_d_11__N_1873[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1871[17]), .B1(d_out_d_11__N_1873[17]), 
          .C1(d_out_d_11__N_1873[1]), .D1(GND_net), .CIN(n11532), .COUT(n11533), 
          .S0(d_out_d_11__N_1875[1]), .S1(d_out_d_11__N_1875[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_597_5.INIT0 = 16'h5aaa;
    defparam add_597_5.INIT1 = 16'h9696;
    defparam add_597_5.INJECT1_0 = "NO";
    defparam add_597_5.INJECT1_1 = "NO";
    CCU2D add_597_3 (.A0(ISquare[18]), .B0(d_out_d_11__N_1873[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11531), .COUT(n11532), .S1(d_out_d_11__N_1875[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_597_3.INIT0 = 16'h5666;
    defparam add_597_3.INIT1 = 16'h5555;
    defparam add_597_3.INJECT1_0 = "NO";
    defparam add_597_3.INJECT1_1 = "NO";
    CCU2D add_597_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1873[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n11531));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_597_1.INIT0 = 16'hF000;
    defparam add_597_1.INIT1 = 16'h0aaa;
    defparam add_597_1.INJECT1_0 = "NO";
    defparam add_597_1.INJECT1_1 = "NO";
    CCU2D add_617_11 (.A0(d_out_d_11__N_1871[17]), .B0(d_out_d_11__N_1870), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1871[17]), .B1(d_out_d_11__N_1870), 
          .C1(GND_net), .D1(GND_net), .CIN(n11525), .S0(d_out_d_11__N_1873[7]), 
          .S1(d_out_d_11__N_1873[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_617_11.INIT0 = 16'h5666;
    defparam add_617_11.INIT1 = 16'h5666;
    defparam add_617_11.INJECT1_0 = "NO";
    defparam add_617_11.INJECT1_1 = "NO";
    CCU2D add_617_9 (.A0(ISquare[31]), .B0(d_out_d_11__N_1871[17]), .C0(d_out_d_11__N_1871[4]), 
          .D0(GND_net), .A1(d_out_d_11__N_1871[5]), .B1(d_out_d_11__N_1871[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11524), .COUT(n11525), .S0(d_out_d_11__N_1873[5]), 
          .S1(d_out_d_11__N_1873[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_617_9.INIT0 = 16'h6969;
    defparam add_617_9.INIT1 = 16'h5999;
    defparam add_617_9.INJECT1_0 = "NO";
    defparam add_617_9.INJECT1_1 = "NO";
    CCU2D add_617_7 (.A0(ISquare[31]), .B0(d_out_d_11__N_1871[17]), .C0(d_out_d_11__N_1871[2]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1871[17]), 
          .C1(d_out_d_11__N_1871[3]), .D1(GND_net), .CIN(n11523), .COUT(n11524), 
          .S0(d_out_d_11__N_1873[3]), .S1(d_out_d_11__N_1873[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_617_7.INIT0 = 16'h6969;
    defparam add_617_7.INIT1 = 16'h6969;
    defparam add_617_7.INJECT1_0 = "NO";
    defparam add_617_7.INJECT1_1 = "NO";
    CCU2D add_617_5 (.A0(n12271), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1871[1]), .B1(d_out_d_11__N_1871[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n11522), .COUT(n11523), .S0(d_out_d_11__N_1873[1]), 
          .S1(d_out_d_11__N_1873[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_617_5.INIT0 = 16'h5aaa;
    defparam add_617_5.INIT1 = 16'h5999;
    defparam add_617_5.INJECT1_0 = "NO";
    defparam add_617_5.INJECT1_1 = "NO";
    CCU2D add_617_3 (.A0(ISquare[20]), .B0(d_out_d_11__N_1871[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11521), .COUT(n11522), .S1(d_out_d_11__N_1873[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_617_3.INIT0 = 16'h5666;
    defparam add_617_3.INIT1 = 16'h5555;
    defparam add_617_3.INJECT1_0 = "NO";
    defparam add_617_3.INJECT1_1 = "NO";
    CCU2D add_617_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1871[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n11521));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_617_1.INIT0 = 16'hF000;
    defparam add_617_1.INIT1 = 16'h0aaa;
    defparam add_617_1.INJECT1_0 = "NO";
    defparam add_617_1.INJECT1_1 = "NO";
    CCU2D add_537_19 (.A0(d_out_d_11__N_1879[17]), .B0(d_out_d_11__N_1878), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1879[17]), .B1(d_out_d_11__N_1878), 
          .C1(GND_net), .D1(GND_net), .CIN(n11515), .S0(d_out_d_11__N_1881[15]), 
          .S1(d_out_d_11__N_1881[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_537_19.INIT0 = 16'h5666;
    defparam add_537_19.INIT1 = 16'h5666;
    defparam add_537_19.INJECT1_0 = "NO";
    defparam add_537_19.INJECT1_1 = "NO";
    CCU2D add_537_17 (.A0(d_out_d_11__N_1879[12]), .B0(d_out_d_11__N_1879[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1879[13]), .B1(d_out_d_11__N_1879[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11514), .COUT(n11515), .S0(d_out_d_11__N_1881[13]), 
          .S1(d_out_d_11__N_1881[14]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_537_17.INIT0 = 16'h5999;
    defparam add_537_17.INIT1 = 16'h5999;
    defparam add_537_17.INJECT1_0 = "NO";
    defparam add_537_17.INJECT1_1 = "NO";
    CCU2D add_537_15 (.A0(d_out_d_11__N_1879[10]), .B0(d_out_d_11__N_1879[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1879[11]), .B1(d_out_d_11__N_1879[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11513), .COUT(n11514), .S0(d_out_d_11__N_1881[11]), 
          .S1(d_out_d_11__N_1881[12]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_537_15.INIT0 = 16'h5999;
    defparam add_537_15.INIT1 = 16'h5999;
    defparam add_537_15.INJECT1_0 = "NO";
    defparam add_537_15.INJECT1_1 = "NO";
    CCU2D add_537_13 (.A0(ISquare[31]), .B0(d_out_d_11__N_1879[17]), .C0(d_out_d_11__N_1879[8]), 
          .D0(GND_net), .A1(d_out_d_11__N_1879[9]), .B1(d_out_d_11__N_1879[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11512), .COUT(n11513), .S0(d_out_d_11__N_1881[9]), 
          .S1(d_out_d_11__N_1881[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_537_13.INIT0 = 16'h6969;
    defparam add_537_13.INIT1 = 16'h5999;
    defparam add_537_13.INJECT1_0 = "NO";
    defparam add_537_13.INJECT1_1 = "NO";
    CCU2D add_537_11 (.A0(ISquare[31]), .B0(d_out_d_11__N_1879[17]), .C0(d_out_d_11__N_1879[6]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1879[17]), 
          .C1(d_out_d_11__N_1879[7]), .D1(GND_net), .CIN(n11511), .COUT(n11512), 
          .S0(d_out_d_11__N_1881[7]), .S1(d_out_d_11__N_1881[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_537_11.INIT0 = 16'h6969;
    defparam add_537_11.INIT1 = 16'h6969;
    defparam add_537_11.INJECT1_0 = "NO";
    defparam add_537_11.INJECT1_1 = "NO";
    CCU2D add_537_9 (.A0(d_out_d_11__N_1871[17]), .B0(d_out_d_11__N_1879[17]), 
          .C0(d_out_d_11__N_1879[4]), .D0(GND_net), .A1(d_out_d_11__N_1879[5]), 
          .B1(d_out_d_11__N_1879[17]), .C1(GND_net), .D1(GND_net), .CIN(n11510), 
          .COUT(n11511), .S0(d_out_d_11__N_1881[5]), .S1(d_out_d_11__N_1881[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_537_9.INIT0 = 16'h9696;
    defparam add_537_9.INIT1 = 16'h5999;
    defparam add_537_9.INJECT1_0 = "NO";
    defparam add_537_9.INJECT1_1 = "NO";
    CCU2D add_537_7 (.A0(d_out_d_11__N_1875[17]), .B0(d_out_d_11__N_1879[17]), 
          .C0(d_out_d_11__N_1879[2]), .D0(GND_net), .A1(d_out_d_11__N_1873[17]), 
          .B1(d_out_d_11__N_1879[17]), .C1(d_out_d_11__N_1879[3]), .D1(GND_net), 
          .CIN(n11509), .COUT(n11510), .S0(d_out_d_11__N_1881[3]), .S1(d_out_d_11__N_1881[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_537_7.INIT0 = 16'h9696;
    defparam add_537_7.INIT1 = 16'h9696;
    defparam add_537_7.INJECT1_0 = "NO";
    defparam add_537_7.INJECT1_1 = "NO";
    CCU2D add_537_5 (.A0(d_out_d_11__N_1879[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1877[17]), .B1(d_out_d_11__N_1879[17]), 
          .C1(d_out_d_11__N_1879[1]), .D1(GND_net), .CIN(n11508), .COUT(n11509), 
          .S0(d_out_d_11__N_1881[1]), .S1(d_out_d_11__N_1881[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_537_5.INIT0 = 16'h5aaa;
    defparam add_537_5.INIT1 = 16'h9696;
    defparam add_537_5.INJECT1_0 = "NO";
    defparam add_537_5.INJECT1_1 = "NO";
    CCU2D add_537_3 (.A0(ISquare[12]), .B0(d_out_d_11__N_1879[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11507), .COUT(n11508), .S1(d_out_d_11__N_1881[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_537_3.INIT0 = 16'h5666;
    defparam add_537_3.INIT1 = 16'h5555;
    defparam add_537_3.INJECT1_0 = "NO";
    defparam add_537_3.INJECT1_1 = "NO";
    CCU2D add_537_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1879[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n11507));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_537_1.INIT0 = 16'hF000;
    defparam add_537_1.INIT1 = 16'h0aaa;
    defparam add_537_1.INJECT1_0 = "NO";
    defparam add_537_1.INJECT1_1 = "NO";
    CCU2D add_477_19 (.A0(d_out_d_11__N_1883[14]), .B0(d_out_d_11__N_1883[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1883[15]), .B1(d_out_d_11__N_1883[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11501), .S0(d_out_d_11__N_1885[15]), 
          .S1(d_out_d_11__N_1885[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_477_19.INIT0 = 16'h5999;
    defparam add_477_19.INIT1 = 16'h5999;
    defparam add_477_19.INJECT1_0 = "NO";
    defparam add_477_19.INJECT1_1 = "NO";
    CCU2D add_477_17 (.A0(d_out_d_11__N_1883[12]), .B0(d_out_d_11__N_1883[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1883[13]), .B1(d_out_d_11__N_1883[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11500), .COUT(n11501), .S0(d_out_d_11__N_1885[13]), 
          .S1(d_out_d_11__N_1885[14]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_477_17.INIT0 = 16'h5999;
    defparam add_477_17.INIT1 = 16'h5999;
    defparam add_477_17.INJECT1_0 = "NO";
    defparam add_477_17.INJECT1_1 = "NO";
    CCU2D add_477_15 (.A0(ISquare[31]), .B0(d_out_d_11__N_1883[17]), .C0(d_out_d_11__N_1883[10]), 
          .D0(GND_net), .A1(d_out_d_11__N_1883[11]), .B1(d_out_d_11__N_1883[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n11499), .COUT(n11500), .S0(d_out_d_11__N_1885[11]), 
          .S1(d_out_d_11__N_1885[12]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_477_15.INIT0 = 16'h6969;
    defparam add_477_15.INIT1 = 16'h5999;
    defparam add_477_15.INJECT1_0 = "NO";
    defparam add_477_15.INJECT1_1 = "NO";
    CCU2D add_477_13 (.A0(ISquare[31]), .B0(d_out_d_11__N_1883[17]), .C0(d_out_d_11__N_1883[8]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1883[17]), 
          .C1(d_out_d_11__N_1883[9]), .D1(GND_net), .CIN(n11498), .COUT(n11499), 
          .S0(d_out_d_11__N_1885[9]), .S1(d_out_d_11__N_1885[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_477_13.INIT0 = 16'h6969;
    defparam add_477_13.INIT1 = 16'h6969;
    defparam add_477_13.INJECT1_0 = "NO";
    defparam add_477_13.INJECT1_1 = "NO";
    CCU2D add_477_11 (.A0(d_out_d_11__N_1871[17]), .B0(d_out_d_11__N_1883[17]), 
          .C0(d_out_d_11__N_1883[6]), .D0(GND_net), .A1(d_out_d_11__N_1883[7]), 
          .B1(d_out_d_11__N_1883[17]), .C1(GND_net), .D1(GND_net), .CIN(n11497), 
          .COUT(n11498), .S0(d_out_d_11__N_1885[7]), .S1(d_out_d_11__N_1885[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_477_11.INIT0 = 16'h9696;
    defparam add_477_11.INIT1 = 16'h5999;
    defparam add_477_11.INJECT1_0 = "NO";
    defparam add_477_11.INJECT1_1 = "NO";
    CCU2D add_477_9 (.A0(d_out_d_11__N_1875[17]), .B0(d_out_d_11__N_1883[17]), 
          .C0(d_out_d_11__N_1883[4]), .D0(GND_net), .A1(d_out_d_11__N_1873[17]), 
          .B1(d_out_d_11__N_1883[17]), .C1(d_out_d_11__N_1883[5]), .D1(GND_net), 
          .CIN(n11496), .COUT(n11497), .S0(d_out_d_11__N_1885[5]), .S1(d_out_d_11__N_1885[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_477_9.INIT0 = 16'h9696;
    defparam add_477_9.INIT1 = 16'h9696;
    defparam add_477_9.INJECT1_0 = "NO";
    defparam add_477_9.INJECT1_1 = "NO";
    CCU2D add_477_7 (.A0(d_out_d_11__N_1879[17]), .B0(d_out_d_11__N_1883[17]), 
          .C0(d_out_d_11__N_1883[2]), .D0(GND_net), .A1(d_out_d_11__N_1877[17]), 
          .B1(d_out_d_11__N_1883[17]), .C1(d_out_d_11__N_1883[3]), .D1(GND_net), 
          .CIN(n11495), .COUT(n11496), .S0(d_out_d_11__N_1885[3]), .S1(d_out_d_11__N_1885[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_477_7.INIT0 = 16'h9696;
    defparam add_477_7.INIT1 = 16'h9696;
    defparam add_477_7.INJECT1_0 = "NO";
    defparam add_477_7.INJECT1_1 = "NO";
    CCU2D add_477_5 (.A0(d_out_d_11__N_1883[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1881[17]), .B1(d_out_d_11__N_1883[17]), 
          .C1(d_out_d_11__N_1883[1]), .D1(GND_net), .CIN(n11494), .COUT(n11495), 
          .S0(d_out_d_11__N_1885[1]), .S1(d_out_d_11__N_1885[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_477_5.INIT0 = 16'h5aaa;
    defparam add_477_5.INIT1 = 16'h9696;
    defparam add_477_5.INJECT1_0 = "NO";
    defparam add_477_5.INJECT1_1 = "NO";
    CCU2D add_477_3 (.A0(ISquare[8]), .B0(d_out_d_11__N_1883[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n11493), .COUT(n11494), .S1(d_out_d_11__N_1885[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_477_3.INIT0 = 16'h5666;
    defparam add_477_3.INIT1 = 16'h5555;
    defparam add_477_3.INJECT1_0 = "NO";
    defparam add_477_3.INJECT1_1 = "NO";
    CCU2D add_477_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1883[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n11493));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_477_1.INIT0 = 16'hF000;
    defparam add_477_1.INIT1 = 16'h0aaa;
    defparam add_477_1.INJECT1_0 = "NO";
    defparam add_477_1.INJECT1_1 = "NO";
    LUT4 mux_74_i1_3_lut (.A(d_out_d_11__N_2334[17]), .B(d_out_d_11__N_2352[17]), 
         .C(d_out_d_11__N_1891[17]), .Z(d_out_d_11__N_1893[17])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam mux_74_i1_3_lut.init = 16'h3535;
    LUT4 i1326_1_lut (.A(ISquare[31]), .Z(n209)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1326_1_lut.init = 16'h5555;
    CCU2D sub_78_add_2_8 (.A0(d_out_d_11__N_1891[4]), .B0(d_out_d_11__N_1883[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1891[5]), .B1(d_out_d_11__N_1881[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12179), .COUT(n12180));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_8.INIT0 = 16'h5666;
    defparam sub_78_add_2_8.INIT1 = 16'h5666;
    defparam sub_78_add_2_8.INJECT1_0 = "NO";
    defparam sub_78_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_6 (.A0(d_out_d_11__N_1891[2]), .B0(d_out_d_11__N_1887[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1891[3]), .B1(d_out_d_11__N_1885[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12178), .COUT(n12179));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_6.INIT0 = 16'h5666;
    defparam sub_78_add_2_6.INIT1 = 16'h5666;
    defparam sub_78_add_2_6.INJECT1_0 = "NO";
    defparam sub_78_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_4 (.A0(d_out_d_11__N_1891[0]), .B0(d_out_d_11__N_1891[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1891[1]), .B1(d_out_d_11__N_1889[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12177), .COUT(n12178));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_4.INIT0 = 16'h5666;
    defparam sub_78_add_2_4.INIT1 = 16'h5666;
    defparam sub_78_add_2_4.INJECT1_0 = "NO";
    defparam sub_78_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_2 (.A0(ISquare[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[1]), .B1(d_out_d_11__N_1891[17]), 
          .C1(GND_net), .D1(GND_net), .COUT(n12177));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[15:27])
    defparam sub_78_add_2_2.INIT0 = 16'h5000;
    defparam sub_78_add_2_2.INIT1 = 16'h5999;
    defparam sub_78_add_2_2.INJECT1_0 = "NO";
    defparam sub_78_add_2_2.INJECT1_1 = "NO";
    CCU2D add_557_17 (.A0(d_out_d_11__N_1877[17]), .B0(d_out_d_11__N_1876), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1877[17]), .B1(d_out_d_11__N_1876), 
          .C1(GND_net), .D1(GND_net), .CIN(n12175), .S0(d_out_d_11__N_1879[13]), 
          .S1(d_out_d_11__N_1879[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_557_17.INIT0 = 16'h5666;
    defparam add_557_17.INIT1 = 16'h5666;
    defparam add_557_17.INJECT1_0 = "NO";
    defparam add_557_17.INJECT1_1 = "NO";
    CCU2D add_557_15 (.A0(d_out_d_11__N_1877[10]), .B0(d_out_d_11__N_1877[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1877[11]), .B1(d_out_d_11__N_1877[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12174), .COUT(n12175), .S0(d_out_d_11__N_1879[11]), 
          .S1(d_out_d_11__N_1879[12]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_557_15.INIT0 = 16'h5999;
    defparam add_557_15.INIT1 = 16'h5999;
    defparam add_557_15.INJECT1_0 = "NO";
    defparam add_557_15.INJECT1_1 = "NO";
    CCU2D add_557_13 (.A0(d_out_d_11__N_1877[8]), .B0(d_out_d_11__N_1877[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1877[9]), .B1(d_out_d_11__N_1877[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12173), .COUT(n12174), .S0(d_out_d_11__N_1879[9]), 
          .S1(d_out_d_11__N_1879[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_557_13.INIT0 = 16'h5999;
    defparam add_557_13.INIT1 = 16'h5999;
    defparam add_557_13.INJECT1_0 = "NO";
    defparam add_557_13.INJECT1_1 = "NO";
    CCU2D add_557_11 (.A0(ISquare[31]), .B0(d_out_d_11__N_1877[17]), .C0(d_out_d_11__N_1877[6]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1877[17]), 
          .C1(d_out_d_11__N_1877[7]), .D1(GND_net), .CIN(n12172), .COUT(n12173), 
          .S0(d_out_d_11__N_1879[7]), .S1(d_out_d_11__N_1879[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_557_11.INIT0 = 16'h6969;
    defparam add_557_11.INIT1 = 16'h6969;
    defparam add_557_11.INJECT1_0 = "NO";
    defparam add_557_11.INJECT1_1 = "NO";
    CCU2D add_557_9 (.A0(d_out_d_11__N_1877[4]), .B0(d_out_d_11__N_1877[17]), 
          .C0(GND_net), .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1877[17]), 
          .C1(d_out_d_11__N_1877[5]), .D1(GND_net), .CIN(n12171), .COUT(n12172), 
          .S0(d_out_d_11__N_1879[5]), .S1(d_out_d_11__N_1879[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_557_9.INIT0 = 16'h5999;
    defparam add_557_9.INIT1 = 16'h6969;
    defparam add_557_9.INJECT1_0 = "NO";
    defparam add_557_9.INJECT1_1 = "NO";
    CCU2D add_557_7 (.A0(d_out_d_11__N_1873[17]), .B0(d_out_d_11__N_1877[17]), 
          .C0(d_out_d_11__N_1877[2]), .D0(GND_net), .A1(d_out_d_11__N_1871[17]), 
          .B1(d_out_d_11__N_1877[17]), .C1(d_out_d_11__N_1877[3]), .D1(GND_net), 
          .CIN(n12170), .COUT(n12171), .S0(d_out_d_11__N_1879[3]), .S1(d_out_d_11__N_1879[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_557_7.INIT0 = 16'h9696;
    defparam add_557_7.INIT1 = 16'h9696;
    defparam add_557_7.INJECT1_0 = "NO";
    defparam add_557_7.INJECT1_1 = "NO";
    CCU2D add_557_5 (.A0(d_out_d_11__N_1877[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1875[17]), .B1(d_out_d_11__N_1877[17]), 
          .C1(d_out_d_11__N_1877[1]), .D1(GND_net), .CIN(n12169), .COUT(n12170), 
          .S0(d_out_d_11__N_1879[1]), .S1(d_out_d_11__N_1879[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_557_5.INIT0 = 16'h5aaa;
    defparam add_557_5.INIT1 = 16'h9696;
    defparam add_557_5.INJECT1_0 = "NO";
    defparam add_557_5.INJECT1_1 = "NO";
    CCU2D add_557_3 (.A0(ISquare[14]), .B0(d_out_d_11__N_1877[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12168), .COUT(n12169), .S1(d_out_d_11__N_1879[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_557_3.INIT0 = 16'h5666;
    defparam add_557_3.INIT1 = 16'h5555;
    defparam add_557_3.INJECT1_0 = "NO";
    defparam add_557_3.INJECT1_1 = "NO";
    CCU2D add_557_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1877[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n12168));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_557_1.INIT0 = 16'hF000;
    defparam add_557_1.INIT1 = 16'h0aaa;
    defparam add_557_1.INJECT1_0 = "NO";
    defparam add_557_1.INJECT1_1 = "NO";
    CCU2D add_497_19 (.A0(d_out_d_11__N_1889[14]), .B0(d_out_d_11__N_1889[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1889[15]), .B1(d_out_d_11__N_1889[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12162), .S0(d_out_d_11__N_1891[15]), 
          .S1(d_out_d_11__N_1891[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_497_19.INIT0 = 16'h5999;
    defparam add_497_19.INIT1 = 16'h5999;
    defparam add_497_19.INJECT1_0 = "NO";
    defparam add_497_19.INJECT1_1 = "NO";
    CCU2D add_497_17 (.A0(ISquare[31]), .B0(d_out_d_11__N_1889[17]), .C0(d_out_d_11__N_1889[12]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1889[17]), 
          .C1(d_out_d_11__N_1889[13]), .D1(GND_net), .CIN(n12161), .COUT(n12162), 
          .S0(d_out_d_11__N_1891[13]), .S1(d_out_d_11__N_1891[14]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_497_17.INIT0 = 16'h6969;
    defparam add_497_17.INIT1 = 16'h6969;
    defparam add_497_17.INJECT1_0 = "NO";
    defparam add_497_17.INJECT1_1 = "NO";
    CCU2D add_497_15 (.A0(d_out_d_11__N_1889[10]), .B0(d_out_d_11__N_1889[17]), 
          .C0(GND_net), .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1889[17]), 
          .C1(d_out_d_11__N_1889[11]), .D1(GND_net), .CIN(n12160), .COUT(n12161), 
          .S0(d_out_d_11__N_1891[11]), .S1(d_out_d_11__N_1891[12]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_497_15.INIT0 = 16'h5999;
    defparam add_497_15.INIT1 = 16'h6969;
    defparam add_497_15.INJECT1_0 = "NO";
    defparam add_497_15.INJECT1_1 = "NO";
    CCU2D add_497_13 (.A0(d_out_d_11__N_1873[17]), .B0(d_out_d_11__N_1889[17]), 
          .C0(d_out_d_11__N_1889[8]), .D0(GND_net), .A1(d_out_d_11__N_1871[17]), 
          .B1(d_out_d_11__N_1889[17]), .C1(d_out_d_11__N_1889[9]), .D1(GND_net), 
          .CIN(n12159), .COUT(n12160), .S0(d_out_d_11__N_1891[9]), .S1(d_out_d_11__N_1891[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_497_13.INIT0 = 16'h9696;
    defparam add_497_13.INIT1 = 16'h9696;
    defparam add_497_13.INJECT1_0 = "NO";
    defparam add_497_13.INJECT1_1 = "NO";
    CCU2D add_497_11 (.A0(d_out_d_11__N_1877[17]), .B0(d_out_d_11__N_1889[17]), 
          .C0(d_out_d_11__N_1889[6]), .D0(GND_net), .A1(d_out_d_11__N_1875[17]), 
          .B1(d_out_d_11__N_1889[17]), .C1(d_out_d_11__N_1889[7]), .D1(GND_net), 
          .CIN(n12158), .COUT(n12159), .S0(d_out_d_11__N_1891[7]), .S1(d_out_d_11__N_1891[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_497_11.INIT0 = 16'h9696;
    defparam add_497_11.INIT1 = 16'h9696;
    defparam add_497_11.INJECT1_0 = "NO";
    defparam add_497_11.INJECT1_1 = "NO";
    CCU2D add_497_9 (.A0(d_out_d_11__N_1881[17]), .B0(d_out_d_11__N_1889[17]), 
          .C0(d_out_d_11__N_1889[4]), .D0(GND_net), .A1(d_out_d_11__N_1879[17]), 
          .B1(d_out_d_11__N_1889[17]), .C1(d_out_d_11__N_1889[5]), .D1(GND_net), 
          .CIN(n12157), .COUT(n12158), .S0(d_out_d_11__N_1891[5]), .S1(d_out_d_11__N_1891[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_497_9.INIT0 = 16'h9696;
    defparam add_497_9.INIT1 = 16'h9696;
    defparam add_497_9.INJECT1_0 = "NO";
    defparam add_497_9.INJECT1_1 = "NO";
    CCU2D add_497_7 (.A0(d_out_d_11__N_1885[17]), .B0(d_out_d_11__N_1889[17]), 
          .C0(d_out_d_11__N_1889[2]), .D0(GND_net), .A1(d_out_d_11__N_1883[17]), 
          .B1(d_out_d_11__N_1889[17]), .C1(d_out_d_11__N_1889[3]), .D1(GND_net), 
          .CIN(n12156), .COUT(n12157), .S0(d_out_d_11__N_1891[3]), .S1(d_out_d_11__N_1891[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_497_7.INIT0 = 16'h9696;
    defparam add_497_7.INIT1 = 16'h9696;
    defparam add_497_7.INJECT1_0 = "NO";
    defparam add_497_7.INJECT1_1 = "NO";
    CCU2D add_497_5 (.A0(d_out_d_11__N_1889[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1887[17]), .B1(d_out_d_11__N_1889[17]), 
          .C1(d_out_d_11__N_1889[1]), .D1(GND_net), .CIN(n12155), .COUT(n12156), 
          .S0(d_out_d_11__N_1891[1]), .S1(d_out_d_11__N_1891[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_497_5.INIT0 = 16'h5aaa;
    defparam add_497_5.INIT1 = 16'h9696;
    defparam add_497_5.INJECT1_0 = "NO";
    defparam add_497_5.INJECT1_1 = "NO";
    CCU2D add_497_3 (.A0(ISquare[2]), .B0(d_out_d_11__N_1889[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12154), .COUT(n12155), .S1(d_out_d_11__N_1891[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_497_3.INIT0 = 16'h5666;
    defparam add_497_3.INIT1 = 16'h5555;
    defparam add_497_3.INJECT1_0 = "NO";
    defparam add_497_3.INJECT1_1 = "NO";
    CCU2D add_497_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1889[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n12154));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_497_1.INIT0 = 16'hF000;
    defparam add_497_1.INIT1 = 16'h0aaa;
    defparam add_497_1.INJECT1_0 = "NO";
    defparam add_497_1.INJECT1_1 = "NO";
    CCU2D add_517_19 (.A0(d_out_d_11__N_1881[14]), .B0(d_out_d_11__N_1881[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1881[15]), .B1(d_out_d_11__N_1881[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12148), .S0(d_out_d_11__N_1883[15]), 
          .S1(d_out_d_11__N_1883[17]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_517_19.INIT0 = 16'h5999;
    defparam add_517_19.INIT1 = 16'h5999;
    defparam add_517_19.INJECT1_0 = "NO";
    defparam add_517_19.INJECT1_1 = "NO";
    CCU2D add_517_17 (.A0(d_out_d_11__N_1881[12]), .B0(d_out_d_11__N_1881[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1881[13]), .B1(d_out_d_11__N_1881[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12147), .COUT(n12148), .S0(d_out_d_11__N_1883[13]), 
          .S1(d_out_d_11__N_1883[14]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_517_17.INIT0 = 16'h5999;
    defparam add_517_17.INIT1 = 16'h5999;
    defparam add_517_17.INJECT1_0 = "NO";
    defparam add_517_17.INJECT1_1 = "NO";
    CCU2D add_517_15 (.A0(d_out_d_11__N_1881[10]), .B0(d_out_d_11__N_1881[17]), 
          .C0(GND_net), .D0(GND_net), .A1(d_out_d_11__N_1881[11]), .B1(d_out_d_11__N_1881[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n12146), .COUT(n12147), .S0(d_out_d_11__N_1883[11]), 
          .S1(d_out_d_11__N_1883[12]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_517_15.INIT0 = 16'h5999;
    defparam add_517_15.INIT1 = 16'h5999;
    defparam add_517_15.INJECT1_0 = "NO";
    defparam add_517_15.INJECT1_1 = "NO";
    CCU2D add_517_13 (.A0(ISquare[31]), .B0(d_out_d_11__N_1881[17]), .C0(d_out_d_11__N_1881[8]), 
          .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1881[17]), 
          .C1(d_out_d_11__N_1881[9]), .D1(GND_net), .CIN(n12145), .COUT(n12146), 
          .S0(d_out_d_11__N_1883[9]), .S1(d_out_d_11__N_1883[10]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_517_13.INIT0 = 16'h6969;
    defparam add_517_13.INIT1 = 16'h6969;
    defparam add_517_13.INJECT1_0 = "NO";
    defparam add_517_13.INJECT1_1 = "NO";
    CCU2D add_517_11 (.A0(d_out_d_11__N_1881[6]), .B0(d_out_d_11__N_1881[17]), 
          .C0(GND_net), .D0(GND_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1881[17]), 
          .C1(d_out_d_11__N_1881[7]), .D1(GND_net), .CIN(n12144), .COUT(n12145), 
          .S0(d_out_d_11__N_1883[7]), .S1(d_out_d_11__N_1883[8]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_517_11.INIT0 = 16'h5999;
    defparam add_517_11.INIT1 = 16'h6969;
    defparam add_517_11.INJECT1_0 = "NO";
    defparam add_517_11.INJECT1_1 = "NO";
    CCU2D add_517_9 (.A0(d_out_d_11__N_1873[17]), .B0(d_out_d_11__N_1881[17]), 
          .C0(d_out_d_11__N_1881[4]), .D0(GND_net), .A1(d_out_d_11__N_1871[17]), 
          .B1(d_out_d_11__N_1881[17]), .C1(d_out_d_11__N_1881[5]), .D1(GND_net), 
          .CIN(n12143), .COUT(n12144), .S0(d_out_d_11__N_1883[5]), .S1(d_out_d_11__N_1883[6]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_517_9.INIT0 = 16'h9696;
    defparam add_517_9.INIT1 = 16'h9696;
    defparam add_517_9.INJECT1_0 = "NO";
    defparam add_517_9.INJECT1_1 = "NO";
    CCU2D add_517_7 (.A0(d_out_d_11__N_1877[17]), .B0(d_out_d_11__N_1881[17]), 
          .C0(d_out_d_11__N_1881[2]), .D0(GND_net), .A1(d_out_d_11__N_1875[17]), 
          .B1(d_out_d_11__N_1881[17]), .C1(d_out_d_11__N_1881[3]), .D1(GND_net), 
          .CIN(n12142), .COUT(n12143), .S0(d_out_d_11__N_1883[3]), .S1(d_out_d_11__N_1883[4]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_517_7.INIT0 = 16'h9696;
    defparam add_517_7.INIT1 = 16'h9696;
    defparam add_517_7.INJECT1_0 = "NO";
    defparam add_517_7.INJECT1_1 = "NO";
    CCU2D add_517_5 (.A0(d_out_d_11__N_1881[0]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(d_out_d_11__N_1879[17]), .B1(d_out_d_11__N_1881[17]), 
          .C1(d_out_d_11__N_1881[1]), .D1(GND_net), .CIN(n12141), .COUT(n12142), 
          .S0(d_out_d_11__N_1883[1]), .S1(d_out_d_11__N_1883[2]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_517_5.INIT0 = 16'h5aaa;
    defparam add_517_5.INIT1 = 16'h9696;
    defparam add_517_5.INJECT1_0 = "NO";
    defparam add_517_5.INJECT1_1 = "NO";
    CCU2D add_517_3 (.A0(ISquare[10]), .B0(d_out_d_11__N_1881[17]), .C0(GND_net), 
          .D0(GND_net), .A1(ISquare[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n12140), .COUT(n12141), .S1(d_out_d_11__N_1883[0]));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_517_3.INIT0 = 16'h5666;
    defparam add_517_3.INIT1 = 16'h5555;
    defparam add_517_3.INJECT1_0 = "NO";
    defparam add_517_3.INJECT1_1 = "NO";
    CCU2D add_517_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(d_out_d_11__N_1881[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n12140));   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(60[11:28])
    defparam add_517_1.INIT0 = 16'hF000;
    defparam add_517_1.INIT1 = 16'h0aaa;
    defparam add_517_1.INJECT1_0 = "NO";
    defparam add_517_1.INJECT1_1 = "NO";
    Multiplier Multiplier2 (.CIC1_out_clkSin(CIC1_out_clkSin), .VCC_net(VCC_net), 
            .GND_net(GND_net), .MultDataC({MultDataC}), .MultResult2({MultResult2})) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    Multiplier_U0 Multiplier1 (.CIC1_out_clkSin(CIC1_out_clkSin), .VCC_net(VCC_net), 
            .GND_net(GND_net), .MultDataB({MultDataB}), .MultResult1({MultResult1})) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    
endmodule
//
// Verilog Description of module Multiplier
//

module Multiplier (CIC1_out_clkSin, VCC_net, GND_net, MultDataC, MultResult2) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input CIC1_out_clkSin;
    input VCC_net;
    input GND_net;
    input [11:0]MultDataC;
    output [23:0]MultResult2;
    
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(67[6:21])
    
    wire Multiplier_0_mult_0_5_n1, regb_b_1, rega_a_11, Multiplier_0_pp_1_2, 
        regb_b_2, regb_b_0, Multiplier_0_mult_2_5_n1, regb_b_3, Multiplier_0_pp_2_4, 
        regb_b_4, Multiplier_0_mult_4_5_n1, regb_b_5, Multiplier_0_pp_3_6, 
        regb_b_6, Multiplier_0_mult_6_5_n1, regb_b_7, Multiplier_0_pp_4_8, 
        regb_b_8, Multiplier_0_mult_8_5_n1, regb_b_9, Multiplier_0_pp_5_10, 
        regb_b_10, Multiplier_0_mult_10_0_n0, regb_b_11, Multiplier_0_mult_10_1_n1, 
        rega_a_3, rega_a_2, Multiplier_0_mult_10_1_n0, Multiplier_0_mult_10_2_n1, 
        rega_a_5, rega_a_4, Multiplier_0_mult_10_2_n0, Multiplier_0_mult_10_3_n1, 
        rega_a_7, rega_a_6, Multiplier_0_mult_10_3_n0, Multiplier_0_mult_10_4_n1, 
        rega_a_9, rega_a_8, Multiplier_0_mult_10_4_n0, Multiplier_0_mult_10_5_n2, 
        rega_a_10, Multiplier_0_mult_10_5_n0, rega_a_1, rego_o_0, rego_o_1, 
        rego_o_2, rego_o_3, rego_o_4, rego_o_5, rego_o_6, rego_o_7, 
        rego_o_8, rego_o_9, rego_o_10, rego_o_11, rego_o_12, rego_o_13, 
        rego_o_14, rego_o_15, rego_o_16, rego_o_17, rego_o_18, rego_o_19, 
        rego_o_20, rego_o_21, rego_o_22, rego_o_23, Multiplier_0_pp_0_0, 
        Multiplier_0_pp_0_1, s_Multiplier_0_0_2, s_Multiplier_0_0_3, s_Multiplier_0_0_4, 
        f_s_Multiplier_0_0_4, s_Multiplier_0_0_5, f_s_Multiplier_0_0_5, 
        s_Multiplier_0_0_6, f_s_Multiplier_0_0_6, s_Multiplier_0_0_7, 
        f_s_Multiplier_0_0_7, s_Multiplier_0_0_8, f_s_Multiplier_0_0_8, 
        s_Multiplier_0_0_9, f_s_Multiplier_0_0_9, s_Multiplier_0_0_10, 
        f_s_Multiplier_0_0_10, s_Multiplier_0_0_11, f_s_Multiplier_0_0_11, 
        s_Multiplier_0_0_12, f_s_Multiplier_0_0_12, s_Multiplier_0_0_13, 
        f_s_Multiplier_0_0_13, s_Multiplier_0_0_14, f_s_Multiplier_0_0_14, 
        s_Multiplier_0_0_15, f_s_Multiplier_0_0_15, s_Multiplier_0_0_16, 
        f_s_Multiplier_0_0_16, s_Multiplier_0_0_17, f_s_Multiplier_0_0_17, 
        f_Multiplier_0_pp_2_4, f_Multiplier_0_pp_2_5, Multiplier_0_pp_2_5, 
        s_Multiplier_0_1_6, f_s_Multiplier_0_1_6, s_Multiplier_0_1_7, 
        f_s_Multiplier_0_1_7, s_Multiplier_0_1_8, f_s_Multiplier_0_1_8, 
        s_Multiplier_0_1_9, f_s_Multiplier_0_1_9, s_Multiplier_0_1_10, 
        f_s_Multiplier_0_1_10, s_Multiplier_0_1_11, f_s_Multiplier_0_1_11, 
        s_Multiplier_0_1_12, f_s_Multiplier_0_1_12, s_Multiplier_0_1_13, 
        f_s_Multiplier_0_1_13, s_Multiplier_0_1_14, f_s_Multiplier_0_1_14, 
        s_Multiplier_0_1_15, f_s_Multiplier_0_1_15, s_Multiplier_0_1_16, 
        f_s_Multiplier_0_1_16, s_Multiplier_0_1_17, f_s_Multiplier_0_1_17, 
        s_Multiplier_0_1_18, f_s_Multiplier_0_1_18, s_Multiplier_0_1_19, 
        f_s_Multiplier_0_1_19, s_Multiplier_0_1_20, f_s_Multiplier_0_1_20, 
        s_Multiplier_0_1_21, f_s_Multiplier_0_1_21, f_Multiplier_0_pp_4_8, 
        f_Multiplier_0_pp_4_9, Multiplier_0_pp_4_9, s_Multiplier_0_2_10, 
        f_s_Multiplier_0_2_10, s_Multiplier_0_2_11, f_s_Multiplier_0_2_11, 
        s_Multiplier_0_2_12, f_s_Multiplier_0_2_12, s_Multiplier_0_2_13, 
        f_s_Multiplier_0_2_13, s_Multiplier_0_2_14, f_s_Multiplier_0_2_14, 
        s_Multiplier_0_2_15, f_s_Multiplier_0_2_15, s_Multiplier_0_2_16, 
        f_s_Multiplier_0_2_16, s_Multiplier_0_2_17, f_s_Multiplier_0_2_17, 
        s_Multiplier_0_2_18, f_s_Multiplier_0_2_18, s_Multiplier_0_2_19, 
        f_s_Multiplier_0_2_19, s_Multiplier_0_2_20, f_s_Multiplier_0_2_20, 
        s_Multiplier_0_2_21, f_s_Multiplier_0_2_21, s_Multiplier_0_2_22, 
        f_s_Multiplier_0_2_22, s_Multiplier_0_2_23, f_s_Multiplier_0_2_23, 
        Multiplier_0_cin_lr_0, Multiplier_0_pp_0_13, mfco, Multiplier_0_cin_lr_2, 
        Multiplier_0_pp_1_15, mfco_1, Multiplier_0_cin_lr_4, Multiplier_0_pp_2_17, 
        mfco_2, Multiplier_0_cin_lr_6, Multiplier_0_pp_3_19, mfco_3, 
        Multiplier_0_cin_lr_8, Multiplier_0_pp_4_21, mfco_4, Multiplier_0_cin_lr_10, 
        Multiplier_0_pp_5_23, mfco_5, co_Multiplier_0_0_1, Multiplier_0_pp_0_2, 
        co_Multiplier_0_0_2, Multiplier_0_pp_0_4, Multiplier_0_pp_0_3, 
        Multiplier_0_pp_1_4, Multiplier_0_pp_1_3, co_Multiplier_0_0_3, 
        Multiplier_0_pp_0_6, Multiplier_0_pp_0_5, Multiplier_0_pp_1_6, 
        Multiplier_0_pp_1_5, co_Multiplier_0_0_4, Multiplier_0_pp_0_8, 
        Multiplier_0_pp_0_7, Multiplier_0_pp_1_8, Multiplier_0_pp_1_7, 
        co_Multiplier_0_0_5, Multiplier_0_pp_0_10, Multiplier_0_pp_0_9, 
        Multiplier_0_pp_1_10, Multiplier_0_pp_1_9, co_Multiplier_0_0_6, 
        Multiplier_0_pp_0_12, Multiplier_0_pp_0_11, Multiplier_0_pp_1_12, 
        Multiplier_0_pp_1_11, co_Multiplier_0_0_7, Multiplier_0_pp_1_14, 
        Multiplier_0_pp_1_13, co_Multiplier_0_0_8, co_Multiplier_0_1_1, 
        Multiplier_0_pp_2_6, co_Multiplier_0_1_2, Multiplier_0_pp_2_8, 
        Multiplier_0_pp_2_7, Multiplier_0_pp_3_8, Multiplier_0_pp_3_7, 
        co_Multiplier_0_1_3, Multiplier_0_pp_2_10, Multiplier_0_pp_2_9, 
        Multiplier_0_pp_3_10, Multiplier_0_pp_3_9, co_Multiplier_0_1_4, 
        Multiplier_0_pp_2_12, Multiplier_0_pp_2_11, Multiplier_0_pp_3_12, 
        Multiplier_0_pp_3_11, co_Multiplier_0_1_5, Multiplier_0_pp_2_14, 
        Multiplier_0_pp_2_13, Multiplier_0_pp_3_14, Multiplier_0_pp_3_13, 
        co_Multiplier_0_1_6, Multiplier_0_pp_2_16, Multiplier_0_pp_2_15, 
        Multiplier_0_pp_3_16, Multiplier_0_pp_3_15, co_Multiplier_0_1_7, 
        Multiplier_0_pp_3_18, Multiplier_0_pp_3_17, co_Multiplier_0_1_8, 
        co_Multiplier_0_2_1, Multiplier_0_pp_4_10, co_Multiplier_0_2_2, 
        Multiplier_0_pp_4_12, Multiplier_0_pp_4_11, Multiplier_0_pp_5_12, 
        Multiplier_0_pp_5_11, co_Multiplier_0_2_3, Multiplier_0_pp_4_14, 
        Multiplier_0_pp_4_13, Multiplier_0_pp_5_14, Multiplier_0_pp_5_13, 
        co_Multiplier_0_2_4, Multiplier_0_pp_4_16, Multiplier_0_pp_4_15, 
        Multiplier_0_pp_5_16, Multiplier_0_pp_5_15, co_Multiplier_0_2_5, 
        Multiplier_0_pp_4_18, Multiplier_0_pp_4_17, Multiplier_0_pp_5_18, 
        Multiplier_0_pp_5_17, co_Multiplier_0_2_6, Multiplier_0_pp_4_20, 
        Multiplier_0_pp_4_19, Multiplier_0_pp_5_20, Multiplier_0_pp_5_19, 
        co_Multiplier_0_2_7, Multiplier_0_pp_5_22, Multiplier_0_pp_5_21, 
        co_Multiplier_0_3_1, co_Multiplier_0_3_2, co_Multiplier_0_3_3, 
        s_Multiplier_0_3_8, co_Multiplier_0_3_4, s_Multiplier_0_3_9, s_Multiplier_0_3_10, 
        co_Multiplier_0_3_5, s_Multiplier_0_3_11, s_Multiplier_0_3_12, 
        co_Multiplier_0_3_6, s_Multiplier_0_3_13, s_Multiplier_0_3_14, 
        co_Multiplier_0_3_7, s_Multiplier_0_3_15, s_Multiplier_0_3_16, 
        co_Multiplier_0_3_8, s_Multiplier_0_3_17, s_Multiplier_0_3_18, 
        co_Multiplier_0_3_9, s_Multiplier_0_3_19, s_Multiplier_0_3_20, 
        co_Multiplier_0_3_10, s_Multiplier_0_3_21, s_Multiplier_0_3_22, 
        s_Multiplier_0_3_23, co_t_Multiplier_0_4_1, co_t_Multiplier_0_4_2, 
        co_t_Multiplier_0_4_3, co_t_Multiplier_0_4_4, co_t_Multiplier_0_4_5, 
        co_t_Multiplier_0_4_6, co_t_Multiplier_0_4_7, co_t_Multiplier_0_4_8, 
        mco, mco_1, mco_2, mco_3, mco_4, Multiplier_0_mult_0_5_n2, 
        mco_5, mco_6, mco_7, mco_8, mco_9, Multiplier_0_mult_2_5_n2, 
        mco_10, mco_11, mco_12, mco_13, mco_14, Multiplier_0_mult_4_5_n2, 
        mco_15, mco_16, mco_17, mco_18, mco_19, Multiplier_0_mult_6_5_n2, 
        mco_20, mco_21, mco_22, mco_23, mco_24, Multiplier_0_mult_8_5_n2, 
        Multiplier_0_mult_10_0_n1, mco_25, mco_26, mco_27, mco_28, 
        mco_29;
    
    ND2 ND2_t25 (.A(rega_a_11), .B(regb_b_1), .Z(Multiplier_0_mult_0_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    AND2 AND2_t24 (.A(regb_b_0), .B(regb_b_2), .Z(Multiplier_0_pp_1_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(382[10:72])
    ND2 ND2_t22 (.A(rega_a_11), .B(regb_b_3), .Z(Multiplier_0_mult_2_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    AND2 AND2_t21 (.A(regb_b_0), .B(regb_b_4), .Z(Multiplier_0_pp_2_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(388[10:72])
    ND2 ND2_t19 (.A(rega_a_11), .B(regb_b_5), .Z(Multiplier_0_mult_4_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    AND2 AND2_t18 (.A(regb_b_0), .B(regb_b_6), .Z(Multiplier_0_pp_3_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(394[10:72])
    ND2 ND2_t16 (.A(rega_a_11), .B(regb_b_7), .Z(Multiplier_0_mult_6_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    AND2 AND2_t15 (.A(regb_b_0), .B(regb_b_8), .Z(Multiplier_0_pp_4_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(400[10:72])
    ND2 ND2_t13 (.A(rega_a_11), .B(regb_b_9), .Z(Multiplier_0_mult_8_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    AND2 AND2_t12 (.A(regb_b_0), .B(regb_b_10), .Z(Multiplier_0_pp_5_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(406[10:74])
    ND2 ND2_t10 (.A(regb_b_0), .B(regb_b_11), .Z(Multiplier_0_mult_10_0_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t9 (.A(rega_a_3), .B(regb_b_11), .Z(Multiplier_0_mult_10_1_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t8 (.A(rega_a_2), .B(regb_b_11), .Z(Multiplier_0_mult_10_1_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t7 (.A(rega_a_5), .B(regb_b_11), .Z(Multiplier_0_mult_10_2_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t6 (.A(rega_a_4), .B(regb_b_11), .Z(Multiplier_0_mult_10_2_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t5 (.A(rega_a_7), .B(regb_b_11), .Z(Multiplier_0_mult_10_3_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t4 (.A(rega_a_6), .B(regb_b_11), .Z(Multiplier_0_mult_10_3_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t3 (.A(rega_a_9), .B(regb_b_11), .Z(Multiplier_0_mult_10_4_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t2 (.A(rega_a_8), .B(regb_b_11), .Z(Multiplier_0_mult_10_4_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t1 (.A(rega_a_11), .B(regb_b_10), .Z(Multiplier_0_mult_10_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t0 (.A(rega_a_10), .B(regb_b_11), .Z(Multiplier_0_mult_10_5_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FD1P3DX FF_98 (.D(MultDataC[1]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(435[13:82])
    defparam FF_98.GSR = "ENABLED";
    FD1P3DX FF_97 (.D(MultDataC[2]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(438[13:82])
    defparam FF_97.GSR = "ENABLED";
    FD1P3DX FF_96 (.D(MultDataC[3]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(441[13:82])
    defparam FF_96.GSR = "ENABLED";
    FD1P3DX FF_95 (.D(MultDataC[4]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(444[13:82])
    defparam FF_95.GSR = "ENABLED";
    FD1P3DX FF_94 (.D(MultDataC[5]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(447[13:82])
    defparam FF_94.GSR = "ENABLED";
    FD1P3DX FF_93 (.D(MultDataC[6]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(450[13:82])
    defparam FF_93.GSR = "ENABLED";
    FD1P3DX FF_92 (.D(MultDataC[7]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(453[13:82])
    defparam FF_92.GSR = "ENABLED";
    FD1P3DX FF_91 (.D(MultDataC[8]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(456[13:82])
    defparam FF_91.GSR = "ENABLED";
    FD1P3DX FF_90 (.D(MultDataC[9]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(459[13:82])
    defparam FF_90.GSR = "ENABLED";
    FD1P3DX FF_89 (.D(MultDataC[10]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(462[13:84])
    defparam FF_89.GSR = "ENABLED";
    FD1P3DX FF_88 (.D(MultDataC[11]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(465[13:84])
    defparam FF_88.GSR = "ENABLED";
    FD1P3DX FF_87 (.D(MultDataC[0]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_0)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(468[13:82])
    defparam FF_87.GSR = "ENABLED";
    FD1P3DX FF_86 (.D(MultDataC[1]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(471[13:82])
    defparam FF_86.GSR = "ENABLED";
    FD1P3DX FF_85 (.D(MultDataC[2]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(474[13:82])
    defparam FF_85.GSR = "ENABLED";
    FD1P3DX FF_84 (.D(MultDataC[3]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(477[13:82])
    defparam FF_84.GSR = "ENABLED";
    FD1P3DX FF_83 (.D(MultDataC[4]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(480[13:82])
    defparam FF_83.GSR = "ENABLED";
    FD1P3DX FF_82 (.D(MultDataC[5]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(483[13:82])
    defparam FF_82.GSR = "ENABLED";
    FD1P3DX FF_81 (.D(MultDataC[6]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(486[13:82])
    defparam FF_81.GSR = "ENABLED";
    FD1P3DX FF_80 (.D(MultDataC[7]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(489[13:82])
    defparam FF_80.GSR = "ENABLED";
    FD1P3DX FF_79 (.D(MultDataC[8]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(492[13:82])
    defparam FF_79.GSR = "ENABLED";
    FD1P3DX FF_78 (.D(MultDataC[9]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(495[13:82])
    defparam FF_78.GSR = "ENABLED";
    FD1P3DX FF_77 (.D(MultDataC[10]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(498[13:84])
    defparam FF_77.GSR = "ENABLED";
    FD1P3DX FF_76 (.D(MultDataC[11]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(501[13:84])
    defparam FF_76.GSR = "ENABLED";
    FD1P3DX FF_75 (.D(rego_o_0), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[0])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(504[13:83])
    defparam FF_75.GSR = "ENABLED";
    FD1P3DX FF_74 (.D(rego_o_1), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[1])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(507[13:83])
    defparam FF_74.GSR = "ENABLED";
    FD1P3DX FF_73 (.D(rego_o_2), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[2])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(510[13:83])
    defparam FF_73.GSR = "ENABLED";
    FD1P3DX FF_72 (.D(rego_o_3), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[3])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(513[13:83])
    defparam FF_72.GSR = "ENABLED";
    FD1P3DX FF_71 (.D(rego_o_4), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[4])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(516[13:83])
    defparam FF_71.GSR = "ENABLED";
    FD1P3DX FF_70 (.D(rego_o_5), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[5])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(519[13:83])
    defparam FF_70.GSR = "ENABLED";
    FD1P3DX FF_69 (.D(rego_o_6), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[6])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(522[13:83])
    defparam FF_69.GSR = "ENABLED";
    FD1P3DX FF_68 (.D(rego_o_7), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[7])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(525[13:83])
    defparam FF_68.GSR = "ENABLED";
    FD1P3DX FF_67 (.D(rego_o_8), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[8])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(528[13:83])
    defparam FF_67.GSR = "ENABLED";
    FD1P3DX FF_66 (.D(rego_o_9), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult2[9])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(531[13:83])
    defparam FF_66.GSR = "ENABLED";
    FD1P3DX FF_65 (.D(rego_o_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[10])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(534[13:85])
    defparam FF_65.GSR = "ENABLED";
    FD1P3DX FF_64 (.D(rego_o_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[11])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(537[13:85])
    defparam FF_64.GSR = "ENABLED";
    FD1P3DX FF_63 (.D(rego_o_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[12])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(540[13:85])
    defparam FF_63.GSR = "ENABLED";
    FD1P3DX FF_62 (.D(rego_o_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[13])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(543[13:85])
    defparam FF_62.GSR = "ENABLED";
    FD1P3DX FF_61 (.D(rego_o_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[14])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(546[13:85])
    defparam FF_61.GSR = "ENABLED";
    FD1P3DX FF_60 (.D(rego_o_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[15])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(549[13:85])
    defparam FF_60.GSR = "ENABLED";
    FD1P3DX FF_59 (.D(rego_o_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[16])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(552[13:85])
    defparam FF_59.GSR = "ENABLED";
    FD1P3DX FF_58 (.D(rego_o_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[17])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(555[13:85])
    defparam FF_58.GSR = "ENABLED";
    FD1P3DX FF_57 (.D(rego_o_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[18])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(558[13:85])
    defparam FF_57.GSR = "ENABLED";
    FD1P3DX FF_56 (.D(rego_o_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[19])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(561[13:85])
    defparam FF_56.GSR = "ENABLED";
    FD1P3DX FF_55 (.D(rego_o_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[20])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(564[13:85])
    defparam FF_55.GSR = "ENABLED";
    FD1P3DX FF_54 (.D(rego_o_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[21])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(567[13:85])
    defparam FF_54.GSR = "ENABLED";
    FD1P3DX FF_53 (.D(rego_o_22), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[22])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(570[13:85])
    defparam FF_53.GSR = "ENABLED";
    FD1P3DX FF_52 (.D(rego_o_23), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult2[23])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(573[13:85])
    defparam FF_52.GSR = "ENABLED";
    FD1P3DX FF_51 (.D(Multiplier_0_pp_0_0), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_0)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(576[13] 577[35])
    defparam FF_51.GSR = "ENABLED";
    FD1P3DX FF_50 (.D(Multiplier_0_pp_0_1), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(580[13] 581[35])
    defparam FF_50.GSR = "ENABLED";
    FD1P3DX FF_49 (.D(s_Multiplier_0_0_2), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(584[13] 585[34])
    defparam FF_49.GSR = "ENABLED";
    FD1P3DX FF_48 (.D(s_Multiplier_0_0_3), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(588[13] 589[34])
    defparam FF_48.GSR = "ENABLED";
    FD1P3DX FF_47 (.D(s_Multiplier_0_0_4), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(592[13] 593[34])
    defparam FF_47.GSR = "ENABLED";
    FD1P3DX FF_46 (.D(s_Multiplier_0_0_5), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(596[13] 597[34])
    defparam FF_46.GSR = "ENABLED";
    FD1P3DX FF_45 (.D(s_Multiplier_0_0_6), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(600[13] 601[34])
    defparam FF_45.GSR = "ENABLED";
    FD1P3DX FF_44 (.D(s_Multiplier_0_0_7), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(604[13] 605[34])
    defparam FF_44.GSR = "ENABLED";
    FD1P3DX FF_43 (.D(s_Multiplier_0_0_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(608[13] 609[34])
    defparam FF_43.GSR = "ENABLED";
    FD1P3DX FF_42 (.D(s_Multiplier_0_0_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(612[13] 613[34])
    defparam FF_42.GSR = "ENABLED";
    FD1P3DX FF_41 (.D(s_Multiplier_0_0_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(616[13] 617[35])
    defparam FF_41.GSR = "ENABLED";
    FD1P3DX FF_40 (.D(s_Multiplier_0_0_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(620[13] 621[35])
    defparam FF_40.GSR = "ENABLED";
    FD1P3DX FF_39 (.D(s_Multiplier_0_0_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(624[13] 625[35])
    defparam FF_39.GSR = "ENABLED";
    FD1P3DX FF_38 (.D(s_Multiplier_0_0_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(628[13] 629[35])
    defparam FF_38.GSR = "ENABLED";
    FD1P3DX FF_37 (.D(s_Multiplier_0_0_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(632[13] 633[35])
    defparam FF_37.GSR = "ENABLED";
    FD1P3DX FF_36 (.D(s_Multiplier_0_0_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(636[13] 637[35])
    defparam FF_36.GSR = "ENABLED";
    FD1P3DX FF_35 (.D(s_Multiplier_0_0_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(640[13] 641[35])
    defparam FF_35.GSR = "ENABLED";
    FD1P3DX FF_34 (.D(s_Multiplier_0_0_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(644[13] 645[35])
    defparam FF_34.GSR = "ENABLED";
    FD1P3DX FF_33 (.D(Multiplier_0_pp_2_4), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_2_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(648[13] 649[35])
    defparam FF_33.GSR = "ENABLED";
    FD1P3DX FF_32 (.D(Multiplier_0_pp_2_5), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_2_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(652[13] 653[35])
    defparam FF_32.GSR = "ENABLED";
    FD1P3DX FF_31 (.D(s_Multiplier_0_1_6), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(656[13] 657[34])
    defparam FF_31.GSR = "ENABLED";
    FD1P3DX FF_30 (.D(s_Multiplier_0_1_7), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(660[13] 661[34])
    defparam FF_30.GSR = "ENABLED";
    FD1P3DX FF_29 (.D(s_Multiplier_0_1_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(664[13] 665[34])
    defparam FF_29.GSR = "ENABLED";
    FD1P3DX FF_28 (.D(s_Multiplier_0_1_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(668[13] 669[34])
    defparam FF_28.GSR = "ENABLED";
    FD1P3DX FF_27 (.D(s_Multiplier_0_1_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(672[13] 673[35])
    defparam FF_27.GSR = "ENABLED";
    FD1P3DX FF_26 (.D(s_Multiplier_0_1_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(676[13] 677[35])
    defparam FF_26.GSR = "ENABLED";
    FD1P3DX FF_25 (.D(s_Multiplier_0_1_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(680[13] 681[35])
    defparam FF_25.GSR = "ENABLED";
    FD1P3DX FF_24 (.D(s_Multiplier_0_1_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(684[13] 685[35])
    defparam FF_24.GSR = "ENABLED";
    FD1P3DX FF_23 (.D(s_Multiplier_0_1_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(688[13] 689[35])
    defparam FF_23.GSR = "ENABLED";
    FD1P3DX FF_22 (.D(s_Multiplier_0_1_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(692[13] 693[35])
    defparam FF_22.GSR = "ENABLED";
    FD1P3DX FF_21 (.D(s_Multiplier_0_1_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(696[13] 697[35])
    defparam FF_21.GSR = "ENABLED";
    FD1P3DX FF_20 (.D(s_Multiplier_0_1_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(700[13] 701[35])
    defparam FF_20.GSR = "ENABLED";
    FD1P3DX FF_19 (.D(s_Multiplier_0_1_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(704[13] 705[35])
    defparam FF_19.GSR = "ENABLED";
    FD1P3DX FF_18 (.D(s_Multiplier_0_1_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(708[13] 709[35])
    defparam FF_18.GSR = "ENABLED";
    FD1P3DX FF_17 (.D(s_Multiplier_0_1_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(712[13] 713[35])
    defparam FF_17.GSR = "ENABLED";
    FD1P3DX FF_16 (.D(s_Multiplier_0_1_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(716[13] 717[35])
    defparam FF_16.GSR = "ENABLED";
    FD1P3DX FF_15 (.D(Multiplier_0_pp_4_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_4_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(720[13] 721[35])
    defparam FF_15.GSR = "ENABLED";
    FD1P3DX FF_14 (.D(Multiplier_0_pp_4_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_4_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(724[13] 725[35])
    defparam FF_14.GSR = "ENABLED";
    FD1P3DX FF_13 (.D(s_Multiplier_0_2_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(728[13] 729[35])
    defparam FF_13.GSR = "ENABLED";
    FD1P3DX FF_12 (.D(s_Multiplier_0_2_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(732[13] 733[35])
    defparam FF_12.GSR = "ENABLED";
    FD1P3DX FF_11 (.D(s_Multiplier_0_2_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(736[13] 737[35])
    defparam FF_11.GSR = "ENABLED";
    FD1P3DX FF_10 (.D(s_Multiplier_0_2_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(740[13] 741[35])
    defparam FF_10.GSR = "ENABLED";
    FD1P3DX FF_9 (.D(s_Multiplier_0_2_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(744[13] 745[35])
    defparam FF_9.GSR = "ENABLED";
    FD1P3DX FF_8 (.D(s_Multiplier_0_2_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(748[13] 749[35])
    defparam FF_8.GSR = "ENABLED";
    FD1P3DX FF_7 (.D(s_Multiplier_0_2_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(752[13] 753[35])
    defparam FF_7.GSR = "ENABLED";
    FD1P3DX FF_6 (.D(s_Multiplier_0_2_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(756[13] 757[35])
    defparam FF_6.GSR = "ENABLED";
    FD1P3DX FF_5 (.D(s_Multiplier_0_2_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(760[13] 761[35])
    defparam FF_5.GSR = "ENABLED";
    FD1P3DX FF_4 (.D(s_Multiplier_0_2_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(764[13] 765[35])
    defparam FF_4.GSR = "ENABLED";
    FD1P3DX FF_3 (.D(s_Multiplier_0_2_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(768[13] 769[35])
    defparam FF_3.GSR = "ENABLED";
    FD1P3DX FF_2 (.D(s_Multiplier_0_2_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(772[13] 773[35])
    defparam FF_2.GSR = "ENABLED";
    FD1P3DX FF_1 (.D(s_Multiplier_0_2_22), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_22)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(776[13] 777[35])
    defparam FF_1.GSR = "ENABLED";
    FD1P3DX FF_0 (.D(s_Multiplier_0_2_23), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_23)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(780[13] 781[35])
    defparam FF_0.GSR = "ENABLED";
    FADD2B Multiplier_0_cin_lr_add_0 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_Cadd_0_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco), .S0(Multiplier_0_pp_0_13)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_cin_lr_add_2 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_Cadd_2_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_1), .S0(Multiplier_0_pp_1_15)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_cin_lr_add_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_Cadd_4_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_2), .S0(Multiplier_0_pp_2_17)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_cin_lr_add_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_Cadd_6_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_3), .S0(Multiplier_0_pp_3_19)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_cin_lr_add_8 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_Cadd_8_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_4), .S0(Multiplier_0_pp_4_21)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_cin_lr_add_10 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_Cadd_10_6 (.A0(VCC_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_5), .S0(Multiplier_0_pp_5_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_Multiplier_0_0_1 (.A0(GND_net), .A1(Multiplier_0_pp_0_2), 
           .B0(GND_net), .B1(Multiplier_0_pp_1_2), .CI(GND_net), .COUT(co_Multiplier_0_0_1), 
           .S1(s_Multiplier_0_0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_0_2 (.A0(Multiplier_0_pp_0_3), .A1(Multiplier_0_pp_0_4), 
           .B0(Multiplier_0_pp_1_3), .B1(Multiplier_0_pp_1_4), .CI(co_Multiplier_0_0_1), 
           .COUT(co_Multiplier_0_0_2), .S0(s_Multiplier_0_0_3), .S1(s_Multiplier_0_0_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_0_3 (.A0(Multiplier_0_pp_0_5), .A1(Multiplier_0_pp_0_6), 
           .B0(Multiplier_0_pp_1_5), .B1(Multiplier_0_pp_1_6), .CI(co_Multiplier_0_0_2), 
           .COUT(co_Multiplier_0_0_3), .S0(s_Multiplier_0_0_5), .S1(s_Multiplier_0_0_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_0_4 (.A0(Multiplier_0_pp_0_7), .A1(Multiplier_0_pp_0_8), 
           .B0(Multiplier_0_pp_1_7), .B1(Multiplier_0_pp_1_8), .CI(co_Multiplier_0_0_3), 
           .COUT(co_Multiplier_0_0_4), .S0(s_Multiplier_0_0_7), .S1(s_Multiplier_0_0_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_0_5 (.A0(Multiplier_0_pp_0_9), .A1(Multiplier_0_pp_0_10), 
           .B0(Multiplier_0_pp_1_9), .B1(Multiplier_0_pp_1_10), .CI(co_Multiplier_0_0_4), 
           .COUT(co_Multiplier_0_0_5), .S0(s_Multiplier_0_0_9), .S1(s_Multiplier_0_0_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_0_6 (.A0(Multiplier_0_pp_0_11), .A1(Multiplier_0_pp_0_12), 
           .B0(Multiplier_0_pp_1_11), .B1(Multiplier_0_pp_1_12), .CI(co_Multiplier_0_0_5), 
           .COUT(co_Multiplier_0_0_6), .S0(s_Multiplier_0_0_11), .S1(s_Multiplier_0_0_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_0_7 (.A0(Multiplier_0_pp_0_13), .A1(GND_net), 
           .B0(Multiplier_0_pp_1_13), .B1(Multiplier_0_pp_1_14), .CI(co_Multiplier_0_0_6), 
           .COUT(co_Multiplier_0_0_7), .S0(s_Multiplier_0_0_13), .S1(s_Multiplier_0_0_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_0_8 (.A0(GND_net), .A1(GND_net), .B0(Multiplier_0_pp_1_15), 
           .B1(GND_net), .CI(co_Multiplier_0_0_7), .COUT(co_Multiplier_0_0_8), 
           .S0(s_Multiplier_0_0_15), .S1(s_Multiplier_0_0_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_Multiplier_0_0_9 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_Multiplier_0_0_8), .S0(s_Multiplier_0_0_17)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_Multiplier_0_1_1 (.A0(GND_net), .A1(Multiplier_0_pp_2_6), 
           .B0(GND_net), .B1(Multiplier_0_pp_3_6), .CI(GND_net), .COUT(co_Multiplier_0_1_1), 
           .S1(s_Multiplier_0_1_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_1_2 (.A0(Multiplier_0_pp_2_7), .A1(Multiplier_0_pp_2_8), 
           .B0(Multiplier_0_pp_3_7), .B1(Multiplier_0_pp_3_8), .CI(co_Multiplier_0_1_1), 
           .COUT(co_Multiplier_0_1_2), .S0(s_Multiplier_0_1_7), .S1(s_Multiplier_0_1_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_1_3 (.A0(Multiplier_0_pp_2_9), .A1(Multiplier_0_pp_2_10), 
           .B0(Multiplier_0_pp_3_9), .B1(Multiplier_0_pp_3_10), .CI(co_Multiplier_0_1_2), 
           .COUT(co_Multiplier_0_1_3), .S0(s_Multiplier_0_1_9), .S1(s_Multiplier_0_1_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_1_4 (.A0(Multiplier_0_pp_2_11), .A1(Multiplier_0_pp_2_12), 
           .B0(Multiplier_0_pp_3_11), .B1(Multiplier_0_pp_3_12), .CI(co_Multiplier_0_1_3), 
           .COUT(co_Multiplier_0_1_4), .S0(s_Multiplier_0_1_11), .S1(s_Multiplier_0_1_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_1_5 (.A0(Multiplier_0_pp_2_13), .A1(Multiplier_0_pp_2_14), 
           .B0(Multiplier_0_pp_3_13), .B1(Multiplier_0_pp_3_14), .CI(co_Multiplier_0_1_4), 
           .COUT(co_Multiplier_0_1_5), .S0(s_Multiplier_0_1_13), .S1(s_Multiplier_0_1_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_1_6 (.A0(Multiplier_0_pp_2_15), .A1(Multiplier_0_pp_2_16), 
           .B0(Multiplier_0_pp_3_15), .B1(Multiplier_0_pp_3_16), .CI(co_Multiplier_0_1_5), 
           .COUT(co_Multiplier_0_1_6), .S0(s_Multiplier_0_1_15), .S1(s_Multiplier_0_1_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_1_7 (.A0(Multiplier_0_pp_2_17), .A1(GND_net), 
           .B0(Multiplier_0_pp_3_17), .B1(Multiplier_0_pp_3_18), .CI(co_Multiplier_0_1_6), 
           .COUT(co_Multiplier_0_1_7), .S0(s_Multiplier_0_1_17), .S1(s_Multiplier_0_1_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_1_8 (.A0(GND_net), .A1(GND_net), .B0(Multiplier_0_pp_3_19), 
           .B1(GND_net), .CI(co_Multiplier_0_1_7), .COUT(co_Multiplier_0_1_8), 
           .S0(s_Multiplier_0_1_19), .S1(s_Multiplier_0_1_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_Multiplier_0_1_9 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_Multiplier_0_1_8), .S0(s_Multiplier_0_1_21)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_Multiplier_0_2_1 (.A0(GND_net), .A1(Multiplier_0_pp_4_10), 
           .B0(GND_net), .B1(Multiplier_0_pp_5_10), .CI(GND_net), .COUT(co_Multiplier_0_2_1), 
           .S1(s_Multiplier_0_2_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_2_2 (.A0(Multiplier_0_pp_4_11), .A1(Multiplier_0_pp_4_12), 
           .B0(Multiplier_0_pp_5_11), .B1(Multiplier_0_pp_5_12), .CI(co_Multiplier_0_2_1), 
           .COUT(co_Multiplier_0_2_2), .S0(s_Multiplier_0_2_11), .S1(s_Multiplier_0_2_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_2_3 (.A0(Multiplier_0_pp_4_13), .A1(Multiplier_0_pp_4_14), 
           .B0(Multiplier_0_pp_5_13), .B1(Multiplier_0_pp_5_14), .CI(co_Multiplier_0_2_2), 
           .COUT(co_Multiplier_0_2_3), .S0(s_Multiplier_0_2_13), .S1(s_Multiplier_0_2_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_2_4 (.A0(Multiplier_0_pp_4_15), .A1(Multiplier_0_pp_4_16), 
           .B0(Multiplier_0_pp_5_15), .B1(Multiplier_0_pp_5_16), .CI(co_Multiplier_0_2_3), 
           .COUT(co_Multiplier_0_2_4), .S0(s_Multiplier_0_2_15), .S1(s_Multiplier_0_2_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_2_5 (.A0(Multiplier_0_pp_4_17), .A1(Multiplier_0_pp_4_18), 
           .B0(Multiplier_0_pp_5_17), .B1(Multiplier_0_pp_5_18), .CI(co_Multiplier_0_2_4), 
           .COUT(co_Multiplier_0_2_5), .S0(s_Multiplier_0_2_17), .S1(s_Multiplier_0_2_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_2_6 (.A0(Multiplier_0_pp_4_19), .A1(Multiplier_0_pp_4_20), 
           .B0(Multiplier_0_pp_5_19), .B1(Multiplier_0_pp_5_20), .CI(co_Multiplier_0_2_5), 
           .COUT(co_Multiplier_0_2_6), .S0(s_Multiplier_0_2_19), .S1(s_Multiplier_0_2_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_2_7 (.A0(Multiplier_0_pp_4_21), .A1(GND_net), 
           .B0(Multiplier_0_pp_5_21), .B1(Multiplier_0_pp_5_22), .CI(co_Multiplier_0_2_6), 
           .COUT(co_Multiplier_0_2_7), .S0(s_Multiplier_0_2_21), .S1(s_Multiplier_0_2_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_2_8 (.A0(GND_net), .A1(GND_net), .B0(Multiplier_0_pp_5_23), 
           .B1(GND_net), .CI(co_Multiplier_0_2_7), .S0(s_Multiplier_0_2_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_Multiplier_0_3_1 (.A0(GND_net), .A1(f_s_Multiplier_0_0_4), 
           .B0(GND_net), .B1(f_Multiplier_0_pp_2_4), .CI(GND_net), .COUT(co_Multiplier_0_3_1), 
           .S1(rego_o_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_2 (.A0(f_s_Multiplier_0_0_5), .A1(f_s_Multiplier_0_0_6), 
           .B0(f_Multiplier_0_pp_2_5), .B1(f_s_Multiplier_0_1_6), .CI(co_Multiplier_0_3_1), 
           .COUT(co_Multiplier_0_3_2), .S0(rego_o_5), .S1(rego_o_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_3 (.A0(f_s_Multiplier_0_0_7), .A1(f_s_Multiplier_0_0_8), 
           .B0(f_s_Multiplier_0_1_7), .B1(f_s_Multiplier_0_1_8), .CI(co_Multiplier_0_3_2), 
           .COUT(co_Multiplier_0_3_3), .S0(rego_o_7), .S1(s_Multiplier_0_3_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_4 (.A0(f_s_Multiplier_0_0_9), .A1(f_s_Multiplier_0_0_10), 
           .B0(f_s_Multiplier_0_1_9), .B1(f_s_Multiplier_0_1_10), .CI(co_Multiplier_0_3_3), 
           .COUT(co_Multiplier_0_3_4), .S0(s_Multiplier_0_3_9), .S1(s_Multiplier_0_3_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_5 (.A0(f_s_Multiplier_0_0_11), .A1(f_s_Multiplier_0_0_12), 
           .B0(f_s_Multiplier_0_1_11), .B1(f_s_Multiplier_0_1_12), .CI(co_Multiplier_0_3_4), 
           .COUT(co_Multiplier_0_3_5), .S0(s_Multiplier_0_3_11), .S1(s_Multiplier_0_3_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_6 (.A0(f_s_Multiplier_0_0_13), .A1(f_s_Multiplier_0_0_14), 
           .B0(f_s_Multiplier_0_1_13), .B1(f_s_Multiplier_0_1_14), .CI(co_Multiplier_0_3_5), 
           .COUT(co_Multiplier_0_3_6), .S0(s_Multiplier_0_3_13), .S1(s_Multiplier_0_3_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_7 (.A0(f_s_Multiplier_0_0_15), .A1(f_s_Multiplier_0_0_16), 
           .B0(f_s_Multiplier_0_1_15), .B1(f_s_Multiplier_0_1_16), .CI(co_Multiplier_0_3_6), 
           .COUT(co_Multiplier_0_3_7), .S0(s_Multiplier_0_3_15), .S1(s_Multiplier_0_3_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_8 (.A0(f_s_Multiplier_0_0_17), .A1(GND_net), 
           .B0(f_s_Multiplier_0_1_17), .B1(f_s_Multiplier_0_1_18), .CI(co_Multiplier_0_3_7), 
           .COUT(co_Multiplier_0_3_8), .S0(s_Multiplier_0_3_17), .S1(s_Multiplier_0_3_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_9 (.A0(GND_net), .A1(GND_net), .B0(f_s_Multiplier_0_1_19), 
           .B1(f_s_Multiplier_0_1_20), .CI(co_Multiplier_0_3_8), .COUT(co_Multiplier_0_3_9), 
           .S0(s_Multiplier_0_3_19), .S1(s_Multiplier_0_3_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Multiplier_0_add_3_10 (.A0(GND_net), .A1(GND_net), .B0(f_s_Multiplier_0_1_21), 
           .B1(GND_net), .CI(co_Multiplier_0_3_9), .COUT(co_Multiplier_0_3_10), 
           .S0(s_Multiplier_0_3_21), .S1(s_Multiplier_0_3_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_Multiplier_0_3_11 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_Multiplier_0_3_10), .S0(s_Multiplier_0_3_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B Cadd_t_Multiplier_0_4_1 (.A0(GND_net), .A1(s_Multiplier_0_3_8), 
           .B0(GND_net), .B1(f_Multiplier_0_pp_4_8), .CI(GND_net), .COUT(co_t_Multiplier_0_4_1), 
           .S1(rego_o_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_2 (.A0(s_Multiplier_0_3_9), .A1(s_Multiplier_0_3_10), 
           .B0(f_Multiplier_0_pp_4_9), .B1(f_s_Multiplier_0_2_10), .CI(co_t_Multiplier_0_4_1), 
           .COUT(co_t_Multiplier_0_4_2), .S0(rego_o_9), .S1(rego_o_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_3 (.A0(s_Multiplier_0_3_11), .A1(s_Multiplier_0_3_12), 
           .B0(f_s_Multiplier_0_2_11), .B1(f_s_Multiplier_0_2_12), .CI(co_t_Multiplier_0_4_2), 
           .COUT(co_t_Multiplier_0_4_3), .S0(rego_o_11), .S1(rego_o_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_4 (.A0(s_Multiplier_0_3_13), .A1(s_Multiplier_0_3_14), 
           .B0(f_s_Multiplier_0_2_13), .B1(f_s_Multiplier_0_2_14), .CI(co_t_Multiplier_0_4_3), 
           .COUT(co_t_Multiplier_0_4_4), .S0(rego_o_13), .S1(rego_o_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_5 (.A0(s_Multiplier_0_3_15), .A1(s_Multiplier_0_3_16), 
           .B0(f_s_Multiplier_0_2_15), .B1(f_s_Multiplier_0_2_16), .CI(co_t_Multiplier_0_4_4), 
           .COUT(co_t_Multiplier_0_4_5), .S0(rego_o_15), .S1(rego_o_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_6 (.A0(s_Multiplier_0_3_17), .A1(s_Multiplier_0_3_18), 
           .B0(f_s_Multiplier_0_2_17), .B1(f_s_Multiplier_0_2_18), .CI(co_t_Multiplier_0_4_5), 
           .COUT(co_t_Multiplier_0_4_6), .S0(rego_o_17), .S1(rego_o_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_7 (.A0(s_Multiplier_0_3_19), .A1(s_Multiplier_0_3_20), 
           .B0(f_s_Multiplier_0_2_19), .B1(f_s_Multiplier_0_2_20), .CI(co_t_Multiplier_0_4_6), 
           .COUT(co_t_Multiplier_0_4_7), .S0(rego_o_19), .S1(rego_o_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_8 (.A0(s_Multiplier_0_3_21), .A1(s_Multiplier_0_3_22), 
           .B0(f_s_Multiplier_0_2_21), .B1(f_s_Multiplier_0_2_22), .CI(co_t_Multiplier_0_4_7), 
           .COUT(co_t_Multiplier_0_4_8), .S0(rego_o_21), .S1(rego_o_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    FADD2B t_Multiplier_0_add_4_9 (.A0(s_Multiplier_0_3_23), .A1(GND_net), 
           .B0(f_s_Multiplier_0_2_23), .B1(GND_net), .CI(co_t_Multiplier_0_4_8), 
           .S0(rego_o_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_0_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(Multiplier_0_cin_lr_0), .CO(mco), .P0(Multiplier_0_pp_0_1), 
          .P1(Multiplier_0_pp_0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_0_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco), .CO(mco_1), .P0(Multiplier_0_pp_0_3), 
          .P1(Multiplier_0_pp_0_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_0_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco_1), .CO(mco_2), .P0(Multiplier_0_pp_0_5), 
          .P1(Multiplier_0_pp_0_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_0_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco_2), .CO(mco_3), .P0(Multiplier_0_pp_0_7), 
          .P1(Multiplier_0_pp_0_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_0_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco_3), .CO(mco_4), .P0(Multiplier_0_pp_0_9), 
          .P1(Multiplier_0_pp_0_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_0_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_0_5_n2), 
          .A2(Multiplier_0_mult_0_5_n1), .A3(VCC_net), .B0(regb_b_1), 
          .B1(VCC_net), .B2(VCC_net), .B3(VCC_net), .CI(mco_4), .CO(mfco), 
          .P0(Multiplier_0_pp_0_11), .P1(Multiplier_0_pp_0_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_2_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(Multiplier_0_cin_lr_2), .CO(mco_5), .P0(Multiplier_0_pp_1_3), 
          .P1(Multiplier_0_pp_1_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_2_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_5), .CO(mco_6), .P0(Multiplier_0_pp_1_5), 
          .P1(Multiplier_0_pp_1_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_2_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_6), .CO(mco_7), .P0(Multiplier_0_pp_1_7), 
          .P1(Multiplier_0_pp_1_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_2_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_7), .CO(mco_8), .P0(Multiplier_0_pp_1_9), 
          .P1(Multiplier_0_pp_1_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_2_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_8), .CO(mco_9), .P0(Multiplier_0_pp_1_11), 
          .P1(Multiplier_0_pp_1_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_2_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_2_5_n2), 
          .A2(Multiplier_0_mult_2_5_n1), .A3(GND_net), .B0(regb_b_3), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_2), .CI(mco_9), .CO(mfco_1), 
          .P0(Multiplier_0_pp_1_13), .P1(Multiplier_0_pp_1_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_4_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(Multiplier_0_cin_lr_4), .CO(mco_10), .P0(Multiplier_0_pp_2_5), 
          .P1(Multiplier_0_pp_2_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_4_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_10), .CO(mco_11), .P0(Multiplier_0_pp_2_7), 
          .P1(Multiplier_0_pp_2_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_4_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_11), .CO(mco_12), .P0(Multiplier_0_pp_2_9), 
          .P1(Multiplier_0_pp_2_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_4_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_12), .CO(mco_13), .P0(Multiplier_0_pp_2_11), 
          .P1(Multiplier_0_pp_2_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_4_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_13), .CO(mco_14), .P0(Multiplier_0_pp_2_13), 
          .P1(Multiplier_0_pp_2_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_4_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_4_5_n2), 
          .A2(Multiplier_0_mult_4_5_n1), .A3(GND_net), .B0(regb_b_5), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_4), .CI(mco_14), .CO(mfco_2), 
          .P0(Multiplier_0_pp_2_15), .P1(Multiplier_0_pp_2_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_6_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(Multiplier_0_cin_lr_6), .CO(mco_15), .P0(Multiplier_0_pp_3_7), 
          .P1(Multiplier_0_pp_3_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_6_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_15), .CO(mco_16), .P0(Multiplier_0_pp_3_9), 
          .P1(Multiplier_0_pp_3_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_6_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_16), .CO(mco_17), .P0(Multiplier_0_pp_3_11), 
          .P1(Multiplier_0_pp_3_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_6_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_17), .CO(mco_18), .P0(Multiplier_0_pp_3_13), 
          .P1(Multiplier_0_pp_3_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_6_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_18), .CO(mco_19), .P0(Multiplier_0_pp_3_15), 
          .P1(Multiplier_0_pp_3_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_6_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_6_5_n2), 
          .A2(Multiplier_0_mult_6_5_n1), .A3(GND_net), .B0(regb_b_7), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_6), .CI(mco_19), .CO(mfco_3), 
          .P0(Multiplier_0_pp_3_17), .P1(Multiplier_0_pp_3_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_8_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(Multiplier_0_cin_lr_8), .CO(mco_20), .P0(Multiplier_0_pp_4_9), 
          .P1(Multiplier_0_pp_4_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_8_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_20), .CO(mco_21), .P0(Multiplier_0_pp_4_11), 
          .P1(Multiplier_0_pp_4_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_8_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_21), .CO(mco_22), .P0(Multiplier_0_pp_4_13), 
          .P1(Multiplier_0_pp_4_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_8_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_22), .CO(mco_23), .P0(Multiplier_0_pp_4_15), 
          .P1(Multiplier_0_pp_4_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_8_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_23), .CO(mco_24), .P0(Multiplier_0_pp_4_17), 
          .P1(Multiplier_0_pp_4_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_8_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_8_5_n2), 
          .A2(Multiplier_0_mult_8_5_n1), .A3(GND_net), .B0(regb_b_9), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_8), .CI(mco_24), .CO(mfco_4), 
          .P0(Multiplier_0_pp_4_19), .P1(Multiplier_0_pp_4_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_10_0 (.A0(Multiplier_0_mult_10_0_n0), .A1(rega_a_1), 
          .A2(Multiplier_0_mult_10_0_n1), .A3(rega_a_2), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(Multiplier_0_cin_lr_10), 
          .CO(mco_25), .P0(Multiplier_0_pp_5_11), .P1(Multiplier_0_pp_5_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_10_1 (.A0(Multiplier_0_mult_10_1_n0), .A1(rega_a_3), 
          .A2(Multiplier_0_mult_10_1_n1), .A3(rega_a_4), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_25), 
          .CO(mco_26), .P0(Multiplier_0_pp_5_13), .P1(Multiplier_0_pp_5_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_10_2 (.A0(Multiplier_0_mult_10_2_n0), .A1(rega_a_5), 
          .A2(Multiplier_0_mult_10_2_n1), .A3(rega_a_6), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_26), 
          .CO(mco_27), .P0(Multiplier_0_pp_5_15), .P1(Multiplier_0_pp_5_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_10_3 (.A0(Multiplier_0_mult_10_3_n0), .A1(rega_a_7), 
          .A2(Multiplier_0_mult_10_3_n1), .A3(rega_a_8), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_27), 
          .CO(mco_28), .P0(Multiplier_0_pp_5_17), .P1(Multiplier_0_pp_5_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_10_4 (.A0(Multiplier_0_mult_10_4_n0), .A1(rega_a_9), 
          .A2(Multiplier_0_mult_10_4_n1), .A3(rega_a_10), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_28), 
          .CO(mco_29), .P0(Multiplier_0_pp_5_19), .P1(Multiplier_0_pp_5_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    MULT2 Multiplier_0_mult_10_5 (.A0(Multiplier_0_mult_10_5_n0), .A1(Multiplier_0_mult_10_5_n2), 
          .A2(rega_a_11), .A3(GND_net), .B0(VCC_net), .B1(VCC_net), 
          .B2(regb_b_11), .B3(regb_b_10), .CI(mco_29), .CO(mfco_5), 
          .P0(Multiplier_0_pp_5_21), .P1(Multiplier_0_pp_5_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    AND2 AND2_t27 (.A(regb_b_0), .B(regb_b_0), .Z(Multiplier_0_pp_0_0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(376[10:72])
    ND2 ND2_t26 (.A(rega_a_11), .B(regb_b_0), .Z(Multiplier_0_mult_0_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t23 (.A(rega_a_11), .B(regb_b_2), .Z(Multiplier_0_mult_2_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t20 (.A(rega_a_11), .B(regb_b_4), .Z(Multiplier_0_mult_4_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t17 (.A(rega_a_11), .B(regb_b_6), .Z(Multiplier_0_mult_6_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t14 (.A(rega_a_11), .B(regb_b_8), .Z(Multiplier_0_mult_8_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    ND2 ND2_t11 (.A(rega_a_1), .B(regb_b_11), .Z(Multiplier_0_mult_10_0_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=77, LSE_RLINE=83 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(77[14] 83[27])
    
endmodule
//
// Verilog Description of module Multiplier_U0
//

module Multiplier_U0 (CIC1_out_clkSin, VCC_net, GND_net, MultDataB, 
            MultResult1) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input CIC1_out_clkSin;
    input VCC_net;
    input GND_net;
    input [11:0]MultDataB;
    output [23:0]MultResult1;
    
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/impl1/source/top.v(67[6:21])
    
    wire Multiplier_0_mult_0_5_n1, regb_b_1, rega_a_11, Multiplier_0_pp_1_2, 
        regb_b_2, regb_b_0, Multiplier_0_mult_2_5_n1, regb_b_3, Multiplier_0_pp_2_4, 
        regb_b_4, Multiplier_0_mult_4_5_n1, regb_b_5, Multiplier_0_pp_3_6, 
        regb_b_6, Multiplier_0_mult_6_5_n1, regb_b_7, Multiplier_0_pp_4_8, 
        regb_b_8, Multiplier_0_mult_8_5_n1, regb_b_9, Multiplier_0_pp_5_10, 
        regb_b_10, Multiplier_0_mult_10_0_n0, regb_b_11, Multiplier_0_mult_10_1_n1, 
        rega_a_3, rega_a_2, Multiplier_0_mult_10_1_n0, Multiplier_0_mult_10_2_n1, 
        rega_a_5, rega_a_4, Multiplier_0_mult_10_2_n0, Multiplier_0_mult_10_3_n1, 
        rega_a_7, rega_a_6, Multiplier_0_mult_10_3_n0, Multiplier_0_mult_10_4_n1, 
        rega_a_9, rega_a_8, Multiplier_0_mult_10_4_n0, Multiplier_0_mult_10_5_n2, 
        rega_a_10, Multiplier_0_mult_10_5_n0, rega_a_1, rego_o_0, rego_o_1, 
        rego_o_2, rego_o_3, rego_o_4, rego_o_5, rego_o_6, rego_o_7, 
        rego_o_8, rego_o_9, rego_o_10, rego_o_11, rego_o_12, rego_o_13, 
        rego_o_14, rego_o_15, rego_o_16, rego_o_17, rego_o_18, rego_o_19, 
        rego_o_20, rego_o_21, rego_o_22, rego_o_23, Multiplier_0_pp_0_0, 
        Multiplier_0_pp_0_1, s_Multiplier_0_0_2, s_Multiplier_0_0_3, s_Multiplier_0_0_4, 
        f_s_Multiplier_0_0_4, s_Multiplier_0_0_5, f_s_Multiplier_0_0_5, 
        s_Multiplier_0_0_6, f_s_Multiplier_0_0_6, s_Multiplier_0_0_7, 
        f_s_Multiplier_0_0_7, s_Multiplier_0_0_8, f_s_Multiplier_0_0_8, 
        s_Multiplier_0_0_9, f_s_Multiplier_0_0_9, s_Multiplier_0_0_10, 
        f_s_Multiplier_0_0_10, s_Multiplier_0_0_11, f_s_Multiplier_0_0_11, 
        s_Multiplier_0_0_12, f_s_Multiplier_0_0_12, s_Multiplier_0_0_13, 
        f_s_Multiplier_0_0_13, s_Multiplier_0_0_14, f_s_Multiplier_0_0_14, 
        s_Multiplier_0_0_15, f_s_Multiplier_0_0_15, s_Multiplier_0_0_16, 
        f_s_Multiplier_0_0_16, s_Multiplier_0_0_17, f_s_Multiplier_0_0_17, 
        f_Multiplier_0_pp_2_4, f_Multiplier_0_pp_2_5, Multiplier_0_pp_2_5, 
        s_Multiplier_0_1_6, f_s_Multiplier_0_1_6, s_Multiplier_0_1_7, 
        f_s_Multiplier_0_1_7, s_Multiplier_0_1_8, f_s_Multiplier_0_1_8, 
        s_Multiplier_0_1_9, f_s_Multiplier_0_1_9, s_Multiplier_0_1_10, 
        f_s_Multiplier_0_1_10, s_Multiplier_0_1_11, f_s_Multiplier_0_1_11, 
        s_Multiplier_0_1_12, f_s_Multiplier_0_1_12, s_Multiplier_0_1_13, 
        f_s_Multiplier_0_1_13, s_Multiplier_0_1_14, f_s_Multiplier_0_1_14, 
        s_Multiplier_0_1_15, f_s_Multiplier_0_1_15, s_Multiplier_0_1_16, 
        f_s_Multiplier_0_1_16, s_Multiplier_0_1_17, f_s_Multiplier_0_1_17, 
        s_Multiplier_0_1_18, f_s_Multiplier_0_1_18, s_Multiplier_0_1_19, 
        f_s_Multiplier_0_1_19, s_Multiplier_0_1_20, f_s_Multiplier_0_1_20, 
        s_Multiplier_0_1_21, f_s_Multiplier_0_1_21, f_Multiplier_0_pp_4_8, 
        f_Multiplier_0_pp_4_9, Multiplier_0_pp_4_9, s_Multiplier_0_2_10, 
        f_s_Multiplier_0_2_10, s_Multiplier_0_2_11, f_s_Multiplier_0_2_11, 
        s_Multiplier_0_2_12, f_s_Multiplier_0_2_12, s_Multiplier_0_2_13, 
        f_s_Multiplier_0_2_13, s_Multiplier_0_2_14, f_s_Multiplier_0_2_14, 
        s_Multiplier_0_2_15, f_s_Multiplier_0_2_15, s_Multiplier_0_2_16, 
        f_s_Multiplier_0_2_16, s_Multiplier_0_2_17, f_s_Multiplier_0_2_17, 
        s_Multiplier_0_2_18, f_s_Multiplier_0_2_18, s_Multiplier_0_2_19, 
        f_s_Multiplier_0_2_19, s_Multiplier_0_2_20, f_s_Multiplier_0_2_20, 
        s_Multiplier_0_2_21, f_s_Multiplier_0_2_21, s_Multiplier_0_2_22, 
        f_s_Multiplier_0_2_22, s_Multiplier_0_2_23, f_s_Multiplier_0_2_23, 
        Multiplier_0_cin_lr_0, Multiplier_0_pp_0_13, mfco, Multiplier_0_cin_lr_2, 
        Multiplier_0_pp_1_15, mfco_1, Multiplier_0_cin_lr_4, Multiplier_0_pp_2_17, 
        mfco_2, Multiplier_0_cin_lr_6, Multiplier_0_pp_3_19, mfco_3, 
        Multiplier_0_cin_lr_8, Multiplier_0_pp_4_21, mfco_4, Multiplier_0_cin_lr_10, 
        Multiplier_0_pp_5_23, mfco_5, co_Multiplier_0_0_1, Multiplier_0_pp_0_2, 
        co_Multiplier_0_0_2, Multiplier_0_pp_0_4, Multiplier_0_pp_0_3, 
        Multiplier_0_pp_1_4, Multiplier_0_pp_1_3, co_Multiplier_0_0_3, 
        Multiplier_0_pp_0_6, Multiplier_0_pp_0_5, Multiplier_0_pp_1_6, 
        Multiplier_0_pp_1_5, co_Multiplier_0_0_4, Multiplier_0_pp_0_8, 
        Multiplier_0_pp_0_7, Multiplier_0_pp_1_8, Multiplier_0_pp_1_7, 
        co_Multiplier_0_0_5, Multiplier_0_pp_0_10, Multiplier_0_pp_0_9, 
        Multiplier_0_pp_1_10, Multiplier_0_pp_1_9, co_Multiplier_0_0_6, 
        Multiplier_0_pp_0_12, Multiplier_0_pp_0_11, Multiplier_0_pp_1_12, 
        Multiplier_0_pp_1_11, co_Multiplier_0_0_7, Multiplier_0_pp_1_14, 
        Multiplier_0_pp_1_13, co_Multiplier_0_0_8, co_Multiplier_0_1_1, 
        Multiplier_0_pp_2_6, co_Multiplier_0_1_2, Multiplier_0_pp_2_8, 
        Multiplier_0_pp_2_7, Multiplier_0_pp_3_8, Multiplier_0_pp_3_7, 
        co_Multiplier_0_1_3, Multiplier_0_pp_2_10, Multiplier_0_pp_2_9, 
        Multiplier_0_pp_3_10, Multiplier_0_pp_3_9, co_Multiplier_0_1_4, 
        Multiplier_0_pp_2_12, Multiplier_0_pp_2_11, Multiplier_0_pp_3_12, 
        Multiplier_0_pp_3_11, co_Multiplier_0_1_5, Multiplier_0_pp_2_14, 
        Multiplier_0_pp_2_13, Multiplier_0_pp_3_14, Multiplier_0_pp_3_13, 
        co_Multiplier_0_1_6, Multiplier_0_pp_2_16, Multiplier_0_pp_2_15, 
        Multiplier_0_pp_3_16, Multiplier_0_pp_3_15, co_Multiplier_0_1_7, 
        Multiplier_0_pp_3_18, Multiplier_0_pp_3_17, co_Multiplier_0_1_8, 
        co_Multiplier_0_2_1, Multiplier_0_pp_4_10, co_Multiplier_0_2_2, 
        Multiplier_0_pp_4_12, Multiplier_0_pp_4_11, Multiplier_0_pp_5_12, 
        Multiplier_0_pp_5_11, co_Multiplier_0_2_3, Multiplier_0_pp_4_14, 
        Multiplier_0_pp_4_13, Multiplier_0_pp_5_14, Multiplier_0_pp_5_13, 
        co_Multiplier_0_2_4, Multiplier_0_pp_4_16, Multiplier_0_pp_4_15, 
        Multiplier_0_pp_5_16, Multiplier_0_pp_5_15, co_Multiplier_0_2_5, 
        Multiplier_0_pp_4_18, Multiplier_0_pp_4_17, Multiplier_0_pp_5_18, 
        Multiplier_0_pp_5_17, co_Multiplier_0_2_6, Multiplier_0_pp_4_20, 
        Multiplier_0_pp_4_19, Multiplier_0_pp_5_20, Multiplier_0_pp_5_19, 
        co_Multiplier_0_2_7, Multiplier_0_pp_5_22, Multiplier_0_pp_5_21, 
        co_Multiplier_0_3_1, co_Multiplier_0_3_2, co_Multiplier_0_3_3, 
        s_Multiplier_0_3_8, co_Multiplier_0_3_4, s_Multiplier_0_3_9, s_Multiplier_0_3_10, 
        co_Multiplier_0_3_5, s_Multiplier_0_3_11, s_Multiplier_0_3_12, 
        co_Multiplier_0_3_6, s_Multiplier_0_3_13, s_Multiplier_0_3_14, 
        co_Multiplier_0_3_7, s_Multiplier_0_3_15, s_Multiplier_0_3_16, 
        co_Multiplier_0_3_8, s_Multiplier_0_3_17, s_Multiplier_0_3_18, 
        co_Multiplier_0_3_9, s_Multiplier_0_3_19, s_Multiplier_0_3_20, 
        co_Multiplier_0_3_10, s_Multiplier_0_3_21, s_Multiplier_0_3_22, 
        s_Multiplier_0_3_23, co_t_Multiplier_0_4_1, co_t_Multiplier_0_4_2, 
        co_t_Multiplier_0_4_3, co_t_Multiplier_0_4_4, co_t_Multiplier_0_4_5, 
        co_t_Multiplier_0_4_6, co_t_Multiplier_0_4_7, co_t_Multiplier_0_4_8, 
        mco, mco_1, mco_2, mco_3, mco_4, Multiplier_0_mult_0_5_n2, 
        mco_5, mco_6, mco_7, mco_8, mco_9, Multiplier_0_mult_2_5_n2, 
        mco_10, mco_11, mco_12, mco_13, mco_14, Multiplier_0_mult_4_5_n2, 
        mco_15, mco_16, mco_17, mco_18, mco_19, Multiplier_0_mult_6_5_n2, 
        mco_20, mco_21, mco_22, mco_23, mco_24, Multiplier_0_mult_8_5_n2, 
        Multiplier_0_mult_10_0_n1, mco_25, mco_26, mco_27, mco_28, 
        mco_29;
    
    ND2 ND2_t25 (.A(rega_a_11), .B(regb_b_1), .Z(Multiplier_0_mult_0_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    AND2 AND2_t24 (.A(regb_b_0), .B(regb_b_2), .Z(Multiplier_0_pp_1_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(382[10:72])
    ND2 ND2_t22 (.A(rega_a_11), .B(regb_b_3), .Z(Multiplier_0_mult_2_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    AND2 AND2_t21 (.A(regb_b_0), .B(regb_b_4), .Z(Multiplier_0_pp_2_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(388[10:72])
    ND2 ND2_t19 (.A(rega_a_11), .B(regb_b_5), .Z(Multiplier_0_mult_4_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    AND2 AND2_t18 (.A(regb_b_0), .B(regb_b_6), .Z(Multiplier_0_pp_3_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(394[10:72])
    ND2 ND2_t16 (.A(rega_a_11), .B(regb_b_7), .Z(Multiplier_0_mult_6_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    AND2 AND2_t15 (.A(regb_b_0), .B(regb_b_8), .Z(Multiplier_0_pp_4_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(400[10:72])
    ND2 ND2_t13 (.A(rega_a_11), .B(regb_b_9), .Z(Multiplier_0_mult_8_5_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    AND2 AND2_t12 (.A(regb_b_0), .B(regb_b_10), .Z(Multiplier_0_pp_5_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(406[10:74])
    ND2 ND2_t10 (.A(regb_b_0), .B(regb_b_11), .Z(Multiplier_0_mult_10_0_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t9 (.A(rega_a_3), .B(regb_b_11), .Z(Multiplier_0_mult_10_1_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t8 (.A(rega_a_2), .B(regb_b_11), .Z(Multiplier_0_mult_10_1_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t7 (.A(rega_a_5), .B(regb_b_11), .Z(Multiplier_0_mult_10_2_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t6 (.A(rega_a_4), .B(regb_b_11), .Z(Multiplier_0_mult_10_2_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t5 (.A(rega_a_7), .B(regb_b_11), .Z(Multiplier_0_mult_10_3_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t4 (.A(rega_a_6), .B(regb_b_11), .Z(Multiplier_0_mult_10_3_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t3 (.A(rega_a_9), .B(regb_b_11), .Z(Multiplier_0_mult_10_4_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t2 (.A(rega_a_8), .B(regb_b_11), .Z(Multiplier_0_mult_10_4_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t1 (.A(rega_a_11), .B(regb_b_10), .Z(Multiplier_0_mult_10_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t0 (.A(rega_a_10), .B(regb_b_11), .Z(Multiplier_0_mult_10_5_n0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FD1P3DX FF_98 (.D(MultDataB[1]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(435[13:82])
    defparam FF_98.GSR = "ENABLED";
    FD1P3DX FF_97 (.D(MultDataB[2]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(438[13:82])
    defparam FF_97.GSR = "ENABLED";
    FD1P3DX FF_96 (.D(MultDataB[3]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(441[13:82])
    defparam FF_96.GSR = "ENABLED";
    FD1P3DX FF_95 (.D(MultDataB[4]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(444[13:82])
    defparam FF_95.GSR = "ENABLED";
    FD1P3DX FF_94 (.D(MultDataB[5]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(447[13:82])
    defparam FF_94.GSR = "ENABLED";
    FD1P3DX FF_93 (.D(MultDataB[6]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(450[13:82])
    defparam FF_93.GSR = "ENABLED";
    FD1P3DX FF_92 (.D(MultDataB[7]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(453[13:82])
    defparam FF_92.GSR = "ENABLED";
    FD1P3DX FF_91 (.D(MultDataB[8]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(456[13:82])
    defparam FF_91.GSR = "ENABLED";
    FD1P3DX FF_90 (.D(MultDataB[9]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(459[13:82])
    defparam FF_90.GSR = "ENABLED";
    FD1P3DX FF_89 (.D(MultDataB[10]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(462[13:84])
    defparam FF_89.GSR = "ENABLED";
    FD1P3DX FF_88 (.D(MultDataB[11]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rega_a_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(465[13:84])
    defparam FF_88.GSR = "ENABLED";
    FD1P3DX FF_87 (.D(MultDataB[0]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_0)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(468[13:82])
    defparam FF_87.GSR = "ENABLED";
    FD1P3DX FF_86 (.D(MultDataB[1]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(471[13:82])
    defparam FF_86.GSR = "ENABLED";
    FD1P3DX FF_85 (.D(MultDataB[2]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(474[13:82])
    defparam FF_85.GSR = "ENABLED";
    FD1P3DX FF_84 (.D(MultDataB[3]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(477[13:82])
    defparam FF_84.GSR = "ENABLED";
    FD1P3DX FF_83 (.D(MultDataB[4]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(480[13:82])
    defparam FF_83.GSR = "ENABLED";
    FD1P3DX FF_82 (.D(MultDataB[5]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(483[13:82])
    defparam FF_82.GSR = "ENABLED";
    FD1P3DX FF_81 (.D(MultDataB[6]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(486[13:82])
    defparam FF_81.GSR = "ENABLED";
    FD1P3DX FF_80 (.D(MultDataB[7]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(489[13:82])
    defparam FF_80.GSR = "ENABLED";
    FD1P3DX FF_79 (.D(MultDataB[8]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(492[13:82])
    defparam FF_79.GSR = "ENABLED";
    FD1P3DX FF_78 (.D(MultDataB[9]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(495[13:82])
    defparam FF_78.GSR = "ENABLED";
    FD1P3DX FF_77 (.D(MultDataB[10]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(498[13:84])
    defparam FF_77.GSR = "ENABLED";
    FD1P3DX FF_76 (.D(MultDataB[11]), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(regb_b_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(501[13:84])
    defparam FF_76.GSR = "ENABLED";
    FD1P3DX FF_75 (.D(rego_o_0), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[0])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(504[13:83])
    defparam FF_75.GSR = "ENABLED";
    FD1P3DX FF_74 (.D(rego_o_1), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[1])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(507[13:83])
    defparam FF_74.GSR = "ENABLED";
    FD1P3DX FF_73 (.D(rego_o_2), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[2])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(510[13:83])
    defparam FF_73.GSR = "ENABLED";
    FD1P3DX FF_72 (.D(rego_o_3), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[3])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(513[13:83])
    defparam FF_72.GSR = "ENABLED";
    FD1P3DX FF_71 (.D(rego_o_4), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[4])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(516[13:83])
    defparam FF_71.GSR = "ENABLED";
    FD1P3DX FF_70 (.D(rego_o_5), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[5])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(519[13:83])
    defparam FF_70.GSR = "ENABLED";
    FD1P3DX FF_69 (.D(rego_o_6), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[6])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(522[13:83])
    defparam FF_69.GSR = "ENABLED";
    FD1P3DX FF_68 (.D(rego_o_7), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[7])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(525[13:83])
    defparam FF_68.GSR = "ENABLED";
    FD1P3DX FF_67 (.D(rego_o_8), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[8])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(528[13:83])
    defparam FF_67.GSR = "ENABLED";
    FD1P3DX FF_66 (.D(rego_o_9), .SP(VCC_net), .CK(CIC1_out_clkSin), .CD(GND_net), 
            .Q(MultResult1[9])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(531[13:83])
    defparam FF_66.GSR = "ENABLED";
    FD1P3DX FF_65 (.D(rego_o_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[10])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(534[13:85])
    defparam FF_65.GSR = "ENABLED";
    FD1P3DX FF_64 (.D(rego_o_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[11])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(537[13:85])
    defparam FF_64.GSR = "ENABLED";
    FD1P3DX FF_63 (.D(rego_o_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[12])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(540[13:85])
    defparam FF_63.GSR = "ENABLED";
    FD1P3DX FF_62 (.D(rego_o_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[13])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(543[13:85])
    defparam FF_62.GSR = "ENABLED";
    FD1P3DX FF_61 (.D(rego_o_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[14])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(546[13:85])
    defparam FF_61.GSR = "ENABLED";
    FD1P3DX FF_60 (.D(rego_o_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[15])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(549[13:85])
    defparam FF_60.GSR = "ENABLED";
    FD1P3DX FF_59 (.D(rego_o_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[16])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(552[13:85])
    defparam FF_59.GSR = "ENABLED";
    FD1P3DX FF_58 (.D(rego_o_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[17])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(555[13:85])
    defparam FF_58.GSR = "ENABLED";
    FD1P3DX FF_57 (.D(rego_o_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[18])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(558[13:85])
    defparam FF_57.GSR = "ENABLED";
    FD1P3DX FF_56 (.D(rego_o_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[19])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(561[13:85])
    defparam FF_56.GSR = "ENABLED";
    FD1P3DX FF_55 (.D(rego_o_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[20])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(564[13:85])
    defparam FF_55.GSR = "ENABLED";
    FD1P3DX FF_54 (.D(rego_o_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[21])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(567[13:85])
    defparam FF_54.GSR = "ENABLED";
    FD1P3DX FF_53 (.D(rego_o_22), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[22])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(570[13:85])
    defparam FF_53.GSR = "ENABLED";
    FD1P3DX FF_52 (.D(rego_o_23), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(MultResult1[23])) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(573[13:85])
    defparam FF_52.GSR = "ENABLED";
    FD1P3DX FF_51 (.D(Multiplier_0_pp_0_0), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_0)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(576[13] 577[35])
    defparam FF_51.GSR = "ENABLED";
    FD1P3DX FF_50 (.D(Multiplier_0_pp_0_1), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(580[13] 581[35])
    defparam FF_50.GSR = "ENABLED";
    FD1P3DX FF_49 (.D(s_Multiplier_0_0_2), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(584[13] 585[34])
    defparam FF_49.GSR = "ENABLED";
    FD1P3DX FF_48 (.D(s_Multiplier_0_0_3), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(rego_o_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(588[13] 589[34])
    defparam FF_48.GSR = "ENABLED";
    FD1P3DX FF_47 (.D(s_Multiplier_0_0_4), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(592[13] 593[34])
    defparam FF_47.GSR = "ENABLED";
    FD1P3DX FF_46 (.D(s_Multiplier_0_0_5), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(596[13] 597[34])
    defparam FF_46.GSR = "ENABLED";
    FD1P3DX FF_45 (.D(s_Multiplier_0_0_6), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(600[13] 601[34])
    defparam FF_45.GSR = "ENABLED";
    FD1P3DX FF_44 (.D(s_Multiplier_0_0_7), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(604[13] 605[34])
    defparam FF_44.GSR = "ENABLED";
    FD1P3DX FF_43 (.D(s_Multiplier_0_0_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(608[13] 609[34])
    defparam FF_43.GSR = "ENABLED";
    FD1P3DX FF_42 (.D(s_Multiplier_0_0_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(612[13] 613[34])
    defparam FF_42.GSR = "ENABLED";
    FD1P3DX FF_41 (.D(s_Multiplier_0_0_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(616[13] 617[35])
    defparam FF_41.GSR = "ENABLED";
    FD1P3DX FF_40 (.D(s_Multiplier_0_0_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(620[13] 621[35])
    defparam FF_40.GSR = "ENABLED";
    FD1P3DX FF_39 (.D(s_Multiplier_0_0_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(624[13] 625[35])
    defparam FF_39.GSR = "ENABLED";
    FD1P3DX FF_38 (.D(s_Multiplier_0_0_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(628[13] 629[35])
    defparam FF_38.GSR = "ENABLED";
    FD1P3DX FF_37 (.D(s_Multiplier_0_0_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(632[13] 633[35])
    defparam FF_37.GSR = "ENABLED";
    FD1P3DX FF_36 (.D(s_Multiplier_0_0_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(636[13] 637[35])
    defparam FF_36.GSR = "ENABLED";
    FD1P3DX FF_35 (.D(s_Multiplier_0_0_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(640[13] 641[35])
    defparam FF_35.GSR = "ENABLED";
    FD1P3DX FF_34 (.D(s_Multiplier_0_0_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_0_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(644[13] 645[35])
    defparam FF_34.GSR = "ENABLED";
    FD1P3DX FF_33 (.D(Multiplier_0_pp_2_4), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_2_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(648[13] 649[35])
    defparam FF_33.GSR = "ENABLED";
    FD1P3DX FF_32 (.D(Multiplier_0_pp_2_5), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_2_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(652[13] 653[35])
    defparam FF_32.GSR = "ENABLED";
    FD1P3DX FF_31 (.D(s_Multiplier_0_1_6), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(656[13] 657[34])
    defparam FF_31.GSR = "ENABLED";
    FD1P3DX FF_30 (.D(s_Multiplier_0_1_7), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(660[13] 661[34])
    defparam FF_30.GSR = "ENABLED";
    FD1P3DX FF_29 (.D(s_Multiplier_0_1_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(664[13] 665[34])
    defparam FF_29.GSR = "ENABLED";
    FD1P3DX FF_28 (.D(s_Multiplier_0_1_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(668[13] 669[34])
    defparam FF_28.GSR = "ENABLED";
    FD1P3DX FF_27 (.D(s_Multiplier_0_1_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(672[13] 673[35])
    defparam FF_27.GSR = "ENABLED";
    FD1P3DX FF_26 (.D(s_Multiplier_0_1_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(676[13] 677[35])
    defparam FF_26.GSR = "ENABLED";
    FD1P3DX FF_25 (.D(s_Multiplier_0_1_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(680[13] 681[35])
    defparam FF_25.GSR = "ENABLED";
    FD1P3DX FF_24 (.D(s_Multiplier_0_1_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(684[13] 685[35])
    defparam FF_24.GSR = "ENABLED";
    FD1P3DX FF_23 (.D(s_Multiplier_0_1_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(688[13] 689[35])
    defparam FF_23.GSR = "ENABLED";
    FD1P3DX FF_22 (.D(s_Multiplier_0_1_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(692[13] 693[35])
    defparam FF_22.GSR = "ENABLED";
    FD1P3DX FF_21 (.D(s_Multiplier_0_1_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(696[13] 697[35])
    defparam FF_21.GSR = "ENABLED";
    FD1P3DX FF_20 (.D(s_Multiplier_0_1_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(700[13] 701[35])
    defparam FF_20.GSR = "ENABLED";
    FD1P3DX FF_19 (.D(s_Multiplier_0_1_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(704[13] 705[35])
    defparam FF_19.GSR = "ENABLED";
    FD1P3DX FF_18 (.D(s_Multiplier_0_1_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(708[13] 709[35])
    defparam FF_18.GSR = "ENABLED";
    FD1P3DX FF_17 (.D(s_Multiplier_0_1_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(712[13] 713[35])
    defparam FF_17.GSR = "ENABLED";
    FD1P3DX FF_16 (.D(s_Multiplier_0_1_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_1_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(716[13] 717[35])
    defparam FF_16.GSR = "ENABLED";
    FD1P3DX FF_15 (.D(Multiplier_0_pp_4_8), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_4_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(720[13] 721[35])
    defparam FF_15.GSR = "ENABLED";
    FD1P3DX FF_14 (.D(Multiplier_0_pp_4_9), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_Multiplier_0_pp_4_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(724[13] 725[35])
    defparam FF_14.GSR = "ENABLED";
    FD1P3DX FF_13 (.D(s_Multiplier_0_2_10), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(728[13] 729[35])
    defparam FF_13.GSR = "ENABLED";
    FD1P3DX FF_12 (.D(s_Multiplier_0_2_11), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(732[13] 733[35])
    defparam FF_12.GSR = "ENABLED";
    FD1P3DX FF_11 (.D(s_Multiplier_0_2_12), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(736[13] 737[35])
    defparam FF_11.GSR = "ENABLED";
    FD1P3DX FF_10 (.D(s_Multiplier_0_2_13), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(740[13] 741[35])
    defparam FF_10.GSR = "ENABLED";
    FD1P3DX FF_9 (.D(s_Multiplier_0_2_14), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(744[13] 745[35])
    defparam FF_9.GSR = "ENABLED";
    FD1P3DX FF_8 (.D(s_Multiplier_0_2_15), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(748[13] 749[35])
    defparam FF_8.GSR = "ENABLED";
    FD1P3DX FF_7 (.D(s_Multiplier_0_2_16), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(752[13] 753[35])
    defparam FF_7.GSR = "ENABLED";
    FD1P3DX FF_6 (.D(s_Multiplier_0_2_17), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(756[13] 757[35])
    defparam FF_6.GSR = "ENABLED";
    FD1P3DX FF_5 (.D(s_Multiplier_0_2_18), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(760[13] 761[35])
    defparam FF_5.GSR = "ENABLED";
    FD1P3DX FF_4 (.D(s_Multiplier_0_2_19), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(764[13] 765[35])
    defparam FF_4.GSR = "ENABLED";
    FD1P3DX FF_3 (.D(s_Multiplier_0_2_20), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(768[13] 769[35])
    defparam FF_3.GSR = "ENABLED";
    FD1P3DX FF_2 (.D(s_Multiplier_0_2_21), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(772[13] 773[35])
    defparam FF_2.GSR = "ENABLED";
    FD1P3DX FF_1 (.D(s_Multiplier_0_2_22), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_22)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(776[13] 777[35])
    defparam FF_1.GSR = "ENABLED";
    FD1P3DX FF_0 (.D(s_Multiplier_0_2_23), .SP(VCC_net), .CK(CIC1_out_clkSin), 
            .CD(GND_net), .Q(f_s_Multiplier_0_2_23)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(780[13] 781[35])
    defparam FF_0.GSR = "ENABLED";
    FADD2B Multiplier_0_cin_lr_add_0 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_Cadd_0_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco), .S0(Multiplier_0_pp_0_13)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_cin_lr_add_2 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_Cadd_2_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_1), .S0(Multiplier_0_pp_1_15)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_cin_lr_add_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_Cadd_4_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_2), .S0(Multiplier_0_pp_2_17)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_cin_lr_add_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_Cadd_6_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_3), .S0(Multiplier_0_pp_3_19)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_cin_lr_add_8 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_Cadd_8_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_4), .S0(Multiplier_0_pp_4_21)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_cin_lr_add_10 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(Multiplier_0_cin_lr_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_Cadd_10_6 (.A0(VCC_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_5), .S0(Multiplier_0_pp_5_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_Multiplier_0_0_1 (.A0(GND_net), .A1(Multiplier_0_pp_0_2), 
           .B0(GND_net), .B1(Multiplier_0_pp_1_2), .CI(GND_net), .COUT(co_Multiplier_0_0_1), 
           .S1(s_Multiplier_0_0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_0_2 (.A0(Multiplier_0_pp_0_3), .A1(Multiplier_0_pp_0_4), 
           .B0(Multiplier_0_pp_1_3), .B1(Multiplier_0_pp_1_4), .CI(co_Multiplier_0_0_1), 
           .COUT(co_Multiplier_0_0_2), .S0(s_Multiplier_0_0_3), .S1(s_Multiplier_0_0_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_0_3 (.A0(Multiplier_0_pp_0_5), .A1(Multiplier_0_pp_0_6), 
           .B0(Multiplier_0_pp_1_5), .B1(Multiplier_0_pp_1_6), .CI(co_Multiplier_0_0_2), 
           .COUT(co_Multiplier_0_0_3), .S0(s_Multiplier_0_0_5), .S1(s_Multiplier_0_0_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_0_4 (.A0(Multiplier_0_pp_0_7), .A1(Multiplier_0_pp_0_8), 
           .B0(Multiplier_0_pp_1_7), .B1(Multiplier_0_pp_1_8), .CI(co_Multiplier_0_0_3), 
           .COUT(co_Multiplier_0_0_4), .S0(s_Multiplier_0_0_7), .S1(s_Multiplier_0_0_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_0_5 (.A0(Multiplier_0_pp_0_9), .A1(Multiplier_0_pp_0_10), 
           .B0(Multiplier_0_pp_1_9), .B1(Multiplier_0_pp_1_10), .CI(co_Multiplier_0_0_4), 
           .COUT(co_Multiplier_0_0_5), .S0(s_Multiplier_0_0_9), .S1(s_Multiplier_0_0_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_0_6 (.A0(Multiplier_0_pp_0_11), .A1(Multiplier_0_pp_0_12), 
           .B0(Multiplier_0_pp_1_11), .B1(Multiplier_0_pp_1_12), .CI(co_Multiplier_0_0_5), 
           .COUT(co_Multiplier_0_0_6), .S0(s_Multiplier_0_0_11), .S1(s_Multiplier_0_0_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_0_7 (.A0(Multiplier_0_pp_0_13), .A1(GND_net), 
           .B0(Multiplier_0_pp_1_13), .B1(Multiplier_0_pp_1_14), .CI(co_Multiplier_0_0_6), 
           .COUT(co_Multiplier_0_0_7), .S0(s_Multiplier_0_0_13), .S1(s_Multiplier_0_0_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_0_8 (.A0(GND_net), .A1(GND_net), .B0(Multiplier_0_pp_1_15), 
           .B1(GND_net), .CI(co_Multiplier_0_0_7), .COUT(co_Multiplier_0_0_8), 
           .S0(s_Multiplier_0_0_15), .S1(s_Multiplier_0_0_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_Multiplier_0_0_9 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_Multiplier_0_0_8), .S0(s_Multiplier_0_0_17)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_Multiplier_0_1_1 (.A0(GND_net), .A1(Multiplier_0_pp_2_6), 
           .B0(GND_net), .B1(Multiplier_0_pp_3_6), .CI(GND_net), .COUT(co_Multiplier_0_1_1), 
           .S1(s_Multiplier_0_1_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_1_2 (.A0(Multiplier_0_pp_2_7), .A1(Multiplier_0_pp_2_8), 
           .B0(Multiplier_0_pp_3_7), .B1(Multiplier_0_pp_3_8), .CI(co_Multiplier_0_1_1), 
           .COUT(co_Multiplier_0_1_2), .S0(s_Multiplier_0_1_7), .S1(s_Multiplier_0_1_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_1_3 (.A0(Multiplier_0_pp_2_9), .A1(Multiplier_0_pp_2_10), 
           .B0(Multiplier_0_pp_3_9), .B1(Multiplier_0_pp_3_10), .CI(co_Multiplier_0_1_2), 
           .COUT(co_Multiplier_0_1_3), .S0(s_Multiplier_0_1_9), .S1(s_Multiplier_0_1_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_1_4 (.A0(Multiplier_0_pp_2_11), .A1(Multiplier_0_pp_2_12), 
           .B0(Multiplier_0_pp_3_11), .B1(Multiplier_0_pp_3_12), .CI(co_Multiplier_0_1_3), 
           .COUT(co_Multiplier_0_1_4), .S0(s_Multiplier_0_1_11), .S1(s_Multiplier_0_1_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_1_5 (.A0(Multiplier_0_pp_2_13), .A1(Multiplier_0_pp_2_14), 
           .B0(Multiplier_0_pp_3_13), .B1(Multiplier_0_pp_3_14), .CI(co_Multiplier_0_1_4), 
           .COUT(co_Multiplier_0_1_5), .S0(s_Multiplier_0_1_13), .S1(s_Multiplier_0_1_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_1_6 (.A0(Multiplier_0_pp_2_15), .A1(Multiplier_0_pp_2_16), 
           .B0(Multiplier_0_pp_3_15), .B1(Multiplier_0_pp_3_16), .CI(co_Multiplier_0_1_5), 
           .COUT(co_Multiplier_0_1_6), .S0(s_Multiplier_0_1_15), .S1(s_Multiplier_0_1_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_1_7 (.A0(Multiplier_0_pp_2_17), .A1(GND_net), 
           .B0(Multiplier_0_pp_3_17), .B1(Multiplier_0_pp_3_18), .CI(co_Multiplier_0_1_6), 
           .COUT(co_Multiplier_0_1_7), .S0(s_Multiplier_0_1_17), .S1(s_Multiplier_0_1_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_1_8 (.A0(GND_net), .A1(GND_net), .B0(Multiplier_0_pp_3_19), 
           .B1(GND_net), .CI(co_Multiplier_0_1_7), .COUT(co_Multiplier_0_1_8), 
           .S0(s_Multiplier_0_1_19), .S1(s_Multiplier_0_1_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_Multiplier_0_1_9 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_Multiplier_0_1_8), .S0(s_Multiplier_0_1_21)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_Multiplier_0_2_1 (.A0(GND_net), .A1(Multiplier_0_pp_4_10), 
           .B0(GND_net), .B1(Multiplier_0_pp_5_10), .CI(GND_net), .COUT(co_Multiplier_0_2_1), 
           .S1(s_Multiplier_0_2_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_2_2 (.A0(Multiplier_0_pp_4_11), .A1(Multiplier_0_pp_4_12), 
           .B0(Multiplier_0_pp_5_11), .B1(Multiplier_0_pp_5_12), .CI(co_Multiplier_0_2_1), 
           .COUT(co_Multiplier_0_2_2), .S0(s_Multiplier_0_2_11), .S1(s_Multiplier_0_2_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_2_3 (.A0(Multiplier_0_pp_4_13), .A1(Multiplier_0_pp_4_14), 
           .B0(Multiplier_0_pp_5_13), .B1(Multiplier_0_pp_5_14), .CI(co_Multiplier_0_2_2), 
           .COUT(co_Multiplier_0_2_3), .S0(s_Multiplier_0_2_13), .S1(s_Multiplier_0_2_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_2_4 (.A0(Multiplier_0_pp_4_15), .A1(Multiplier_0_pp_4_16), 
           .B0(Multiplier_0_pp_5_15), .B1(Multiplier_0_pp_5_16), .CI(co_Multiplier_0_2_3), 
           .COUT(co_Multiplier_0_2_4), .S0(s_Multiplier_0_2_15), .S1(s_Multiplier_0_2_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_2_5 (.A0(Multiplier_0_pp_4_17), .A1(Multiplier_0_pp_4_18), 
           .B0(Multiplier_0_pp_5_17), .B1(Multiplier_0_pp_5_18), .CI(co_Multiplier_0_2_4), 
           .COUT(co_Multiplier_0_2_5), .S0(s_Multiplier_0_2_17), .S1(s_Multiplier_0_2_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_2_6 (.A0(Multiplier_0_pp_4_19), .A1(Multiplier_0_pp_4_20), 
           .B0(Multiplier_0_pp_5_19), .B1(Multiplier_0_pp_5_20), .CI(co_Multiplier_0_2_5), 
           .COUT(co_Multiplier_0_2_6), .S0(s_Multiplier_0_2_19), .S1(s_Multiplier_0_2_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_2_7 (.A0(Multiplier_0_pp_4_21), .A1(GND_net), 
           .B0(Multiplier_0_pp_5_21), .B1(Multiplier_0_pp_5_22), .CI(co_Multiplier_0_2_6), 
           .COUT(co_Multiplier_0_2_7), .S0(s_Multiplier_0_2_21), .S1(s_Multiplier_0_2_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_2_8 (.A0(GND_net), .A1(GND_net), .B0(Multiplier_0_pp_5_23), 
           .B1(GND_net), .CI(co_Multiplier_0_2_7), .S0(s_Multiplier_0_2_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_Multiplier_0_3_1 (.A0(GND_net), .A1(f_s_Multiplier_0_0_4), 
           .B0(GND_net), .B1(f_Multiplier_0_pp_2_4), .CI(GND_net), .COUT(co_Multiplier_0_3_1), 
           .S1(rego_o_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_2 (.A0(f_s_Multiplier_0_0_5), .A1(f_s_Multiplier_0_0_6), 
           .B0(f_Multiplier_0_pp_2_5), .B1(f_s_Multiplier_0_1_6), .CI(co_Multiplier_0_3_1), 
           .COUT(co_Multiplier_0_3_2), .S0(rego_o_5), .S1(rego_o_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_3 (.A0(f_s_Multiplier_0_0_7), .A1(f_s_Multiplier_0_0_8), 
           .B0(f_s_Multiplier_0_1_7), .B1(f_s_Multiplier_0_1_8), .CI(co_Multiplier_0_3_2), 
           .COUT(co_Multiplier_0_3_3), .S0(rego_o_7), .S1(s_Multiplier_0_3_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_4 (.A0(f_s_Multiplier_0_0_9), .A1(f_s_Multiplier_0_0_10), 
           .B0(f_s_Multiplier_0_1_9), .B1(f_s_Multiplier_0_1_10), .CI(co_Multiplier_0_3_3), 
           .COUT(co_Multiplier_0_3_4), .S0(s_Multiplier_0_3_9), .S1(s_Multiplier_0_3_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_5 (.A0(f_s_Multiplier_0_0_11), .A1(f_s_Multiplier_0_0_12), 
           .B0(f_s_Multiplier_0_1_11), .B1(f_s_Multiplier_0_1_12), .CI(co_Multiplier_0_3_4), 
           .COUT(co_Multiplier_0_3_5), .S0(s_Multiplier_0_3_11), .S1(s_Multiplier_0_3_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_6 (.A0(f_s_Multiplier_0_0_13), .A1(f_s_Multiplier_0_0_14), 
           .B0(f_s_Multiplier_0_1_13), .B1(f_s_Multiplier_0_1_14), .CI(co_Multiplier_0_3_5), 
           .COUT(co_Multiplier_0_3_6), .S0(s_Multiplier_0_3_13), .S1(s_Multiplier_0_3_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_7 (.A0(f_s_Multiplier_0_0_15), .A1(f_s_Multiplier_0_0_16), 
           .B0(f_s_Multiplier_0_1_15), .B1(f_s_Multiplier_0_1_16), .CI(co_Multiplier_0_3_6), 
           .COUT(co_Multiplier_0_3_7), .S0(s_Multiplier_0_3_15), .S1(s_Multiplier_0_3_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_8 (.A0(f_s_Multiplier_0_0_17), .A1(GND_net), 
           .B0(f_s_Multiplier_0_1_17), .B1(f_s_Multiplier_0_1_18), .CI(co_Multiplier_0_3_7), 
           .COUT(co_Multiplier_0_3_8), .S0(s_Multiplier_0_3_17), .S1(s_Multiplier_0_3_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_9 (.A0(GND_net), .A1(GND_net), .B0(f_s_Multiplier_0_1_19), 
           .B1(f_s_Multiplier_0_1_20), .CI(co_Multiplier_0_3_8), .COUT(co_Multiplier_0_3_9), 
           .S0(s_Multiplier_0_3_19), .S1(s_Multiplier_0_3_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Multiplier_0_add_3_10 (.A0(GND_net), .A1(GND_net), .B0(f_s_Multiplier_0_1_21), 
           .B1(GND_net), .CI(co_Multiplier_0_3_9), .COUT(co_Multiplier_0_3_10), 
           .S0(s_Multiplier_0_3_21), .S1(s_Multiplier_0_3_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_Multiplier_0_3_11 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_Multiplier_0_3_10), .S0(s_Multiplier_0_3_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B Cadd_t_Multiplier_0_4_1 (.A0(GND_net), .A1(s_Multiplier_0_3_8), 
           .B0(GND_net), .B1(f_Multiplier_0_pp_4_8), .CI(GND_net), .COUT(co_t_Multiplier_0_4_1), 
           .S1(rego_o_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_2 (.A0(s_Multiplier_0_3_9), .A1(s_Multiplier_0_3_10), 
           .B0(f_Multiplier_0_pp_4_9), .B1(f_s_Multiplier_0_2_10), .CI(co_t_Multiplier_0_4_1), 
           .COUT(co_t_Multiplier_0_4_2), .S0(rego_o_9), .S1(rego_o_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_3 (.A0(s_Multiplier_0_3_11), .A1(s_Multiplier_0_3_12), 
           .B0(f_s_Multiplier_0_2_11), .B1(f_s_Multiplier_0_2_12), .CI(co_t_Multiplier_0_4_2), 
           .COUT(co_t_Multiplier_0_4_3), .S0(rego_o_11), .S1(rego_o_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_4 (.A0(s_Multiplier_0_3_13), .A1(s_Multiplier_0_3_14), 
           .B0(f_s_Multiplier_0_2_13), .B1(f_s_Multiplier_0_2_14), .CI(co_t_Multiplier_0_4_3), 
           .COUT(co_t_Multiplier_0_4_4), .S0(rego_o_13), .S1(rego_o_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_5 (.A0(s_Multiplier_0_3_15), .A1(s_Multiplier_0_3_16), 
           .B0(f_s_Multiplier_0_2_15), .B1(f_s_Multiplier_0_2_16), .CI(co_t_Multiplier_0_4_4), 
           .COUT(co_t_Multiplier_0_4_5), .S0(rego_o_15), .S1(rego_o_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_6 (.A0(s_Multiplier_0_3_17), .A1(s_Multiplier_0_3_18), 
           .B0(f_s_Multiplier_0_2_17), .B1(f_s_Multiplier_0_2_18), .CI(co_t_Multiplier_0_4_5), 
           .COUT(co_t_Multiplier_0_4_6), .S0(rego_o_17), .S1(rego_o_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_7 (.A0(s_Multiplier_0_3_19), .A1(s_Multiplier_0_3_20), 
           .B0(f_s_Multiplier_0_2_19), .B1(f_s_Multiplier_0_2_20), .CI(co_t_Multiplier_0_4_6), 
           .COUT(co_t_Multiplier_0_4_7), .S0(rego_o_19), .S1(rego_o_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_8 (.A0(s_Multiplier_0_3_21), .A1(s_Multiplier_0_3_22), 
           .B0(f_s_Multiplier_0_2_21), .B1(f_s_Multiplier_0_2_22), .CI(co_t_Multiplier_0_4_7), 
           .COUT(co_t_Multiplier_0_4_8), .S0(rego_o_21), .S1(rego_o_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    FADD2B t_Multiplier_0_add_4_9 (.A0(s_Multiplier_0_3_23), .A1(GND_net), 
           .B0(f_s_Multiplier_0_2_23), .B1(GND_net), .CI(co_t_Multiplier_0_4_8), 
           .S0(rego_o_23)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_0_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(Multiplier_0_cin_lr_0), .CO(mco), .P0(Multiplier_0_pp_0_1), 
          .P1(Multiplier_0_pp_0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_0_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco), .CO(mco_1), .P0(Multiplier_0_pp_0_3), 
          .P1(Multiplier_0_pp_0_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_0_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco_1), .CO(mco_2), .P0(Multiplier_0_pp_0_5), 
          .P1(Multiplier_0_pp_0_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_0_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco_2), .CO(mco_3), .P0(Multiplier_0_pp_0_7), 
          .P1(Multiplier_0_pp_0_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_0_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_1), .B1(regb_b_0), .B2(regb_b_1), 
          .B3(regb_b_0), .CI(mco_3), .CO(mco_4), .P0(Multiplier_0_pp_0_9), 
          .P1(Multiplier_0_pp_0_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_0_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_0_5_n2), 
          .A2(Multiplier_0_mult_0_5_n1), .A3(VCC_net), .B0(regb_b_1), 
          .B1(VCC_net), .B2(VCC_net), .B3(VCC_net), .CI(mco_4), .CO(mfco), 
          .P0(Multiplier_0_pp_0_11), .P1(Multiplier_0_pp_0_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_2_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(Multiplier_0_cin_lr_2), .CO(mco_5), .P0(Multiplier_0_pp_1_3), 
          .P1(Multiplier_0_pp_1_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_2_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_5), .CO(mco_6), .P0(Multiplier_0_pp_1_5), 
          .P1(Multiplier_0_pp_1_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_2_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_6), .CO(mco_7), .P0(Multiplier_0_pp_1_7), 
          .P1(Multiplier_0_pp_1_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_2_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_7), .CO(mco_8), .P0(Multiplier_0_pp_1_9), 
          .P1(Multiplier_0_pp_1_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_2_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_3), .B1(regb_b_2), .B2(regb_b_3), 
          .B3(regb_b_2), .CI(mco_8), .CO(mco_9), .P0(Multiplier_0_pp_1_11), 
          .P1(Multiplier_0_pp_1_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_2_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_2_5_n2), 
          .A2(Multiplier_0_mult_2_5_n1), .A3(GND_net), .B0(regb_b_3), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_2), .CI(mco_9), .CO(mfco_1), 
          .P0(Multiplier_0_pp_1_13), .P1(Multiplier_0_pp_1_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_4_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(Multiplier_0_cin_lr_4), .CO(mco_10), .P0(Multiplier_0_pp_2_5), 
          .P1(Multiplier_0_pp_2_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_4_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_10), .CO(mco_11), .P0(Multiplier_0_pp_2_7), 
          .P1(Multiplier_0_pp_2_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_4_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_11), .CO(mco_12), .P0(Multiplier_0_pp_2_9), 
          .P1(Multiplier_0_pp_2_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_4_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_12), .CO(mco_13), .P0(Multiplier_0_pp_2_11), 
          .P1(Multiplier_0_pp_2_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_4_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_5), .B1(regb_b_4), .B2(regb_b_5), 
          .B3(regb_b_4), .CI(mco_13), .CO(mco_14), .P0(Multiplier_0_pp_2_13), 
          .P1(Multiplier_0_pp_2_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_4_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_4_5_n2), 
          .A2(Multiplier_0_mult_4_5_n1), .A3(GND_net), .B0(regb_b_5), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_4), .CI(mco_14), .CO(mfco_2), 
          .P0(Multiplier_0_pp_2_15), .P1(Multiplier_0_pp_2_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_6_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(Multiplier_0_cin_lr_6), .CO(mco_15), .P0(Multiplier_0_pp_3_7), 
          .P1(Multiplier_0_pp_3_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_6_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_15), .CO(mco_16), .P0(Multiplier_0_pp_3_9), 
          .P1(Multiplier_0_pp_3_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_6_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_16), .CO(mco_17), .P0(Multiplier_0_pp_3_11), 
          .P1(Multiplier_0_pp_3_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_6_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_17), .CO(mco_18), .P0(Multiplier_0_pp_3_13), 
          .P1(Multiplier_0_pp_3_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_6_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_7), .B1(regb_b_6), .B2(regb_b_7), 
          .B3(regb_b_6), .CI(mco_18), .CO(mco_19), .P0(Multiplier_0_pp_3_15), 
          .P1(Multiplier_0_pp_3_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_6_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_6_5_n2), 
          .A2(Multiplier_0_mult_6_5_n1), .A3(GND_net), .B0(regb_b_7), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_6), .CI(mco_19), .CO(mfco_3), 
          .P0(Multiplier_0_pp_3_17), .P1(Multiplier_0_pp_3_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_8_0 (.A0(regb_b_0), .A1(rega_a_1), .A2(rega_a_1), 
          .A3(rega_a_2), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(Multiplier_0_cin_lr_8), .CO(mco_20), .P0(Multiplier_0_pp_4_9), 
          .P1(Multiplier_0_pp_4_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_8_1 (.A0(rega_a_2), .A1(rega_a_3), .A2(rega_a_3), 
          .A3(rega_a_4), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_20), .CO(mco_21), .P0(Multiplier_0_pp_4_11), 
          .P1(Multiplier_0_pp_4_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_8_2 (.A0(rega_a_4), .A1(rega_a_5), .A2(rega_a_5), 
          .A3(rega_a_6), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_21), .CO(mco_22), .P0(Multiplier_0_pp_4_13), 
          .P1(Multiplier_0_pp_4_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_8_3 (.A0(rega_a_6), .A1(rega_a_7), .A2(rega_a_7), 
          .A3(rega_a_8), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_22), .CO(mco_23), .P0(Multiplier_0_pp_4_15), 
          .P1(Multiplier_0_pp_4_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_8_4 (.A0(rega_a_8), .A1(rega_a_9), .A2(rega_a_9), 
          .A3(rega_a_10), .B0(regb_b_9), .B1(regb_b_8), .B2(regb_b_9), 
          .B3(regb_b_8), .CI(mco_23), .CO(mco_24), .P0(Multiplier_0_pp_4_17), 
          .P1(Multiplier_0_pp_4_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_8_5 (.A0(rega_a_10), .A1(Multiplier_0_mult_8_5_n2), 
          .A2(Multiplier_0_mult_8_5_n1), .A3(GND_net), .B0(regb_b_9), 
          .B1(VCC_net), .B2(VCC_net), .B3(regb_b_8), .CI(mco_24), .CO(mfco_4), 
          .P0(Multiplier_0_pp_4_19), .P1(Multiplier_0_pp_4_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_10_0 (.A0(Multiplier_0_mult_10_0_n0), .A1(rega_a_1), 
          .A2(Multiplier_0_mult_10_0_n1), .A3(rega_a_2), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(Multiplier_0_cin_lr_10), 
          .CO(mco_25), .P0(Multiplier_0_pp_5_11), .P1(Multiplier_0_pp_5_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_10_1 (.A0(Multiplier_0_mult_10_1_n0), .A1(rega_a_3), 
          .A2(Multiplier_0_mult_10_1_n1), .A3(rega_a_4), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_25), 
          .CO(mco_26), .P0(Multiplier_0_pp_5_13), .P1(Multiplier_0_pp_5_14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_10_2 (.A0(Multiplier_0_mult_10_2_n0), .A1(rega_a_5), 
          .A2(Multiplier_0_mult_10_2_n1), .A3(rega_a_6), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_26), 
          .CO(mco_27), .P0(Multiplier_0_pp_5_15), .P1(Multiplier_0_pp_5_16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_10_3 (.A0(Multiplier_0_mult_10_3_n0), .A1(rega_a_7), 
          .A2(Multiplier_0_mult_10_3_n1), .A3(rega_a_8), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_27), 
          .CO(mco_28), .P0(Multiplier_0_pp_5_17), .P1(Multiplier_0_pp_5_18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_10_4 (.A0(Multiplier_0_mult_10_4_n0), .A1(rega_a_9), 
          .A2(Multiplier_0_mult_10_4_n1), .A3(rega_a_10), .B0(VCC_net), 
          .B1(regb_b_10), .B2(VCC_net), .B3(regb_b_10), .CI(mco_28), 
          .CO(mco_29), .P0(Multiplier_0_pp_5_19), .P1(Multiplier_0_pp_5_20)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    MULT2 Multiplier_0_mult_10_5 (.A0(Multiplier_0_mult_10_5_n0), .A1(Multiplier_0_mult_10_5_n2), 
          .A2(rega_a_11), .A3(GND_net), .B0(VCC_net), .B1(VCC_net), 
          .B2(regb_b_11), .B3(regb_b_10), .CI(mco_29), .CO(mfco_5), 
          .P0(Multiplier_0_pp_5_21), .P1(Multiplier_0_pp_5_22)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t26 (.A(rega_a_11), .B(regb_b_0), .Z(Multiplier_0_mult_0_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    AND2 AND2_t27 (.A(regb_b_0), .B(regb_b_0), .Z(Multiplier_0_pp_0_0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/multiplier.v(376[10:72])
    ND2 ND2_t23 (.A(rega_a_11), .B(regb_b_2), .Z(Multiplier_0_mult_2_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t20 (.A(rega_a_11), .B(regb_b_4), .Z(Multiplier_0_mult_4_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t17 (.A(rega_a_11), .B(regb_b_6), .Z(Multiplier_0_mult_6_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t14 (.A(rega_a_11), .B(regb_b_8), .Z(Multiplier_0_mult_8_5_n2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    ND2 ND2_t11 (.A(rega_a_1), .B(regb_b_11), .Z(Multiplier_0_mult_10_0_n1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=69, LSE_RLINE=75 */ ;   // c:/users/user/lattice/1bitadcfpgasdr/amdemod.v(69[14] 75[27])
    
endmodule
